module sha256_unrolled_pipelined (clk,
    ready,
    reset,
    hashvalue,
    message);
 input clk;
 output ready;
 input reset;
 output [255:0] hashvalue;
 input [0:511] message;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire net629;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire net557;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire net556;
 wire net555;
 wire net554;
 wire net553;
 wire net552;
 wire net551;
 wire net550;
 wire net549;
 wire net548;
 wire _02714_;
 wire net547;
 wire net546;
 wire _02717_;
 wire _02718_;
 wire net545;
 wire net544;
 wire net543;
 wire _02722_;
 wire net542;
 wire net541;
 wire net540;
 wire net539;
 wire net538;
 wire _02728_;
 wire _02729_;
 wire net537;
 wire net536;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire net535;
 wire net534;
 wire _02738_;
 wire net533;
 wire net532;
 wire net531;
 wire _02742_;
 wire net530;
 wire net529;
 wire _02745_;
 wire net528;
 wire net527;
 wire _02748_;
 wire net526;
 wire net525;
 wire _02751_;
 wire net524;
 wire net523;
 wire _02754_;
 wire net522;
 wire _02756_;
 wire net521;
 wire net520;
 wire _02759_;
 wire net519;
 wire net518;
 wire _02762_;
 wire net517;
 wire net516;
 wire _02765_;
 wire net515;
 wire net514;
 wire _02768_;
 wire net513;
 wire _02770_;
 wire net512;
 wire _02772_;
 wire net511;
 wire net510;
 wire _02775_;
 wire _02776_;
 wire net509;
 wire net508;
 wire _02779_;
 wire net507;
 wire net506;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire net505;
 wire net504;
 wire net503;
 wire net502;
 wire net501;
 wire net500;
 wire net499;
 wire net498;
 wire net497;
 wire _02799_;
 wire net496;
 wire net495;
 wire net494;
 wire net493;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire net492;
 wire net491;
 wire net490;
 wire net489;
 wire net488;
 wire _02812_;
 wire _02813_;
 wire net487;
 wire net486;
 wire net485;
 wire net484;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire net483;
 wire net482;
 wire _02824_;
 wire net481;
 wire net480;
 wire _02827_;
 wire net479;
 wire net478;
 wire _02830_;
 wire net477;
 wire net476;
 wire _02833_;
 wire net475;
 wire net474;
 wire _02836_;
 wire net473;
 wire net472;
 wire _02839_;
 wire _02840_;
 wire net471;
 wire _02842_;
 wire net470;
 wire net469;
 wire _02845_;
 wire net468;
 wire net467;
 wire _02848_;
 wire net466;
 wire net465;
 wire _02851_;
 wire net464;
 wire _02853_;
 wire net463;
 wire net462;
 wire _02856_;
 wire net461;
 wire net460;
 wire _02859_;
 wire net459;
 wire _02861_;
 wire net458;
 wire _02863_;
 wire net457;
 wire net456;
 wire _02866_;
 wire net455;
 wire net454;
 wire _02869_;
 wire net453;
 wire net452;
 wire _02872_;
 wire net451;
 wire net450;
 wire _02875_;
 wire net449;
 wire net448;
 wire _02878_;
 wire net447;
 wire net446;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire net445;
 wire net444;
 wire net443;
 wire net442;
 wire net441;
 wire net440;
 wire net439;
 wire net438;
 wire _02892_;
 wire net437;
 wire net436;
 wire net435;
 wire net434;
 wire _02897_;
 wire net433;
 wire net432;
 wire _02900_;
 wire net431;
 wire net430;
 wire net429;
 wire _02904_;
 wire net428;
 wire net427;
 wire net426;
 wire net425;
 wire net424;
 wire _02910_;
 wire net423;
 wire net422;
 wire _02913_;
 wire net421;
 wire net420;
 wire _02916_;
 wire net419;
 wire net418;
 wire _02919_;
 wire net417;
 wire net416;
 wire _02922_;
 wire net415;
 wire net414;
 wire _02925_;
 wire net413;
 wire net412;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire net411;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire net410;
 wire _02947_;
 wire _02948_;
 wire net409;
 wire _02950_;
 wire net408;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire net407;
 wire net406;
 wire _02980_;
 wire _02981_;
 wire net405;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire net404;
 wire net403;
 wire _02989_;
 wire net402;
 wire net401;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire net400;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire net399;
 wire net398;
 wire net397;
 wire net396;
 wire net395;
 wire net394;
 wire net393;
 wire net392;
 wire _03026_;
 wire net391;
 wire net390;
 wire net389;
 wire net388;
 wire _03031_;
 wire net387;
 wire net386;
 wire _03034_;
 wire net385;
 wire net384;
 wire net383;
 wire _03038_;
 wire net382;
 wire net381;
 wire net380;
 wire net379;
 wire net378;
 wire _03044_;
 wire net377;
 wire net376;
 wire _03047_;
 wire net375;
 wire net374;
 wire _03050_;
 wire net373;
 wire net372;
 wire _03053_;
 wire net371;
 wire net370;
 wire _03056_;
 wire net369;
 wire net368;
 wire _03059_;
 wire net367;
 wire net366;
 wire net365;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire net364;
 wire _03072_;
 wire net363;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire net362;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire net361;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire net360;
 wire net359;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire net358;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire net357;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire net356;
 wire net355;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire net354;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire net353;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire net352;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire net351;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire net350;
 wire _03283_;
 wire _03284_;
 wire net349;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire net348;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire net347;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire net346;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire net345;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire net344;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire net343;
 wire _03425_;
 wire net342;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire net341;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire net340;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire net339;
 wire _03484_;
 wire net338;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire net337;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire net336;
 wire _03537_;
 wire net335;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire net334;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire net333;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire net332;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire net331;
 wire _03604_;
 wire net330;
 wire _03606_;
 wire net329;
 wire _03608_;
 wire net328;
 wire _03610_;
 wire net327;
 wire _03612_;
 wire net326;
 wire _03614_;
 wire net325;
 wire _03616_;
 wire net324;
 wire _03618_;
 wire net323;
 wire _03620_;
 wire net322;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire net321;
 wire net320;
 wire _03670_;
 wire net319;
 wire _03672_;
 wire net318;
 wire _03674_;
 wire net317;
 wire _03676_;
 wire _03677_;
 wire net316;
 wire _03679_;
 wire net315;
 wire _03681_;
 wire net314;
 wire _03683_;
 wire net313;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire net312;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire net311;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire net310;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire net309;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire net308;
 wire net307;
 wire _03781_;
 wire net306;
 wire net305;
 wire _03784_;
 wire net304;
 wire net303;
 wire _03787_;
 wire net302;
 wire net301;
 wire _03790_;
 wire net300;
 wire net299;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire net298;
 wire net297;
 wire _03798_;
 wire net296;
 wire net295;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire net294;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire net293;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire net292;
 wire _03853_;
 wire net291;
 wire net290;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03872_;
 wire _03873_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03968_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04005_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04036_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04081_;
 wire _04083_;
 wire _04085_;
 wire net1143;
 wire _04087_;
 wire net1142;
 wire _04089_;
 wire net1141;
 wire _04091_;
 wire net1140;
 wire _04093_;
 wire net1139;
 wire _04095_;
 wire net1138;
 wire _04097_;
 wire net1137;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire net1136;
 wire net1135;
 wire _04125_;
 wire net1134;
 wire _04127_;
 wire net1133;
 wire _04129_;
 wire net1132;
 wire _04131_;
 wire _04132_;
 wire net1131;
 wire _04134_;
 wire net1130;
 wire _04136_;
 wire net1129;
 wire _04138_;
 wire net1123;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire net1114;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire net1113;
 wire net1106;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire net1105;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire net1104;
 wire net1103;
 wire net1075;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire net1074;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire net1073;
 wire _04389_;
 wire net1102;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire net1101;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire net1100;
 wire _04439_;
 wire net1099;
 wire net1098;
 wire _04442_;
 wire net1097;
 wire net1096;
 wire net1095;
 wire _04446_;
 wire net1094;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire net1093;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire net1092;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire net1091;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire net1090;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire net1089;
 wire net1085;
 wire net1084;
 wire net1083;
 wire net1082;
 wire _04784_;
 wire net1081;
 wire _04786_;
 wire net1112;
 wire net1079;
 wire net1078;
 wire _04790_;
 wire net1072;
 wire net1071;
 wire _04793_;
 wire _04794_;
 wire net1070;
 wire _04796_;
 wire _04797_;
 wire net1069;
 wire net1068;
 wire _04800_;
 wire _04801_;
 wire net1067;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire net1066;
 wire _04807_;
 wire _04808_;
 wire net1065;
 wire _04810_;
 wire net1064;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire net1063;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire net1062;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire net1061;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire net1060;
 wire _04845_;
 wire net1059;
 wire net1058;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire net1057;
 wire _04854_;
 wire net1056;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire net1055;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire net1054;
 wire net1053;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire net1052;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire net1051;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire net1050;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire net1049;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire net1048;
 wire _04913_;
 wire net1047;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire net1046;
 wire _04925_;
 wire net1045;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire clknet_5_31__leaf_clk;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire clknet_5_30__leaf_clk;
 wire _04941_;
 wire clknet_5_29__leaf_clk;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire clknet_5_28__leaf_clk;
 wire _04953_;
 wire clknet_5_27__leaf_clk;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire _04963_;
 wire clknet_5_24__leaf_clk;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire clknet_5_23__leaf_clk;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire clknet_5_22__leaf_clk;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire clknet_5_21__leaf_clk;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire clknet_5_20__leaf_clk;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire clknet_5_19__leaf_clk;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire clknet_5_18__leaf_clk;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire clknet_5_17__leaf_clk;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire clknet_5_16__leaf_clk;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire clknet_5_15__leaf_clk;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire clknet_5_14__leaf_clk;
 wire _05062_;
 wire _05063_;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire clknet_5_9__leaf_clk;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire clknet_5_8__leaf_clk;
 wire _05080_;
 wire _05081_;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire clknet_5_3__leaf_clk;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire clknet_5_2__leaf_clk;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire clknet_5_1__leaf_clk;
 wire _05118_;
 wire clknet_5_0__leaf_clk;
 wire clknet_2_3_0_clk;
 wire _05121_;
 wire _05122_;
 wire clknet_2_2_0_clk;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire clknet_2_1_0_clk;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire clknet_2_0_0_clk;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire clknet_0_clk;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire clknet_leaf_288_clk;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire clknet_leaf_287_clk;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire clknet_leaf_286_clk;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire clknet_leaf_285_clk;
 wire _05175_;
 wire clknet_leaf_284_clk;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire clknet_leaf_283_clk;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_281_clk;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire clknet_leaf_280_clk;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire clknet_leaf_279_clk;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire clknet_leaf_278_clk;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire clknet_leaf_277_clk;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire clknet_leaf_276_clk;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire clknet_leaf_275_clk;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire clknet_leaf_274_clk;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire clknet_leaf_273_clk;
 wire _05269_;
 wire clknet_leaf_272_clk;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire clknet_leaf_271_clk;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_269_clk;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire clknet_leaf_268_clk;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire clknet_leaf_267_clk;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire clknet_leaf_266_clk;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire clknet_leaf_265_clk;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire clknet_leaf_264_clk;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire clknet_leaf_263_clk;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire clknet_leaf_262_clk;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire clknet_leaf_261_clk;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire clknet_leaf_260_clk;
 wire _05382_;
 wire clknet_leaf_259_clk;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire clknet_leaf_258_clk;
 wire _05432_;
 wire _05433_;
 wire clknet_leaf_257_clk;
 wire _05435_;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_255_clk;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire clknet_leaf_254_clk;
 wire _05447_;
 wire _05448_;
 wire clknet_leaf_253_clk;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire clknet_leaf_252_clk;
 wire _05459_;
 wire _05460_;
 wire clknet_leaf_251_clk;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_249_clk;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire clknet_leaf_248_clk;
 wire _05488_;
 wire clknet_leaf_247_clk;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire clknet_leaf_246_clk;
 wire _05500_;
 wire clknet_leaf_245_clk;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_243_clk;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire clknet_leaf_242_clk;
 wire _05518_;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_240_clk;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire clknet_leaf_239_clk;
 wire _05530_;
 wire _05531_;
 wire clknet_leaf_238_clk;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire clknet_leaf_237_clk;
 wire _05542_;
 wire _05543_;
 wire clknet_leaf_236_clk;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_234_clk;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire clknet_leaf_233_clk;
 wire _05571_;
 wire clknet_leaf_232_clk;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire clknet_leaf_231_clk;
 wire _05583_;
 wire clknet_leaf_230_clk;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire clknet_leaf_229_clk;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire clknet_leaf_228_clk;
 wire _05600_;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_226_clk;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire clknet_leaf_225_clk;
 wire _05612_;
 wire _05613_;
 wire clknet_leaf_224_clk;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire clknet_leaf_223_clk;
 wire _05624_;
 wire _05625_;
 wire clknet_leaf_222_clk;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_220_clk;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire clknet_leaf_219_clk;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire clknet_leaf_218_clk;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire clknet_leaf_217_clk;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_215_clk;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire clknet_leaf_214_clk;
 wire _05690_;
 wire _05691_;
 wire clknet_leaf_213_clk;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire clknet_leaf_212_clk;
 wire _05702_;
 wire _05703_;
 wire clknet_leaf_211_clk;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_209_clk;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire clknet_leaf_208_clk;
 wire _05730_;
 wire clknet_leaf_207_clk;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire clknet_leaf_206_clk;
 wire _05742_;
 wire clknet_leaf_205_clk;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_203_clk;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire clknet_leaf_202_clk;
 wire _05768_;
 wire _05769_;
 wire clknet_leaf_201_clk;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire clknet_leaf_200_clk;
 wire _05780_;
 wire _05781_;
 wire clknet_leaf_199_clk;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_197_clk;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire clknet_leaf_196_clk;
 wire _05808_;
 wire clknet_leaf_195_clk;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire clknet_leaf_194_clk;
 wire _05820_;
 wire clknet_leaf_193_clk;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_191_clk;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire clknet_leaf_190_clk;
 wire _05846_;
 wire _05847_;
 wire clknet_leaf_189_clk;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire clknet_leaf_188_clk;
 wire _05858_;
 wire _05859_;
 wire clknet_leaf_187_clk;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_185_clk;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire clknet_leaf_184_clk;
 wire _05886_;
 wire clknet_leaf_183_clk;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire clknet_leaf_182_clk;
 wire _05898_;
 wire clknet_leaf_181_clk;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_179_clk;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire clknet_leaf_178_clk;
 wire _05924_;
 wire _05925_;
 wire clknet_leaf_177_clk;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire clknet_leaf_176_clk;
 wire _05936_;
 wire _05937_;
 wire clknet_leaf_175_clk;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_173_clk;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire clknet_leaf_172_clk;
 wire _05965_;
 wire clknet_leaf_171_clk;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire clknet_leaf_170_clk;
 wire _05977_;
 wire clknet_leaf_169_clk;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_162_clk;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_158_clk;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire clknet_leaf_155_clk;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire clknet_leaf_154_clk;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire clknet_leaf_151_clk;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire clknet_leaf_147_clk;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire clknet_leaf_145_clk;
 wire _06237_;
 wire clknet_leaf_144_clk;
 wire _06239_;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_141_clk;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_138_clk;
 wire _06275_;
 wire _06276_;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_136_clk;
 wire _06279_;
 wire _06280_;
 wire clknet_leaf_133_clk;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_124_clk;
 wire _06294_;
 wire clknet_leaf_123_clk;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire clknet_leaf_122_clk;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire clknet_leaf_120_clk;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire clknet_leaf_119_clk;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_117_clk;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire clknet_leaf_116_clk;
 wire _06433_;
 wire clknet_leaf_115_clk;
 wire _06435_;
 wire _06436_;
 wire clknet_leaf_114_clk;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire clknet_leaf_112_clk;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire clknet_leaf_111_clk;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire clknet_leaf_110_clk;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire clknet_leaf_109_clk;
 wire _06462_;
 wire _06463_;
 wire clknet_leaf_108_clk;
 wire _06465_;
 wire clknet_leaf_107_clk;
 wire _06467_;
 wire _06468_;
 wire clknet_leaf_105_clk;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire clknet_leaf_104_clk;
 wire _06474_;
 wire _06475_;
 wire clknet_leaf_103_clk;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire clknet_leaf_102_clk;
 wire _06481_;
 wire _06482_;
 wire clknet_leaf_101_clk;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire clknet_leaf_99_clk;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire clknet_leaf_98_clk;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire clknet_leaf_97_clk;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire clknet_leaf_96_clk;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire clknet_leaf_87_clk;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire clknet_leaf_86_clk;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire clknet_leaf_85_clk;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire clknet_leaf_84_clk;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire clknet_leaf_83_clk;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire clknet_leaf_82_clk;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire clknet_leaf_81_clk;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_77_clk;
 wire _07139_;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_73_clk;
 wire _07144_;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_71_clk;
 wire _07147_;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_68_clk;
 wire _07151_;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_64_clk;
 wire _07156_;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_62_clk;
 wire _07159_;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_60_clk;
 wire _07162_;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_58_clk;
 wire _07165_;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_56_clk;
 wire _07168_;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_54_clk;
 wire _07171_;
 wire clknet_leaf_53_clk;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire clknet_leaf_52_clk;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire clknet_leaf_51_clk;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire clknet_leaf_50_clk;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire clknet_leaf_49_clk;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire clknet_leaf_48_clk;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire clknet_leaf_47_clk;
 wire _07214_;
 wire _07215_;
 wire clknet_leaf_46_clk;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire clknet_leaf_45_clk;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire clknet_leaf_44_clk;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire clknet_leaf_43_clk;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire clknet_leaf_42_clk;
 wire _07242_;
 wire clknet_leaf_41_clk;
 wire _07244_;
 wire clknet_leaf_40_clk;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire clknet_leaf_39_clk;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire clknet_leaf_38_clk;
 wire _07256_;
 wire clknet_leaf_37_clk;
 wire _07258_;
 wire clknet_leaf_36_clk;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire clknet_leaf_35_clk;
 wire _07264_;
 wire clknet_leaf_34_clk;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire clknet_leaf_33_clk;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire clknet_leaf_32_clk;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire clknet_leaf_31_clk;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire clknet_leaf_30_clk;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire clknet_leaf_29_clk;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire clknet_leaf_28_clk;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire clknet_leaf_27_clk;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire clknet_leaf_26_clk;
 wire _07335_;
 wire _07336_;
 wire clknet_leaf_25_clk;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire clknet_leaf_24_clk;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire clknet_leaf_23_clk;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire clknet_leaf_22_clk;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire clknet_leaf_21_clk;
 wire _07363_;
 wire clknet_leaf_20_clk;
 wire _07365_;
 wire clknet_leaf_19_clk;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire clknet_leaf_18_clk;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire clknet_leaf_17_clk;
 wire _07377_;
 wire clknet_leaf_16_clk;
 wire _07379_;
 wire clknet_leaf_15_clk;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire clknet_leaf_14_clk;
 wire _07385_;
 wire clknet_leaf_13_clk;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire clknet_leaf_12_clk;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire clknet_leaf_11_clk;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire clknet_leaf_10_clk;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_6_clk;
 wire _07520_;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_2_clk;
 wire _07525_;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_0_clk;
 wire _07528_;
 wire net1044;
 wire net1043;
 wire net1042;
 wire _07532_;
 wire _07537_;
 wire _07540_;
 wire _07543_;
 wire _07546_;
 wire _07549_;
 wire _07552_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07595_;
 wire _07596_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07623_;
 wire _07625_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07637_;
 wire _07639_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07645_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07716_;
 wire _07717_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07744_;
 wire _07746_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07758_;
 wire _07760_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07766_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08264_;
 wire _08266_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08283_;
 wire _08284_;
 wire _08288_;
 wire _08289_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08301_;
 wire _08302_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08310_;
 wire _08311_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08374_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08573_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08581_;
 wire _08582_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08599_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08622_;
 wire _08623_;
 wire _08625_;
 wire _08626_;
 wire _08629_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08866_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08905_;
 wire _08940_;
 wire _08944_;
 wire _08948_;
 wire _08952_;
 wire _08956_;
 wire _08960_;
 wire _08965_;
 wire _08969_;
 wire _08973_;
 wire _08977_;
 wire _08981_;
 wire _08985_;
 wire _08989_;
 wire _08993_;
 wire _08997_;
 wire _09001_;
 wire _09005_;
 wire _09009_;
 wire _09014_;
 wire net784;
 wire net783;
 wire net782;
 wire net781;
 wire net780;
 wire net779;
 wire net778;
 wire net777;
 wire net776;
 wire net775;
 wire net774;
 wire net773;
 wire net772;
 wire net771;
 wire net770;
 wire net769;
 wire net768;
 wire net767;
 wire net766;
 wire net765;
 wire net764;
 wire net763;
 wire net762;
 wire net761;
 wire net760;
 wire _09050_;
 wire net759;
 wire net758;
 wire net757;
 wire net756;
 wire net755;
 wire net754;
 wire net753;
 wire net752;
 wire net751;
 wire net750;
 wire net749;
 wire net748;
 wire net747;
 wire net746;
 wire net745;
 wire net744;
 wire net743;
 wire net742;
 wire net741;
 wire net740;
 wire net739;
 wire net738;
 wire net737;
 wire net736;
 wire net735;
 wire net734;
 wire net733;
 wire net732;
 wire net731;
 wire net730;
 wire net729;
 wire net728;
 wire net727;
 wire net726;
 wire _09085_;
 wire net725;
 wire net724;
 wire net723;
 wire _09089_;
 wire net722;
 wire net721;
 wire net720;
 wire net719;
 wire _09094_;
 wire net718;
 wire net717;
 wire net716;
 wire _09098_;
 wire net715;
 wire net714;
 wire net713;
 wire _09102_;
 wire net712;
 wire net711;
 wire net710;
 wire _09106_;
 wire net709;
 wire net708;
 wire net707;
 wire _09110_;
 wire net706;
 wire net705;
 wire net704;
 wire _09114_;
 wire net703;
 wire net702;
 wire net701;
 wire _09118_;
 wire net700;
 wire net699;
 wire net698;
 wire _09122_;
 wire net697;
 wire net696;
 wire net695;
 wire _09126_;
 wire net694;
 wire net693;
 wire net692;
 wire _09130_;
 wire net691;
 wire net690;
 wire net689;
 wire _09134_;
 wire net688;
 wire net687;
 wire net686;
 wire _09138_;
 wire net685;
 wire net684;
 wire net683;
 wire _09142_;
 wire net682;
 wire net681;
 wire net680;
 wire _09146_;
 wire net679;
 wire net678;
 wire net677;
 wire _09150_;
 wire net676;
 wire net675;
 wire net674;
 wire _09154_;
 wire net673;
 wire net672;
 wire net671;
 wire net670;
 wire _09159_;
 wire net669;
 wire net668;
 wire net667;
 wire _09163_;
 wire net666;
 wire net665;
 wire net664;
 wire _09167_;
 wire net663;
 wire net662;
 wire net661;
 wire _09171_;
 wire net660;
 wire net659;
 wire net658;
 wire _09175_;
 wire net657;
 wire net656;
 wire net655;
 wire _09179_;
 wire net654;
 wire net653;
 wire net652;
 wire _09183_;
 wire net651;
 wire net650;
 wire net649;
 wire _09187_;
 wire net648;
 wire net647;
 wire net646;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire net645;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire net644;
 wire net643;
 wire net642;
 wire net641;
 wire net640;
 wire net639;
 wire net638;
 wire net637;
 wire net636;
 wire net635;
 wire net634;
 wire net633;
 wire _09726_;
 wire _09727_;
 wire net632;
 wire net631;
 wire net630;
 wire _09731_;
 wire net628;
 wire net627;
 wire net626;
 wire _09735_;
 wire _09736_;
 wire net625;
 wire net624;
 wire _09739_;
 wire _09740_;
 wire net623;
 wire _09742_;
 wire net622;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire net621;
 wire net620;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire net619;
 wire _09766_;
 wire _09767_;
 wire net618;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire net617;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire net616;
 wire _09780_;
 wire net615;
 wire net614;
 wire net613;
 wire _09784_;
 wire net612;
 wire _09786_;
 wire _09787_;
 wire net611;
 wire net610;
 wire _09790_;
 wire _09791_;
 wire net609;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire net608;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire net607;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire net606;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire net605;
 wire _09836_;
 wire net604;
 wire _09838_;
 wire net603;
 wire net602;
 wire net601;
 wire net600;
 wire net599;
 wire _09844_;
 wire net598;
 wire net597;
 wire _09847_;
 wire _09848_;
 wire net596;
 wire net595;
 wire net594;
 wire _09852_;
 wire net593;
 wire _09854_;
 wire net592;
 wire _09856_;
 wire _09857_;
 wire net591;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire net590;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire net589;
 wire net588;
 wire _09870_;
 wire net587;
 wire net586;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire net585;
 wire net584;
 wire net583;
 wire _09879_;
 wire net582;
 wire net581;
 wire net580;
 wire net579;
 wire _09884_;
 wire net578;
 wire net577;
 wire _09887_;
 wire net576;
 wire net575;
 wire _09890_;
 wire net574;
 wire net573;
 wire _09893_;
 wire net572;
 wire net571;
 wire _09896_;
 wire net570;
 wire net569;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire net568;
 wire net567;
 wire _09904_;
 wire net566;
 wire net565;
 wire net564;
 wire _09908_;
 wire net563;
 wire _09910_;
 wire _09911_;
 wire net562;
 wire _09913_;
 wire net561;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire net289;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire net288;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire net287;
 wire _09936_;
 wire _09937_;
 wire net286;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire net285;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire net284;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire net283;
 wire net282;
 wire net281;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire net280;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire net279;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire net278;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire net277;
 wire _09987_;
 wire _09988_;
 wire net276;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire net275;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire net274;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire net273;
 wire net272;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire net271;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire net270;
 wire _10024_;
 wire _10025_;
 wire net269;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire net268;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire net267;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire net266;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire net265;
 wire _10059_;
 wire net264;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire net263;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire net262;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire net261;
 wire _10082_;
 wire _10083_;
 wire net260;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire net259;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire net258;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire net257;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire net256;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire net255;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire net254;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire net253;
 wire _10131_;
 wire _10132_;
 wire net252;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire net251;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire net250;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire net249;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire net248;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire net247;
 wire _10167_;
 wire _10168_;
 wire net246;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire net245;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire net244;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire net243;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire net242;
 wire _10202_;
 wire net241;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire net240;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire net239;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire net238;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire net237;
 wire net236;
 wire net235;
 wire net234;
 wire net233;
 wire net232;
 wire net231;
 wire _10333_;
 wire net230;
 wire net229;
 wire net228;
 wire net227;
 wire _10338_;
 wire net226;
 wire net225;
 wire _10341_;
 wire net224;
 wire net223;
 wire net222;
 wire net221;
 wire _10346_;
 wire net220;
 wire _10348_;
 wire net219;
 wire net218;
 wire _10351_;
 wire _10352_;
 wire net217;
 wire net216;
 wire _10355_;
 wire net215;
 wire net214;
 wire _10358_;
 wire net213;
 wire net212;
 wire _10361_;
 wire net211;
 wire net210;
 wire _10364_;
 wire net209;
 wire net208;
 wire _10367_;
 wire net207;
 wire net206;
 wire net205;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire net204;
 wire net203;
 wire net202;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire net201;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire net200;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire net199;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire net198;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire net197;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire net196;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire net195;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire net194;
 wire _10439_;
 wire _10440_;
 wire net193;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire net192;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire net191;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire net190;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire net189;
 wire _10463_;
 wire _10464_;
 wire net188;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire net187;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire net186;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire net185;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire net184;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire net183;
 wire net182;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire net181;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire net180;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire net179;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire net178;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire net177;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire net176;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire net175;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire net174;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire net173;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire net172;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire net171;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire net170;
 wire _10583_;
 wire _10584_;
 wire net169;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire net168;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire net167;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire net166;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire net165;
 wire _10607_;
 wire _10608_;
 wire net164;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire net163;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire net162;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire net161;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire net160;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire net159;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire net158;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire net157;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire net156;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire net155;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire net154;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire net153;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire net152;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire net151;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire net150;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire net149;
 wire net148;
 wire net147;
 wire net146;
 wire net145;
 wire net144;
 wire net143;
 wire net142;
 wire net141;
 wire _10812_;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire net136;
 wire net135;
 wire net134;
 wire net133;
 wire net132;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire net131;
 wire net130;
 wire _10833_;
 wire net129;
 wire net128;
 wire net127;
 wire _10837_;
 wire net126;
 wire net125;
 wire _10840_;
 wire net124;
 wire net123;
 wire _10843_;
 wire net122;
 wire net121;
 wire _10846_;
 wire net120;
 wire net119;
 wire _10849_;
 wire net118;
 wire _10851_;
 wire net117;
 wire net116;
 wire _10854_;
 wire net115;
 wire net114;
 wire _10857_;
 wire net113;
 wire net112;
 wire _10860_;
 wire net111;
 wire net110;
 wire _10863_;
 wire net109;
 wire _10865_;
 wire net108;
 wire net107;
 wire _10868_;
 wire net106;
 wire net105;
 wire _10871_;
 wire net104;
 wire _10873_;
 wire net103;
 wire _10875_;
 wire net102;
 wire net101;
 wire _10878_;
 wire net100;
 wire net99;
 wire _10881_;
 wire net98;
 wire net97;
 wire _10884_;
 wire net96;
 wire _10886_;
 wire net95;
 wire net94;
 wire _10889_;
 wire net93;
 wire net92;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire net91;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire _10940_;
 wire net80;
 wire net79;
 wire _10943_;
 wire _10944_;
 wire net78;
 wire net77;
 wire _10947_;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire _10953_;
 wire _10954_;
 wire net71;
 wire net70;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire net69;
 wire net68;
 wire _10963_;
 wire net67;
 wire net66;
 wire net65;
 wire _10967_;
 wire net64;
 wire net63;
 wire _10970_;
 wire net62;
 wire net61;
 wire _10973_;
 wire net60;
 wire net59;
 wire _10976_;
 wire net58;
 wire net57;
 wire _10979_;
 wire net56;
 wire net55;
 wire _10982_;
 wire net54;
 wire _10984_;
 wire net53;
 wire net52;
 wire _10987_;
 wire net51;
 wire net50;
 wire _10990_;
 wire net49;
 wire net48;
 wire _10993_;
 wire net47;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire net46;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire net45;
 wire _11017_;
 wire net44;
 wire net43;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire net42;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire net41;
 wire _11059_;
 wire _11060_;
 wire net40;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire net39;
 wire _11070_;
 wire _11071_;
 wire net38;
 wire _11073_;
 wire net37;
 wire _11075_;
 wire _11076_;
 wire net36;
 wire net35;
 wire _11079_;
 wire net34;
 wire net33;
 wire _11082_;
 wire _11083_;
 wire net32;
 wire net31;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire net30;
 wire net29;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire net28;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire net27;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire net26;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire net25;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire net24;
 wire net23;
 wire _11140_;
 wire _11141_;
 wire net22;
 wire _11143_;
 wire net21;
 wire _11145_;
 wire net20;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire net19;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire net18;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire net17;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire net16;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire net15;
 wire net14;
 wire _11515_;
 wire net13;
 wire net12;
 wire _11518_;
 wire net11;
 wire net10;
 wire _11521_;
 wire net9;
 wire net8;
 wire _11524_;
 wire net7;
 wire net6;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire net5;
 wire net4;
 wire _11532_;
 wire net3;
 wire net2;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire net1;
 wire net560;
 wire _11541_;
 wire net559;
 wire net558;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire clknet_leaf_121_clk;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire clknet_leaf_88_clk;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire clknet_leaf_129_clk;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire \count15_1[1] ;
 wire \count15_1[2] ;
 wire \count15_1[3] ;
 wire \count15_1[4] ;
 wire \count15_1[5] ;
 wire \count15_2[1] ;
 wire \count15_2[2] ;
 wire \count15_2[3] ;
 wire \count15_2[4] ;
 wire \count15_2[5] ;
 wire \count16_1[1] ;
 wire \count16_1[2] ;
 wire \count16_1[3] ;
 wire \count16_1[4] ;
 wire \count16_1[5] ;
 wire \count16_2[1] ;
 wire \count16_2[2] ;
 wire \count16_2[3] ;
 wire \count16_2[4] ;
 wire \count16_2[5] ;
 wire \count2_1[1] ;
 wire \count2_1[2] ;
 wire \count2_1[3] ;
 wire \count2_1[4] ;
 wire \count2_1[5] ;
 wire \count2_2[1] ;
 wire \count2_2[2] ;
 wire \count2_2[3] ;
 wire \count2_2[4] ;
 wire \count2_2[5] ;
 wire \count7_1[1] ;
 wire \count7_1[2] ;
 wire \count7_1[3] ;
 wire \count7_1[4] ;
 wire \count7_1[5] ;
 wire \count7_2[1] ;
 wire \count7_2[2] ;
 wire \count7_2[3] ;
 wire \count7_2[4] ;
 wire \count7_2[5] ;
 wire \count_1[1] ;
 wire \count_1[2] ;
 wire \count_1[3] ;
 wire \count_1[4] ;
 wire \count_1[5] ;
 wire \count_2[1] ;
 wire \count_2[2] ;
 wire \count_2[3] ;
 wire \count_2[4] ;
 wire \count_2[5] ;
 wire \count_2[6] ;
 wire \count_hash1[1] ;
 wire \count_hash1[2] ;
 wire \count_hash1[3] ;
 wire \count_hash1[4] ;
 wire \count_hash1[5] ;
 wire \count_hash1[6] ;
 wire \count_hash2[1] ;
 wire \count_hash2[2] ;
 wire \count_hash2[3] ;
 wire \count_hash2[4] ;
 wire \count_hash2[5] ;
 wire done;
 wire \hash.CA1.S0.X[0] ;
 wire \hash.CA1.S0.X[10] ;
 wire \hash.CA1.S0.X[11] ;
 wire \hash.CA1.S0.X[12] ;
 wire \hash.CA1.S0.X[13] ;
 wire \hash.CA1.S0.X[14] ;
 wire \hash.CA1.S0.X[15] ;
 wire \hash.CA1.S0.X[16] ;
 wire \hash.CA1.S0.X[17] ;
 wire \hash.CA1.S0.X[18] ;
 wire \hash.CA1.S0.X[19] ;
 wire \hash.CA1.S0.X[1] ;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_152_clk;
 wire \hash.CA1.S0.X[22] ;
 wire \hash.CA1.S0.X[23] ;
 wire clknet_leaf_150_clk;
 wire \hash.CA1.S0.X[25] ;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_148_clk;
 wire \hash.CA1.S0.X[28] ;
 wire \hash.CA1.S0.X[29] ;
 wire \hash.CA1.S0.X[2] ;
 wire clknet_leaf_146_clk;
 wire \hash.CA1.S0.X[31] ;
 wire \hash.CA1.S0.X[3] ;
 wire clknet_leaf_157_clk;
 wire \hash.CA1.S0.X[5] ;
 wire \hash.CA1.S0.X[6] ;
 wire \hash.CA1.S0.X[7] ;
 wire clknet_leaf_156_clk;
 wire \hash.CA1.S0.X[9] ;
 wire \hash.CA1.S1.X[0] ;
 wire \hash.CA1.S1.X[10] ;
 wire clknet_leaf_94_clk;
 wire \hash.CA1.S1.X[12] ;
 wire \hash.CA1.S1.X[13] ;
 wire \hash.CA1.S1.X[14] ;
 wire clknet_leaf_93_clk;
 wire \hash.CA1.S1.X[16] ;
 wire \hash.CA1.S1.X[17] ;
 wire \hash.CA1.S1.X[18] ;
 wire \hash.CA1.S1.X[19] ;
 wire \hash.CA1.S1.X[1] ;
 wire \hash.CA1.S1.X[20] ;
 wire \hash.CA1.S1.X[21] ;
 wire \hash.CA1.S1.X[22] ;
 wire \hash.CA1.S1.X[23] ;
 wire \hash.CA1.S1.X[24] ;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_89_clk;
 wire \hash.CA1.S1.X[29] ;
 wire \hash.CA1.S1.X[2] ;
 wire \hash.CA1.S1.X[30] ;
 wire \hash.CA1.S1.X[31] ;
 wire \hash.CA1.S1.X[3] ;
 wire \hash.CA1.S1.X[4] ;
 wire \hash.CA1.S1.X[5] ;
 wire \hash.CA1.S1.X[6] ;
 wire \hash.CA1.S1.X[7] ;
 wire clknet_leaf_95_clk;
 wire \hash.CA1.S1.X[9] ;
 wire \hash.CA1.b[0] ;
 wire \hash.CA1.b[10] ;
 wire \hash.CA1.b[11] ;
 wire clknet_leaf_132_clk;
 wire \hash.CA1.b[13] ;
 wire \hash.CA1.b[14] ;
 wire \hash.CA1.b[15] ;
 wire \hash.CA1.b[16] ;
 wire \hash.CA1.b[17] ;
 wire \hash.CA1.b[18] ;
 wire clknet_leaf_131_clk;
 wire \hash.CA1.b[1] ;
 wire \hash.CA1.b[20] ;
 wire \hash.CA1.b[21] ;
 wire \hash.CA1.b[22] ;
 wire clknet_leaf_130_clk;
 wire \hash.CA1.b[24] ;
 wire \hash.CA1.b[25] ;
 wire \hash.CA1.b[26] ;
 wire \hash.CA1.b[27] ;
 wire \hash.CA1.b[28] ;
 wire \hash.CA1.b[29] ;
 wire \hash.CA1.b[2] ;
 wire \hash.CA1.b[30] ;
 wire \hash.CA1.b[31] ;
 wire \hash.CA1.b[3] ;
 wire \hash.CA1.b[4] ;
 wire \hash.CA1.b[5] ;
 wire \hash.CA1.b[6] ;
 wire \hash.CA1.b[7] ;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_134_clk;
 wire \hash.CA1.c[0] ;
 wire \hash.CA1.d[0] ;
 wire \hash.CA1.f[0] ;
 wire \hash.CA1.f[10] ;
 wire \hash.CA1.f[11] ;
 wire \hash.CA1.f[12] ;
 wire \hash.CA1.f[13] ;
 wire \hash.CA1.f[14] ;
 wire \hash.CA1.f[15] ;
 wire \hash.CA1.f[16] ;
 wire \hash.CA1.f[17] ;
 wire clknet_leaf_106_clk;
 wire \hash.CA1.f[19] ;
 wire \hash.CA1.f[1] ;
 wire \hash.CA1.f[20] ;
 wire \hash.CA1.f[21] ;
 wire \hash.CA1.f[22] ;
 wire \hash.CA1.f[23] ;
 wire clknet_leaf_100_clk;
 wire \hash.CA1.f[25] ;
 wire \hash.CA1.f[26] ;
 wire \hash.CA1.f[27] ;
 wire \hash.CA1.f[28] ;
 wire \hash.CA1.f[29] ;
 wire \hash.CA1.f[2] ;
 wire \hash.CA1.f[30] ;
 wire \hash.CA1.f[31] ;
 wire \hash.CA1.f[3] ;
 wire \hash.CA1.f[4] ;
 wire \hash.CA1.f[5] ;
 wire \hash.CA1.f[6] ;
 wire \hash.CA1.f[7] ;
 wire \hash.CA1.f[8] ;
 wire clknet_leaf_113_clk;
 wire \hash.CA1.k_i1[0] ;
 wire \hash.CA1.k_i1[10] ;
 wire \hash.CA1.k_i1[11] ;
 wire \hash.CA1.k_i1[12] ;
 wire \hash.CA1.k_i1[13] ;
 wire \hash.CA1.k_i1[14] ;
 wire \hash.CA1.k_i1[15] ;
 wire \hash.CA1.k_i1[16] ;
 wire \hash.CA1.k_i1[17] ;
 wire \hash.CA1.k_i1[18] ;
 wire \hash.CA1.k_i1[19] ;
 wire \hash.CA1.k_i1[1] ;
 wire \hash.CA1.k_i1[20] ;
 wire \hash.CA1.k_i1[21] ;
 wire \hash.CA1.k_i1[22] ;
 wire \hash.CA1.k_i1[23] ;
 wire \hash.CA1.k_i1[24] ;
 wire \hash.CA1.k_i1[25] ;
 wire \hash.CA1.k_i1[26] ;
 wire \hash.CA1.k_i1[27] ;
 wire \hash.CA1.k_i1[28] ;
 wire \hash.CA1.k_i1[29] ;
 wire \hash.CA1.k_i1[2] ;
 wire \hash.CA1.k_i1[30] ;
 wire \hash.CA1.k_i1[31] ;
 wire \hash.CA1.k_i1[3] ;
 wire \hash.CA1.k_i1[4] ;
 wire \hash.CA1.k_i1[5] ;
 wire \hash.CA1.k_i1[6] ;
 wire \hash.CA1.k_i1[7] ;
 wire \hash.CA1.k_i1[8] ;
 wire \hash.CA1.k_i1[9] ;
 wire \hash.CA1.k_i2[0] ;
 wire \hash.CA1.k_i2[10] ;
 wire \hash.CA1.k_i2[11] ;
 wire \hash.CA1.k_i2[12] ;
 wire \hash.CA1.k_i2[13] ;
 wire \hash.CA1.k_i2[14] ;
 wire \hash.CA1.k_i2[15] ;
 wire \hash.CA1.k_i2[16] ;
 wire \hash.CA1.k_i2[17] ;
 wire \hash.CA1.k_i2[18] ;
 wire \hash.CA1.k_i2[19] ;
 wire \hash.CA1.k_i2[1] ;
 wire \hash.CA1.k_i2[20] ;
 wire \hash.CA1.k_i2[21] ;
 wire \hash.CA1.k_i2[22] ;
 wire \hash.CA1.k_i2[23] ;
 wire \hash.CA1.k_i2[24] ;
 wire \hash.CA1.k_i2[25] ;
 wire \hash.CA1.k_i2[26] ;
 wire \hash.CA1.k_i2[27] ;
 wire \hash.CA1.k_i2[28] ;
 wire \hash.CA1.k_i2[29] ;
 wire \hash.CA1.k_i2[2] ;
 wire \hash.CA1.k_i2[30] ;
 wire \hash.CA1.k_i2[31] ;
 wire \hash.CA1.k_i2[3] ;
 wire \hash.CA1.k_i2[4] ;
 wire \hash.CA1.k_i2[5] ;
 wire \hash.CA1.k_i2[6] ;
 wire \hash.CA1.k_i2[7] ;
 wire \hash.CA1.k_i2[8] ;
 wire \hash.CA1.k_i2[9] ;
 wire \hash.CA1.p1[0] ;
 wire \hash.CA1.p1[10] ;
 wire \hash.CA1.p1[11] ;
 wire \hash.CA1.p1[12] ;
 wire \hash.CA1.p1[13] ;
 wire \hash.CA1.p1[14] ;
 wire \hash.CA1.p1[15] ;
 wire \hash.CA1.p1[16] ;
 wire \hash.CA1.p1[17] ;
 wire \hash.CA1.p1[18] ;
 wire \hash.CA1.p1[19] ;
 wire \hash.CA1.p1[1] ;
 wire \hash.CA1.p1[20] ;
 wire \hash.CA1.p1[21] ;
 wire \hash.CA1.p1[22] ;
 wire \hash.CA1.p1[23] ;
 wire \hash.CA1.p1[24] ;
 wire \hash.CA1.p1[25] ;
 wire \hash.CA1.p1[26] ;
 wire \hash.CA1.p1[27] ;
 wire \hash.CA1.p1[28] ;
 wire \hash.CA1.p1[29] ;
 wire \hash.CA1.p1[2] ;
 wire \hash.CA1.p1[30] ;
 wire \hash.CA1.p1[31] ;
 wire \hash.CA1.p1[3] ;
 wire \hash.CA1.p1[4] ;
 wire \hash.CA1.p1[5] ;
 wire \hash.CA1.p1[6] ;
 wire \hash.CA1.p1[7] ;
 wire \hash.CA1.p1[8] ;
 wire \hash.CA1.p1[9] ;
 wire \hash.CA1.p2[0] ;
 wire \hash.CA1.p2[10] ;
 wire \hash.CA1.p2[11] ;
 wire \hash.CA1.p2[12] ;
 wire \hash.CA1.p2[13] ;
 wire \hash.CA1.p2[14] ;
 wire \hash.CA1.p2[15] ;
 wire \hash.CA1.p2[16] ;
 wire \hash.CA1.p2[17] ;
 wire \hash.CA1.p2[18] ;
 wire \hash.CA1.p2[19] ;
 wire \hash.CA1.p2[1] ;
 wire \hash.CA1.p2[20] ;
 wire \hash.CA1.p2[21] ;
 wire \hash.CA1.p2[22] ;
 wire \hash.CA1.p2[23] ;
 wire \hash.CA1.p2[24] ;
 wire \hash.CA1.p2[25] ;
 wire \hash.CA1.p2[26] ;
 wire \hash.CA1.p2[27] ;
 wire \hash.CA1.p2[28] ;
 wire \hash.CA1.p2[29] ;
 wire \hash.CA1.p2[2] ;
 wire \hash.CA1.p2[30] ;
 wire \hash.CA1.p2[31] ;
 wire \hash.CA1.p2[3] ;
 wire \hash.CA1.p2[4] ;
 wire \hash.CA1.p2[5] ;
 wire \hash.CA1.p2[6] ;
 wire \hash.CA1.p2[7] ;
 wire \hash.CA1.p2[8] ;
 wire \hash.CA1.p2[9] ;
 wire \hash.CA1.p3[0] ;
 wire \hash.CA1.p3[10] ;
 wire \hash.CA1.p3[11] ;
 wire \hash.CA1.p3[12] ;
 wire \hash.CA1.p3[13] ;
 wire \hash.CA1.p3[14] ;
 wire \hash.CA1.p3[15] ;
 wire \hash.CA1.p3[16] ;
 wire \hash.CA1.p3[17] ;
 wire \hash.CA1.p3[18] ;
 wire \hash.CA1.p3[19] ;
 wire \hash.CA1.p3[1] ;
 wire \hash.CA1.p3[20] ;
 wire \hash.CA1.p3[21] ;
 wire \hash.CA1.p3[22] ;
 wire \hash.CA1.p3[23] ;
 wire \hash.CA1.p3[24] ;
 wire \hash.CA1.p3[25] ;
 wire \hash.CA1.p3[26] ;
 wire \hash.CA1.p3[27] ;
 wire \hash.CA1.p3[28] ;
 wire \hash.CA1.p3[29] ;
 wire \hash.CA1.p3[2] ;
 wire \hash.CA1.p3[30] ;
 wire \hash.CA1.p3[31] ;
 wire \hash.CA1.p3[3] ;
 wire \hash.CA1.p3[4] ;
 wire \hash.CA1.p3[5] ;
 wire \hash.CA1.p3[6] ;
 wire \hash.CA1.p3[7] ;
 wire \hash.CA1.p3[8] ;
 wire \hash.CA1.p3[9] ;
 wire \hash.CA1.p4[0] ;
 wire \hash.CA1.p4[10] ;
 wire \hash.CA1.p4[11] ;
 wire \hash.CA1.p4[12] ;
 wire \hash.CA1.p4[13] ;
 wire \hash.CA1.p4[14] ;
 wire \hash.CA1.p4[15] ;
 wire \hash.CA1.p4[16] ;
 wire \hash.CA1.p4[17] ;
 wire \hash.CA1.p4[18] ;
 wire \hash.CA1.p4[19] ;
 wire \hash.CA1.p4[1] ;
 wire \hash.CA1.p4[20] ;
 wire \hash.CA1.p4[21] ;
 wire \hash.CA1.p4[22] ;
 wire \hash.CA1.p4[23] ;
 wire \hash.CA1.p4[24] ;
 wire \hash.CA1.p4[25] ;
 wire \hash.CA1.p4[26] ;
 wire \hash.CA1.p4[27] ;
 wire \hash.CA1.p4[28] ;
 wire \hash.CA1.p4[29] ;
 wire \hash.CA1.p4[2] ;
 wire \hash.CA1.p4[30] ;
 wire \hash.CA1.p4[31] ;
 wire \hash.CA1.p4[3] ;
 wire \hash.CA1.p4[4] ;
 wire \hash.CA1.p4[5] ;
 wire \hash.CA1.p4[6] ;
 wire \hash.CA1.p4[7] ;
 wire \hash.CA1.p4[8] ;
 wire \hash.CA1.p4[9] ;
 wire \hash.CA1.p5[0] ;
 wire \hash.CA1.p5[10] ;
 wire \hash.CA1.p5[11] ;
 wire \hash.CA1.p5[12] ;
 wire \hash.CA1.p5[13] ;
 wire \hash.CA1.p5[14] ;
 wire \hash.CA1.p5[15] ;
 wire \hash.CA1.p5[16] ;
 wire \hash.CA1.p5[17] ;
 wire \hash.CA1.p5[18] ;
 wire \hash.CA1.p5[19] ;
 wire \hash.CA1.p5[1] ;
 wire \hash.CA1.p5[20] ;
 wire \hash.CA1.p5[21] ;
 wire \hash.CA1.p5[22] ;
 wire \hash.CA1.p5[23] ;
 wire \hash.CA1.p5[24] ;
 wire \hash.CA1.p5[25] ;
 wire \hash.CA1.p5[26] ;
 wire \hash.CA1.p5[27] ;
 wire \hash.CA1.p5[28] ;
 wire \hash.CA1.p5[29] ;
 wire \hash.CA1.p5[2] ;
 wire \hash.CA1.p5[30] ;
 wire \hash.CA1.p5[31] ;
 wire \hash.CA1.p5[3] ;
 wire \hash.CA1.p5[4] ;
 wire \hash.CA1.p5[5] ;
 wire \hash.CA1.p5[6] ;
 wire \hash.CA1.p5[7] ;
 wire \hash.CA1.p5[8] ;
 wire \hash.CA1.p5[9] ;
 wire \hash.CA1.w_i1[0] ;
 wire \hash.CA1.w_i1[10] ;
 wire \hash.CA1.w_i1[11] ;
 wire \hash.CA1.w_i1[12] ;
 wire \hash.CA1.w_i1[13] ;
 wire \hash.CA1.w_i1[14] ;
 wire \hash.CA1.w_i1[15] ;
 wire \hash.CA1.w_i1[16] ;
 wire \hash.CA1.w_i1[17] ;
 wire \hash.CA1.w_i1[18] ;
 wire \hash.CA1.w_i1[19] ;
 wire \hash.CA1.w_i1[1] ;
 wire \hash.CA1.w_i1[20] ;
 wire \hash.CA1.w_i1[21] ;
 wire \hash.CA1.w_i1[22] ;
 wire \hash.CA1.w_i1[23] ;
 wire \hash.CA1.w_i1[24] ;
 wire \hash.CA1.w_i1[25] ;
 wire \hash.CA1.w_i1[26] ;
 wire \hash.CA1.w_i1[27] ;
 wire \hash.CA1.w_i1[28] ;
 wire \hash.CA1.w_i1[29] ;
 wire \hash.CA1.w_i1[2] ;
 wire \hash.CA1.w_i1[30] ;
 wire \hash.CA1.w_i1[31] ;
 wire \hash.CA1.w_i1[3] ;
 wire \hash.CA1.w_i1[4] ;
 wire \hash.CA1.w_i1[5] ;
 wire \hash.CA1.w_i1[6] ;
 wire \hash.CA1.w_i1[7] ;
 wire \hash.CA1.w_i1[8] ;
 wire \hash.CA1.w_i1[9] ;
 wire \hash.CA1.w_i2[0] ;
 wire \hash.CA1.w_i2[10] ;
 wire \hash.CA1.w_i2[11] ;
 wire \hash.CA1.w_i2[12] ;
 wire \hash.CA1.w_i2[13] ;
 wire \hash.CA1.w_i2[14] ;
 wire \hash.CA1.w_i2[15] ;
 wire \hash.CA1.w_i2[16] ;
 wire \hash.CA1.w_i2[17] ;
 wire \hash.CA1.w_i2[18] ;
 wire \hash.CA1.w_i2[19] ;
 wire \hash.CA1.w_i2[1] ;
 wire \hash.CA1.w_i2[20] ;
 wire \hash.CA1.w_i2[21] ;
 wire \hash.CA1.w_i2[22] ;
 wire \hash.CA1.w_i2[23] ;
 wire \hash.CA1.w_i2[24] ;
 wire \hash.CA1.w_i2[25] ;
 wire \hash.CA1.w_i2[26] ;
 wire \hash.CA1.w_i2[27] ;
 wire \hash.CA1.w_i2[28] ;
 wire \hash.CA1.w_i2[29] ;
 wire \hash.CA1.w_i2[2] ;
 wire \hash.CA1.w_i2[30] ;
 wire \hash.CA1.w_i2[31] ;
 wire \hash.CA1.w_i2[3] ;
 wire \hash.CA1.w_i2[4] ;
 wire \hash.CA1.w_i2[5] ;
 wire \hash.CA1.w_i2[6] ;
 wire \hash.CA1.w_i2[7] ;
 wire \hash.CA1.w_i2[8] ;
 wire \hash.CA1.w_i2[9] ;
 wire \hash.CA2.S1.X[0] ;
 wire \hash.CA2.S1.X[10] ;
 wire \hash.CA2.S1.X[11] ;
 wire \hash.CA2.S1.X[12] ;
 wire \hash.CA2.S1.X[13] ;
 wire \hash.CA2.S1.X[14] ;
 wire \hash.CA2.S1.X[15] ;
 wire \hash.CA2.S1.X[16] ;
 wire \hash.CA2.S1.X[17] ;
 wire \hash.CA2.S1.X[18] ;
 wire \hash.CA2.S1.X[19] ;
 wire \hash.CA2.S1.X[1] ;
 wire \hash.CA2.S1.X[20] ;
 wire \hash.CA2.S1.X[21] ;
 wire \hash.CA2.S1.X[22] ;
 wire \hash.CA2.S1.X[23] ;
 wire \hash.CA2.S1.X[24] ;
 wire \hash.CA2.S1.X[25] ;
 wire \hash.CA2.S1.X[26] ;
 wire \hash.CA2.S1.X[27] ;
 wire \hash.CA2.S1.X[28] ;
 wire \hash.CA2.S1.X[29] ;
 wire \hash.CA2.S1.X[2] ;
 wire \hash.CA2.S1.X[30] ;
 wire \hash.CA2.S1.X[31] ;
 wire \hash.CA2.S1.X[3] ;
 wire \hash.CA2.S1.X[4] ;
 wire \hash.CA2.S1.X[5] ;
 wire \hash.CA2.S1.X[6] ;
 wire \hash.CA2.S1.X[7] ;
 wire \hash.CA2.S1.X[8] ;
 wire \hash.CA2.S1.X[9] ;
 wire \hash.CA2.a_dash[0] ;
 wire \hash.CA2.a_dash[10] ;
 wire \hash.CA2.a_dash[11] ;
 wire \hash.CA2.a_dash[12] ;
 wire \hash.CA2.a_dash[13] ;
 wire \hash.CA2.a_dash[14] ;
 wire \hash.CA2.a_dash[15] ;
 wire \hash.CA2.a_dash[16] ;
 wire \hash.CA2.a_dash[17] ;
 wire \hash.CA2.a_dash[18] ;
 wire \hash.CA2.a_dash[19] ;
 wire \hash.CA2.a_dash[1] ;
 wire \hash.CA2.a_dash[20] ;
 wire \hash.CA2.a_dash[21] ;
 wire \hash.CA2.a_dash[22] ;
 wire \hash.CA2.a_dash[23] ;
 wire \hash.CA2.a_dash[24] ;
 wire \hash.CA2.a_dash[25] ;
 wire \hash.CA2.a_dash[26] ;
 wire \hash.CA2.a_dash[27] ;
 wire \hash.CA2.a_dash[28] ;
 wire \hash.CA2.a_dash[29] ;
 wire \hash.CA2.a_dash[2] ;
 wire \hash.CA2.a_dash[30] ;
 wire \hash.CA2.a_dash[31] ;
 wire \hash.CA2.a_dash[3] ;
 wire \hash.CA2.a_dash[4] ;
 wire \hash.CA2.a_dash[5] ;
 wire \hash.CA2.a_dash[6] ;
 wire \hash.CA2.a_dash[7] ;
 wire \hash.CA2.a_dash[8] ;
 wire \hash.CA2.a_dash[9] ;
 wire \hash.CA2.b_dash[0] ;
 wire \hash.CA2.b_dash[10] ;
 wire \hash.CA2.b_dash[11] ;
 wire \hash.CA2.b_dash[12] ;
 wire \hash.CA2.b_dash[13] ;
 wire \hash.CA2.b_dash[14] ;
 wire \hash.CA2.b_dash[15] ;
 wire \hash.CA2.b_dash[16] ;
 wire \hash.CA2.b_dash[17] ;
 wire \hash.CA2.b_dash[18] ;
 wire \hash.CA2.b_dash[19] ;
 wire \hash.CA2.b_dash[1] ;
 wire \hash.CA2.b_dash[20] ;
 wire \hash.CA2.b_dash[21] ;
 wire \hash.CA2.b_dash[22] ;
 wire \hash.CA2.b_dash[23] ;
 wire \hash.CA2.b_dash[24] ;
 wire \hash.CA2.b_dash[25] ;
 wire \hash.CA2.b_dash[26] ;
 wire \hash.CA2.b_dash[27] ;
 wire \hash.CA2.b_dash[28] ;
 wire \hash.CA2.b_dash[29] ;
 wire \hash.CA2.b_dash[2] ;
 wire \hash.CA2.b_dash[30] ;
 wire \hash.CA2.b_dash[31] ;
 wire \hash.CA2.b_dash[3] ;
 wire \hash.CA2.b_dash[4] ;
 wire \hash.CA2.b_dash[5] ;
 wire \hash.CA2.b_dash[6] ;
 wire \hash.CA2.b_dash[7] ;
 wire \hash.CA2.b_dash[8] ;
 wire \hash.CA2.b_dash[9] ;
 wire \hash.CA2.e_dash[0] ;
 wire \hash.CA2.e_dash[10] ;
 wire \hash.CA2.e_dash[11] ;
 wire \hash.CA2.e_dash[12] ;
 wire \hash.CA2.e_dash[13] ;
 wire \hash.CA2.e_dash[14] ;
 wire \hash.CA2.e_dash[15] ;
 wire \hash.CA2.e_dash[16] ;
 wire \hash.CA2.e_dash[17] ;
 wire \hash.CA2.e_dash[18] ;
 wire \hash.CA2.e_dash[19] ;
 wire \hash.CA2.e_dash[1] ;
 wire \hash.CA2.e_dash[20] ;
 wire \hash.CA2.e_dash[21] ;
 wire \hash.CA2.e_dash[22] ;
 wire \hash.CA2.e_dash[23] ;
 wire \hash.CA2.e_dash[24] ;
 wire \hash.CA2.e_dash[25] ;
 wire \hash.CA2.e_dash[26] ;
 wire \hash.CA2.e_dash[27] ;
 wire \hash.CA2.e_dash[28] ;
 wire \hash.CA2.e_dash[29] ;
 wire \hash.CA2.e_dash[2] ;
 wire \hash.CA2.e_dash[30] ;
 wire \hash.CA2.e_dash[31] ;
 wire \hash.CA2.e_dash[3] ;
 wire \hash.CA2.e_dash[4] ;
 wire \hash.CA2.e_dash[5] ;
 wire \hash.CA2.e_dash[6] ;
 wire \hash.CA2.e_dash[7] ;
 wire \hash.CA2.e_dash[8] ;
 wire \hash.CA2.e_dash[9] ;
 wire \hash.CA2.f_dash[0] ;
 wire \hash.CA2.f_dash[10] ;
 wire \hash.CA2.f_dash[11] ;
 wire \hash.CA2.f_dash[12] ;
 wire \hash.CA2.f_dash[13] ;
 wire \hash.CA2.f_dash[14] ;
 wire \hash.CA2.f_dash[15] ;
 wire \hash.CA2.f_dash[16] ;
 wire \hash.CA2.f_dash[17] ;
 wire \hash.CA2.f_dash[18] ;
 wire \hash.CA2.f_dash[19] ;
 wire \hash.CA2.f_dash[1] ;
 wire \hash.CA2.f_dash[20] ;
 wire \hash.CA2.f_dash[21] ;
 wire \hash.CA2.f_dash[22] ;
 wire \hash.CA2.f_dash[23] ;
 wire \hash.CA2.f_dash[24] ;
 wire \hash.CA2.f_dash[25] ;
 wire \hash.CA2.f_dash[26] ;
 wire \hash.CA2.f_dash[27] ;
 wire \hash.CA2.f_dash[28] ;
 wire \hash.CA2.f_dash[29] ;
 wire \hash.CA2.f_dash[2] ;
 wire \hash.CA2.f_dash[30] ;
 wire \hash.CA2.f_dash[31] ;
 wire \hash.CA2.f_dash[3] ;
 wire \hash.CA2.f_dash[4] ;
 wire \hash.CA2.f_dash[5] ;
 wire \hash.CA2.f_dash[6] ;
 wire \hash.CA2.f_dash[7] ;
 wire \hash.CA2.f_dash[8] ;
 wire \hash.CA2.f_dash[9] ;
 wire \hash.CA2.p1[0] ;
 wire \hash.CA2.p1[10] ;
 wire \hash.CA2.p1[11] ;
 wire \hash.CA2.p1[12] ;
 wire \hash.CA2.p1[13] ;
 wire \hash.CA2.p1[14] ;
 wire \hash.CA2.p1[15] ;
 wire \hash.CA2.p1[16] ;
 wire \hash.CA2.p1[17] ;
 wire \hash.CA2.p1[18] ;
 wire \hash.CA2.p1[19] ;
 wire \hash.CA2.p1[1] ;
 wire \hash.CA2.p1[20] ;
 wire \hash.CA2.p1[21] ;
 wire \hash.CA2.p1[22] ;
 wire \hash.CA2.p1[23] ;
 wire \hash.CA2.p1[24] ;
 wire \hash.CA2.p1[25] ;
 wire \hash.CA2.p1[26] ;
 wire \hash.CA2.p1[27] ;
 wire \hash.CA2.p1[28] ;
 wire \hash.CA2.p1[29] ;
 wire \hash.CA2.p1[2] ;
 wire \hash.CA2.p1[30] ;
 wire \hash.CA2.p1[31] ;
 wire \hash.CA2.p1[3] ;
 wire \hash.CA2.p1[4] ;
 wire \hash.CA2.p1[5] ;
 wire \hash.CA2.p1[6] ;
 wire \hash.CA2.p1[7] ;
 wire \hash.CA2.p1[8] ;
 wire \hash.CA2.p1[9] ;
 wire \hash.CA2.p3[0] ;
 wire \hash.CA2.p3[10] ;
 wire \hash.CA2.p3[11] ;
 wire \hash.CA2.p3[12] ;
 wire \hash.CA2.p3[13] ;
 wire \hash.CA2.p3[14] ;
 wire \hash.CA2.p3[15] ;
 wire \hash.CA2.p3[16] ;
 wire \hash.CA2.p3[17] ;
 wire \hash.CA2.p3[18] ;
 wire \hash.CA2.p3[19] ;
 wire \hash.CA2.p3[1] ;
 wire \hash.CA2.p3[20] ;
 wire \hash.CA2.p3[21] ;
 wire \hash.CA2.p3[22] ;
 wire \hash.CA2.p3[23] ;
 wire \hash.CA2.p3[24] ;
 wire \hash.CA2.p3[25] ;
 wire \hash.CA2.p3[26] ;
 wire \hash.CA2.p3[27] ;
 wire \hash.CA2.p3[28] ;
 wire \hash.CA2.p3[29] ;
 wire \hash.CA2.p3[2] ;
 wire \hash.CA2.p3[30] ;
 wire \hash.CA2.p3[31] ;
 wire \hash.CA2.p3[3] ;
 wire \hash.CA2.p3[4] ;
 wire \hash.CA2.p3[5] ;
 wire \hash.CA2.p3[6] ;
 wire \hash.CA2.p3[7] ;
 wire \hash.CA2.p3[8] ;
 wire \hash.CA2.p3[9] ;
 wire \hash.CA2.p4[0] ;
 wire \hash.CA2.p4[10] ;
 wire \hash.CA2.p4[11] ;
 wire \hash.CA2.p4[12] ;
 wire \hash.CA2.p4[13] ;
 wire \hash.CA2.p4[14] ;
 wire \hash.CA2.p4[15] ;
 wire \hash.CA2.p4[16] ;
 wire \hash.CA2.p4[17] ;
 wire \hash.CA2.p4[18] ;
 wire \hash.CA2.p4[19] ;
 wire \hash.CA2.p4[1] ;
 wire \hash.CA2.p4[20] ;
 wire \hash.CA2.p4[21] ;
 wire \hash.CA2.p4[22] ;
 wire \hash.CA2.p4[23] ;
 wire \hash.CA2.p4[24] ;
 wire \hash.CA2.p4[25] ;
 wire \hash.CA2.p4[26] ;
 wire \hash.CA2.p4[27] ;
 wire \hash.CA2.p4[28] ;
 wire \hash.CA2.p4[29] ;
 wire \hash.CA2.p4[2] ;
 wire \hash.CA2.p4[30] ;
 wire \hash.CA2.p4[31] ;
 wire \hash.CA2.p4[3] ;
 wire \hash.CA2.p4[4] ;
 wire \hash.CA2.p4[5] ;
 wire \hash.CA2.p4[6] ;
 wire \hash.CA2.p4[7] ;
 wire \hash.CA2.p4[8] ;
 wire \hash.CA2.p4[9] ;
 wire \hash.CA2.p5[0] ;
 wire \hash.CA2.p5[10] ;
 wire \hash.CA2.p5[11] ;
 wire \hash.CA2.p5[12] ;
 wire \hash.CA2.p5[13] ;
 wire \hash.CA2.p5[14] ;
 wire \hash.CA2.p5[15] ;
 wire \hash.CA2.p5[16] ;
 wire \hash.CA2.p5[17] ;
 wire \hash.CA2.p5[18] ;
 wire \hash.CA2.p5[19] ;
 wire \hash.CA2.p5[1] ;
 wire \hash.CA2.p5[20] ;
 wire \hash.CA2.p5[21] ;
 wire \hash.CA2.p5[22] ;
 wire \hash.CA2.p5[23] ;
 wire \hash.CA2.p5[24] ;
 wire \hash.CA2.p5[25] ;
 wire \hash.CA2.p5[26] ;
 wire \hash.CA2.p5[27] ;
 wire \hash.CA2.p5[28] ;
 wire \hash.CA2.p5[29] ;
 wire \hash.CA2.p5[2] ;
 wire \hash.CA2.p5[30] ;
 wire \hash.CA2.p5[31] ;
 wire \hash.CA2.p5[3] ;
 wire \hash.CA2.p5[4] ;
 wire \hash.CA2.p5[5] ;
 wire \hash.CA2.p5[6] ;
 wire \hash.CA2.p5[7] ;
 wire \hash.CA2.p5[8] ;
 wire \hash.CA2.p5[9] ;
 wire \hash.reset ;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire ready_dash;
 wire reset_hash;
 wire \w[0][0] ;
 wire \w[0][10] ;
 wire \w[0][11] ;
 wire \w[0][12] ;
 wire \w[0][13] ;
 wire \w[0][14] ;
 wire \w[0][15] ;
 wire \w[0][16] ;
 wire \w[0][17] ;
 wire \w[0][18] ;
 wire \w[0][19] ;
 wire \w[0][1] ;
 wire \w[0][20] ;
 wire \w[0][21] ;
 wire \w[0][22] ;
 wire \w[0][23] ;
 wire \w[0][24] ;
 wire \w[0][25] ;
 wire \w[0][26] ;
 wire \w[0][27] ;
 wire \w[0][28] ;
 wire \w[0][29] ;
 wire \w[0][2] ;
 wire \w[0][30] ;
 wire \w[0][31] ;
 wire \w[0][3] ;
 wire \w[0][4] ;
 wire \w[0][5] ;
 wire \w[0][6] ;
 wire \w[0][7] ;
 wire \w[0][8] ;
 wire \w[0][9] ;
 wire \w[10][0] ;
 wire \w[10][10] ;
 wire \w[10][11] ;
 wire \w[10][12] ;
 wire \w[10][13] ;
 wire \w[10][14] ;
 wire \w[10][15] ;
 wire \w[10][16] ;
 wire \w[10][17] ;
 wire \w[10][18] ;
 wire \w[10][19] ;
 wire \w[10][1] ;
 wire \w[10][20] ;
 wire \w[10][21] ;
 wire \w[10][22] ;
 wire \w[10][23] ;
 wire \w[10][24] ;
 wire \w[10][25] ;
 wire \w[10][26] ;
 wire \w[10][27] ;
 wire \w[10][28] ;
 wire \w[10][29] ;
 wire \w[10][2] ;
 wire \w[10][30] ;
 wire \w[10][31] ;
 wire \w[10][3] ;
 wire \w[10][4] ;
 wire \w[10][5] ;
 wire \w[10][6] ;
 wire \w[10][7] ;
 wire \w[10][8] ;
 wire \w[10][9] ;
 wire \w[11][0] ;
 wire \w[11][10] ;
 wire \w[11][11] ;
 wire \w[11][12] ;
 wire \w[11][13] ;
 wire \w[11][14] ;
 wire \w[11][15] ;
 wire \w[11][16] ;
 wire \w[11][17] ;
 wire \w[11][18] ;
 wire \w[11][19] ;
 wire \w[11][1] ;
 wire \w[11][20] ;
 wire \w[11][21] ;
 wire \w[11][22] ;
 wire \w[11][23] ;
 wire \w[11][24] ;
 wire \w[11][25] ;
 wire \w[11][26] ;
 wire \w[11][27] ;
 wire \w[11][28] ;
 wire \w[11][29] ;
 wire \w[11][2] ;
 wire \w[11][30] ;
 wire \w[11][31] ;
 wire \w[11][3] ;
 wire \w[11][4] ;
 wire \w[11][5] ;
 wire \w[11][6] ;
 wire \w[11][7] ;
 wire \w[11][8] ;
 wire \w[11][9] ;
 wire \w[12][0] ;
 wire \w[12][10] ;
 wire \w[12][11] ;
 wire \w[12][12] ;
 wire \w[12][13] ;
 wire \w[12][14] ;
 wire \w[12][15] ;
 wire \w[12][16] ;
 wire \w[12][17] ;
 wire \w[12][18] ;
 wire \w[12][19] ;
 wire \w[12][1] ;
 wire \w[12][20] ;
 wire \w[12][21] ;
 wire \w[12][22] ;
 wire \w[12][23] ;
 wire \w[12][24] ;
 wire \w[12][25] ;
 wire \w[12][26] ;
 wire \w[12][27] ;
 wire \w[12][28] ;
 wire \w[12][29] ;
 wire \w[12][2] ;
 wire \w[12][30] ;
 wire \w[12][31] ;
 wire \w[12][3] ;
 wire \w[12][4] ;
 wire \w[12][5] ;
 wire \w[12][6] ;
 wire \w[12][7] ;
 wire \w[12][8] ;
 wire \w[12][9] ;
 wire \w[13][0] ;
 wire \w[13][10] ;
 wire \w[13][11] ;
 wire \w[13][12] ;
 wire \w[13][13] ;
 wire \w[13][14] ;
 wire \w[13][15] ;
 wire \w[13][16] ;
 wire \w[13][17] ;
 wire \w[13][18] ;
 wire \w[13][19] ;
 wire \w[13][1] ;
 wire \w[13][20] ;
 wire \w[13][21] ;
 wire \w[13][22] ;
 wire \w[13][23] ;
 wire \w[13][24] ;
 wire \w[13][25] ;
 wire \w[13][26] ;
 wire \w[13][27] ;
 wire \w[13][28] ;
 wire \w[13][29] ;
 wire \w[13][2] ;
 wire \w[13][30] ;
 wire \w[13][31] ;
 wire \w[13][3] ;
 wire \w[13][4] ;
 wire \w[13][5] ;
 wire \w[13][6] ;
 wire \w[13][7] ;
 wire \w[13][8] ;
 wire \w[13][9] ;
 wire \w[14][0] ;
 wire \w[14][10] ;
 wire \w[14][11] ;
 wire \w[14][12] ;
 wire \w[14][13] ;
 wire \w[14][14] ;
 wire \w[14][15] ;
 wire \w[14][16] ;
 wire \w[14][17] ;
 wire \w[14][18] ;
 wire \w[14][19] ;
 wire \w[14][1] ;
 wire \w[14][20] ;
 wire \w[14][21] ;
 wire \w[14][22] ;
 wire \w[14][23] ;
 wire \w[14][24] ;
 wire \w[14][25] ;
 wire \w[14][26] ;
 wire \w[14][27] ;
 wire \w[14][28] ;
 wire \w[14][29] ;
 wire \w[14][2] ;
 wire \w[14][30] ;
 wire \w[14][31] ;
 wire \w[14][3] ;
 wire \w[14][4] ;
 wire \w[14][5] ;
 wire \w[14][6] ;
 wire \w[14][7] ;
 wire \w[14][8] ;
 wire \w[14][9] ;
 wire \w[15][0] ;
 wire \w[15][10] ;
 wire \w[15][11] ;
 wire \w[15][12] ;
 wire \w[15][13] ;
 wire \w[15][14] ;
 wire \w[15][15] ;
 wire \w[15][16] ;
 wire \w[15][17] ;
 wire \w[15][18] ;
 wire \w[15][19] ;
 wire \w[15][1] ;
 wire \w[15][20] ;
 wire \w[15][21] ;
 wire \w[15][22] ;
 wire \w[15][23] ;
 wire \w[15][24] ;
 wire \w[15][25] ;
 wire \w[15][26] ;
 wire \w[15][27] ;
 wire \w[15][28] ;
 wire \w[15][29] ;
 wire \w[15][2] ;
 wire \w[15][30] ;
 wire \w[15][31] ;
 wire \w[15][3] ;
 wire \w[15][4] ;
 wire \w[15][5] ;
 wire \w[15][6] ;
 wire \w[15][7] ;
 wire \w[15][8] ;
 wire \w[15][9] ;
 wire \w[16][0] ;
 wire \w[16][10] ;
 wire \w[16][11] ;
 wire \w[16][12] ;
 wire \w[16][13] ;
 wire \w[16][14] ;
 wire \w[16][15] ;
 wire \w[16][16] ;
 wire \w[16][17] ;
 wire \w[16][18] ;
 wire \w[16][19] ;
 wire \w[16][1] ;
 wire \w[16][20] ;
 wire \w[16][21] ;
 wire \w[16][22] ;
 wire \w[16][23] ;
 wire \w[16][24] ;
 wire \w[16][25] ;
 wire \w[16][26] ;
 wire \w[16][27] ;
 wire \w[16][28] ;
 wire \w[16][29] ;
 wire \w[16][2] ;
 wire \w[16][30] ;
 wire \w[16][31] ;
 wire \w[16][3] ;
 wire \w[16][4] ;
 wire \w[16][5] ;
 wire \w[16][6] ;
 wire \w[16][7] ;
 wire \w[16][8] ;
 wire \w[16][9] ;
 wire \w[17][0] ;
 wire \w[17][10] ;
 wire \w[17][11] ;
 wire \w[17][12] ;
 wire \w[17][13] ;
 wire \w[17][14] ;
 wire \w[17][15] ;
 wire \w[17][16] ;
 wire \w[17][17] ;
 wire \w[17][18] ;
 wire \w[17][19] ;
 wire \w[17][1] ;
 wire \w[17][20] ;
 wire \w[17][21] ;
 wire \w[17][22] ;
 wire \w[17][23] ;
 wire \w[17][24] ;
 wire \w[17][25] ;
 wire \w[17][26] ;
 wire \w[17][27] ;
 wire \w[17][28] ;
 wire \w[17][29] ;
 wire \w[17][2] ;
 wire \w[17][30] ;
 wire \w[17][31] ;
 wire \w[17][3] ;
 wire \w[17][4] ;
 wire \w[17][5] ;
 wire \w[17][6] ;
 wire \w[17][7] ;
 wire \w[17][8] ;
 wire \w[17][9] ;
 wire \w[18][0] ;
 wire \w[18][10] ;
 wire \w[18][11] ;
 wire \w[18][12] ;
 wire \w[18][13] ;
 wire \w[18][14] ;
 wire \w[18][15] ;
 wire \w[18][16] ;
 wire \w[18][17] ;
 wire \w[18][18] ;
 wire \w[18][19] ;
 wire \w[18][1] ;
 wire \w[18][20] ;
 wire \w[18][21] ;
 wire \w[18][22] ;
 wire \w[18][23] ;
 wire \w[18][24] ;
 wire \w[18][25] ;
 wire \w[18][26] ;
 wire \w[18][27] ;
 wire \w[18][28] ;
 wire \w[18][29] ;
 wire \w[18][2] ;
 wire \w[18][30] ;
 wire \w[18][31] ;
 wire \w[18][3] ;
 wire \w[18][4] ;
 wire \w[18][5] ;
 wire \w[18][6] ;
 wire \w[18][7] ;
 wire \w[18][8] ;
 wire \w[18][9] ;
 wire \w[19][0] ;
 wire \w[19][10] ;
 wire \w[19][11] ;
 wire \w[19][12] ;
 wire \w[19][13] ;
 wire \w[19][14] ;
 wire \w[19][15] ;
 wire \w[19][16] ;
 wire \w[19][17] ;
 wire \w[19][18] ;
 wire \w[19][19] ;
 wire \w[19][1] ;
 wire \w[19][20] ;
 wire \w[19][21] ;
 wire \w[19][22] ;
 wire \w[19][23] ;
 wire \w[19][24] ;
 wire \w[19][25] ;
 wire \w[19][26] ;
 wire \w[19][27] ;
 wire \w[19][28] ;
 wire \w[19][29] ;
 wire \w[19][2] ;
 wire \w[19][30] ;
 wire \w[19][31] ;
 wire \w[19][3] ;
 wire \w[19][4] ;
 wire \w[19][5] ;
 wire \w[19][6] ;
 wire \w[19][7] ;
 wire \w[19][8] ;
 wire \w[19][9] ;
 wire \w[1][0] ;
 wire \w[1][10] ;
 wire \w[1][11] ;
 wire \w[1][12] ;
 wire \w[1][13] ;
 wire \w[1][14] ;
 wire \w[1][15] ;
 wire \w[1][16] ;
 wire \w[1][17] ;
 wire \w[1][18] ;
 wire \w[1][19] ;
 wire \w[1][1] ;
 wire \w[1][20] ;
 wire \w[1][21] ;
 wire \w[1][22] ;
 wire \w[1][23] ;
 wire \w[1][24] ;
 wire \w[1][25] ;
 wire \w[1][26] ;
 wire \w[1][27] ;
 wire \w[1][28] ;
 wire \w[1][29] ;
 wire \w[1][2] ;
 wire \w[1][30] ;
 wire \w[1][31] ;
 wire \w[1][3] ;
 wire \w[1][4] ;
 wire \w[1][5] ;
 wire \w[1][6] ;
 wire \w[1][7] ;
 wire \w[1][8] ;
 wire \w[1][9] ;
 wire \w[20][0] ;
 wire \w[20][10] ;
 wire \w[20][11] ;
 wire \w[20][12] ;
 wire \w[20][13] ;
 wire \w[20][14] ;
 wire \w[20][15] ;
 wire \w[20][16] ;
 wire \w[20][17] ;
 wire \w[20][18] ;
 wire \w[20][19] ;
 wire \w[20][1] ;
 wire \w[20][20] ;
 wire \w[20][21] ;
 wire \w[20][22] ;
 wire \w[20][23] ;
 wire \w[20][24] ;
 wire \w[20][25] ;
 wire \w[20][26] ;
 wire \w[20][27] ;
 wire \w[20][28] ;
 wire \w[20][29] ;
 wire \w[20][2] ;
 wire \w[20][30] ;
 wire \w[20][31] ;
 wire \w[20][3] ;
 wire \w[20][4] ;
 wire \w[20][5] ;
 wire \w[20][6] ;
 wire \w[20][7] ;
 wire \w[20][8] ;
 wire \w[20][9] ;
 wire \w[21][0] ;
 wire \w[21][10] ;
 wire \w[21][11] ;
 wire \w[21][12] ;
 wire \w[21][13] ;
 wire \w[21][14] ;
 wire \w[21][15] ;
 wire \w[21][16] ;
 wire \w[21][17] ;
 wire \w[21][18] ;
 wire \w[21][19] ;
 wire \w[21][1] ;
 wire \w[21][20] ;
 wire \w[21][21] ;
 wire \w[21][22] ;
 wire \w[21][23] ;
 wire \w[21][24] ;
 wire \w[21][25] ;
 wire \w[21][26] ;
 wire \w[21][27] ;
 wire \w[21][28] ;
 wire \w[21][29] ;
 wire \w[21][2] ;
 wire \w[21][30] ;
 wire \w[21][31] ;
 wire \w[21][3] ;
 wire \w[21][4] ;
 wire \w[21][5] ;
 wire \w[21][6] ;
 wire \w[21][7] ;
 wire \w[21][8] ;
 wire \w[21][9] ;
 wire \w[22][0] ;
 wire \w[22][10] ;
 wire \w[22][11] ;
 wire \w[22][12] ;
 wire \w[22][13] ;
 wire \w[22][14] ;
 wire \w[22][15] ;
 wire \w[22][16] ;
 wire \w[22][17] ;
 wire \w[22][18] ;
 wire \w[22][19] ;
 wire \w[22][1] ;
 wire \w[22][20] ;
 wire \w[22][21] ;
 wire \w[22][22] ;
 wire \w[22][23] ;
 wire \w[22][24] ;
 wire \w[22][25] ;
 wire \w[22][26] ;
 wire \w[22][27] ;
 wire \w[22][28] ;
 wire \w[22][29] ;
 wire \w[22][2] ;
 wire \w[22][30] ;
 wire \w[22][31] ;
 wire \w[22][3] ;
 wire \w[22][4] ;
 wire \w[22][5] ;
 wire \w[22][6] ;
 wire \w[22][7] ;
 wire \w[22][8] ;
 wire \w[22][9] ;
 wire \w[23][0] ;
 wire \w[23][10] ;
 wire \w[23][11] ;
 wire \w[23][12] ;
 wire \w[23][13] ;
 wire \w[23][14] ;
 wire \w[23][15] ;
 wire \w[23][16] ;
 wire \w[23][17] ;
 wire \w[23][18] ;
 wire \w[23][19] ;
 wire \w[23][1] ;
 wire \w[23][20] ;
 wire \w[23][21] ;
 wire \w[23][22] ;
 wire \w[23][23] ;
 wire \w[23][24] ;
 wire \w[23][25] ;
 wire \w[23][26] ;
 wire \w[23][27] ;
 wire \w[23][28] ;
 wire \w[23][29] ;
 wire \w[23][2] ;
 wire \w[23][30] ;
 wire \w[23][31] ;
 wire \w[23][3] ;
 wire \w[23][4] ;
 wire \w[23][5] ;
 wire \w[23][6] ;
 wire \w[23][7] ;
 wire \w[23][8] ;
 wire \w[23][9] ;
 wire \w[24][0] ;
 wire \w[24][10] ;
 wire \w[24][11] ;
 wire \w[24][12] ;
 wire \w[24][13] ;
 wire \w[24][14] ;
 wire \w[24][15] ;
 wire \w[24][16] ;
 wire \w[24][17] ;
 wire \w[24][18] ;
 wire \w[24][19] ;
 wire \w[24][1] ;
 wire \w[24][20] ;
 wire \w[24][21] ;
 wire \w[24][22] ;
 wire \w[24][23] ;
 wire \w[24][24] ;
 wire \w[24][25] ;
 wire \w[24][26] ;
 wire \w[24][27] ;
 wire \w[24][28] ;
 wire \w[24][29] ;
 wire \w[24][2] ;
 wire \w[24][30] ;
 wire \w[24][31] ;
 wire \w[24][3] ;
 wire \w[24][4] ;
 wire \w[24][5] ;
 wire \w[24][6] ;
 wire \w[24][7] ;
 wire \w[24][8] ;
 wire \w[24][9] ;
 wire \w[25][0] ;
 wire \w[25][10] ;
 wire \w[25][11] ;
 wire \w[25][12] ;
 wire \w[25][13] ;
 wire \w[25][14] ;
 wire \w[25][15] ;
 wire \w[25][16] ;
 wire \w[25][17] ;
 wire \w[25][18] ;
 wire \w[25][19] ;
 wire \w[25][1] ;
 wire \w[25][20] ;
 wire \w[25][21] ;
 wire \w[25][22] ;
 wire \w[25][23] ;
 wire \w[25][24] ;
 wire \w[25][25] ;
 wire \w[25][26] ;
 wire \w[25][27] ;
 wire \w[25][28] ;
 wire \w[25][29] ;
 wire \w[25][2] ;
 wire \w[25][30] ;
 wire \w[25][31] ;
 wire \w[25][3] ;
 wire \w[25][4] ;
 wire \w[25][5] ;
 wire \w[25][6] ;
 wire \w[25][7] ;
 wire \w[25][8] ;
 wire \w[25][9] ;
 wire \w[26][0] ;
 wire \w[26][10] ;
 wire \w[26][11] ;
 wire \w[26][12] ;
 wire \w[26][13] ;
 wire \w[26][14] ;
 wire \w[26][15] ;
 wire \w[26][16] ;
 wire \w[26][17] ;
 wire \w[26][18] ;
 wire \w[26][19] ;
 wire \w[26][1] ;
 wire \w[26][20] ;
 wire \w[26][21] ;
 wire \w[26][22] ;
 wire \w[26][23] ;
 wire \w[26][24] ;
 wire \w[26][25] ;
 wire \w[26][26] ;
 wire \w[26][27] ;
 wire \w[26][28] ;
 wire \w[26][29] ;
 wire \w[26][2] ;
 wire \w[26][30] ;
 wire \w[26][31] ;
 wire \w[26][3] ;
 wire \w[26][4] ;
 wire \w[26][5] ;
 wire \w[26][6] ;
 wire \w[26][7] ;
 wire \w[26][8] ;
 wire \w[26][9] ;
 wire \w[27][0] ;
 wire \w[27][10] ;
 wire \w[27][11] ;
 wire \w[27][12] ;
 wire \w[27][13] ;
 wire \w[27][14] ;
 wire \w[27][15] ;
 wire \w[27][16] ;
 wire \w[27][17] ;
 wire \w[27][18] ;
 wire \w[27][19] ;
 wire \w[27][1] ;
 wire \w[27][20] ;
 wire \w[27][21] ;
 wire \w[27][22] ;
 wire \w[27][23] ;
 wire \w[27][24] ;
 wire \w[27][25] ;
 wire \w[27][26] ;
 wire \w[27][27] ;
 wire \w[27][28] ;
 wire \w[27][29] ;
 wire \w[27][2] ;
 wire \w[27][30] ;
 wire \w[27][31] ;
 wire \w[27][3] ;
 wire \w[27][4] ;
 wire \w[27][5] ;
 wire \w[27][6] ;
 wire \w[27][7] ;
 wire \w[27][8] ;
 wire \w[27][9] ;
 wire \w[28][0] ;
 wire \w[28][10] ;
 wire \w[28][11] ;
 wire \w[28][12] ;
 wire \w[28][13] ;
 wire \w[28][14] ;
 wire \w[28][15] ;
 wire \w[28][16] ;
 wire \w[28][17] ;
 wire \w[28][18] ;
 wire \w[28][19] ;
 wire \w[28][1] ;
 wire \w[28][20] ;
 wire \w[28][21] ;
 wire \w[28][22] ;
 wire \w[28][23] ;
 wire \w[28][24] ;
 wire \w[28][25] ;
 wire \w[28][26] ;
 wire \w[28][27] ;
 wire \w[28][28] ;
 wire \w[28][29] ;
 wire \w[28][2] ;
 wire \w[28][30] ;
 wire \w[28][31] ;
 wire \w[28][3] ;
 wire \w[28][4] ;
 wire \w[28][5] ;
 wire \w[28][6] ;
 wire \w[28][7] ;
 wire \w[28][8] ;
 wire \w[28][9] ;
 wire \w[29][0] ;
 wire \w[29][10] ;
 wire \w[29][11] ;
 wire \w[29][12] ;
 wire \w[29][13] ;
 wire \w[29][14] ;
 wire \w[29][15] ;
 wire \w[29][16] ;
 wire \w[29][17] ;
 wire \w[29][18] ;
 wire \w[29][19] ;
 wire \w[29][1] ;
 wire \w[29][20] ;
 wire \w[29][21] ;
 wire \w[29][22] ;
 wire \w[29][23] ;
 wire \w[29][24] ;
 wire \w[29][25] ;
 wire \w[29][26] ;
 wire \w[29][27] ;
 wire \w[29][28] ;
 wire \w[29][29] ;
 wire \w[29][2] ;
 wire \w[29][30] ;
 wire \w[29][31] ;
 wire \w[29][3] ;
 wire \w[29][4] ;
 wire \w[29][5] ;
 wire \w[29][6] ;
 wire \w[29][7] ;
 wire \w[29][8] ;
 wire \w[29][9] ;
 wire \w[2][0] ;
 wire \w[2][10] ;
 wire \w[2][11] ;
 wire \w[2][12] ;
 wire \w[2][13] ;
 wire \w[2][14] ;
 wire \w[2][15] ;
 wire \w[2][16] ;
 wire \w[2][17] ;
 wire \w[2][18] ;
 wire \w[2][19] ;
 wire \w[2][1] ;
 wire \w[2][20] ;
 wire \w[2][21] ;
 wire \w[2][22] ;
 wire \w[2][23] ;
 wire \w[2][24] ;
 wire \w[2][25] ;
 wire \w[2][26] ;
 wire \w[2][27] ;
 wire \w[2][28] ;
 wire \w[2][29] ;
 wire \w[2][2] ;
 wire \w[2][30] ;
 wire \w[2][31] ;
 wire \w[2][3] ;
 wire \w[2][4] ;
 wire \w[2][5] ;
 wire \w[2][6] ;
 wire \w[2][7] ;
 wire \w[2][8] ;
 wire \w[2][9] ;
 wire \w[30][0] ;
 wire \w[30][10] ;
 wire \w[30][11] ;
 wire \w[30][12] ;
 wire \w[30][13] ;
 wire \w[30][14] ;
 wire \w[30][15] ;
 wire \w[30][16] ;
 wire \w[30][17] ;
 wire \w[30][18] ;
 wire \w[30][19] ;
 wire \w[30][1] ;
 wire \w[30][20] ;
 wire \w[30][21] ;
 wire \w[30][22] ;
 wire \w[30][23] ;
 wire \w[30][24] ;
 wire \w[30][25] ;
 wire \w[30][26] ;
 wire \w[30][27] ;
 wire \w[30][28] ;
 wire \w[30][29] ;
 wire \w[30][2] ;
 wire \w[30][30] ;
 wire \w[30][31] ;
 wire \w[30][3] ;
 wire \w[30][4] ;
 wire \w[30][5] ;
 wire \w[30][6] ;
 wire \w[30][7] ;
 wire \w[30][8] ;
 wire \w[30][9] ;
 wire \w[31][0] ;
 wire \w[31][10] ;
 wire \w[31][11] ;
 wire \w[31][12] ;
 wire \w[31][13] ;
 wire \w[31][14] ;
 wire \w[31][15] ;
 wire \w[31][16] ;
 wire \w[31][17] ;
 wire \w[31][18] ;
 wire \w[31][19] ;
 wire \w[31][1] ;
 wire \w[31][20] ;
 wire \w[31][21] ;
 wire \w[31][22] ;
 wire \w[31][23] ;
 wire \w[31][24] ;
 wire \w[31][25] ;
 wire \w[31][26] ;
 wire \w[31][27] ;
 wire \w[31][28] ;
 wire \w[31][29] ;
 wire \w[31][2] ;
 wire \w[31][30] ;
 wire \w[31][31] ;
 wire \w[31][3] ;
 wire \w[31][4] ;
 wire \w[31][5] ;
 wire \w[31][6] ;
 wire \w[31][7] ;
 wire \w[31][8] ;
 wire \w[31][9] ;
 wire \w[32][0] ;
 wire \w[32][10] ;
 wire \w[32][11] ;
 wire \w[32][12] ;
 wire \w[32][13] ;
 wire \w[32][14] ;
 wire \w[32][15] ;
 wire \w[32][16] ;
 wire \w[32][17] ;
 wire \w[32][18] ;
 wire \w[32][19] ;
 wire \w[32][1] ;
 wire \w[32][20] ;
 wire \w[32][21] ;
 wire \w[32][22] ;
 wire \w[32][23] ;
 wire \w[32][24] ;
 wire \w[32][25] ;
 wire \w[32][26] ;
 wire \w[32][27] ;
 wire \w[32][28] ;
 wire \w[32][29] ;
 wire \w[32][2] ;
 wire \w[32][30] ;
 wire \w[32][31] ;
 wire \w[32][3] ;
 wire \w[32][4] ;
 wire \w[32][5] ;
 wire \w[32][6] ;
 wire \w[32][7] ;
 wire \w[32][8] ;
 wire \w[32][9] ;
 wire \w[33][0] ;
 wire \w[33][10] ;
 wire \w[33][11] ;
 wire \w[33][12] ;
 wire \w[33][13] ;
 wire \w[33][14] ;
 wire \w[33][15] ;
 wire \w[33][16] ;
 wire \w[33][17] ;
 wire \w[33][18] ;
 wire \w[33][19] ;
 wire \w[33][1] ;
 wire \w[33][20] ;
 wire \w[33][21] ;
 wire \w[33][22] ;
 wire \w[33][23] ;
 wire \w[33][24] ;
 wire \w[33][25] ;
 wire \w[33][26] ;
 wire \w[33][27] ;
 wire \w[33][28] ;
 wire \w[33][29] ;
 wire \w[33][2] ;
 wire \w[33][30] ;
 wire \w[33][31] ;
 wire \w[33][3] ;
 wire \w[33][4] ;
 wire \w[33][5] ;
 wire \w[33][6] ;
 wire \w[33][7] ;
 wire \w[33][8] ;
 wire \w[33][9] ;
 wire \w[34][0] ;
 wire \w[34][10] ;
 wire \w[34][11] ;
 wire \w[34][12] ;
 wire \w[34][13] ;
 wire \w[34][14] ;
 wire \w[34][15] ;
 wire \w[34][16] ;
 wire \w[34][17] ;
 wire \w[34][18] ;
 wire \w[34][19] ;
 wire \w[34][1] ;
 wire \w[34][20] ;
 wire \w[34][21] ;
 wire \w[34][22] ;
 wire \w[34][23] ;
 wire \w[34][24] ;
 wire \w[34][25] ;
 wire \w[34][26] ;
 wire \w[34][27] ;
 wire \w[34][28] ;
 wire \w[34][29] ;
 wire \w[34][2] ;
 wire \w[34][30] ;
 wire \w[34][31] ;
 wire \w[34][3] ;
 wire \w[34][4] ;
 wire \w[34][5] ;
 wire \w[34][6] ;
 wire \w[34][7] ;
 wire \w[34][8] ;
 wire \w[34][9] ;
 wire \w[35][0] ;
 wire \w[35][10] ;
 wire \w[35][11] ;
 wire \w[35][12] ;
 wire \w[35][13] ;
 wire \w[35][14] ;
 wire \w[35][15] ;
 wire \w[35][16] ;
 wire \w[35][17] ;
 wire \w[35][18] ;
 wire \w[35][19] ;
 wire \w[35][1] ;
 wire \w[35][20] ;
 wire \w[35][21] ;
 wire \w[35][22] ;
 wire \w[35][23] ;
 wire \w[35][24] ;
 wire \w[35][25] ;
 wire \w[35][26] ;
 wire \w[35][27] ;
 wire \w[35][28] ;
 wire \w[35][29] ;
 wire \w[35][2] ;
 wire \w[35][30] ;
 wire \w[35][31] ;
 wire \w[35][3] ;
 wire \w[35][4] ;
 wire \w[35][5] ;
 wire \w[35][6] ;
 wire \w[35][7] ;
 wire \w[35][8] ;
 wire \w[35][9] ;
 wire \w[36][0] ;
 wire \w[36][10] ;
 wire \w[36][11] ;
 wire \w[36][12] ;
 wire \w[36][13] ;
 wire \w[36][14] ;
 wire \w[36][15] ;
 wire \w[36][16] ;
 wire \w[36][17] ;
 wire \w[36][18] ;
 wire \w[36][19] ;
 wire \w[36][1] ;
 wire \w[36][20] ;
 wire \w[36][21] ;
 wire \w[36][22] ;
 wire \w[36][23] ;
 wire \w[36][24] ;
 wire \w[36][25] ;
 wire \w[36][26] ;
 wire \w[36][27] ;
 wire \w[36][28] ;
 wire \w[36][29] ;
 wire \w[36][2] ;
 wire \w[36][30] ;
 wire \w[36][31] ;
 wire \w[36][3] ;
 wire \w[36][4] ;
 wire \w[36][5] ;
 wire \w[36][6] ;
 wire \w[36][7] ;
 wire \w[36][8] ;
 wire \w[36][9] ;
 wire \w[37][0] ;
 wire \w[37][10] ;
 wire \w[37][11] ;
 wire \w[37][12] ;
 wire \w[37][13] ;
 wire \w[37][14] ;
 wire \w[37][15] ;
 wire \w[37][16] ;
 wire \w[37][17] ;
 wire \w[37][18] ;
 wire \w[37][19] ;
 wire \w[37][1] ;
 wire \w[37][20] ;
 wire \w[37][21] ;
 wire \w[37][22] ;
 wire \w[37][23] ;
 wire \w[37][24] ;
 wire \w[37][25] ;
 wire \w[37][26] ;
 wire \w[37][27] ;
 wire \w[37][28] ;
 wire \w[37][29] ;
 wire \w[37][2] ;
 wire \w[37][30] ;
 wire \w[37][31] ;
 wire \w[37][3] ;
 wire \w[37][4] ;
 wire \w[37][5] ;
 wire \w[37][6] ;
 wire \w[37][7] ;
 wire \w[37][8] ;
 wire \w[37][9] ;
 wire \w[38][0] ;
 wire \w[38][10] ;
 wire \w[38][11] ;
 wire \w[38][12] ;
 wire \w[38][13] ;
 wire \w[38][14] ;
 wire \w[38][15] ;
 wire \w[38][16] ;
 wire \w[38][17] ;
 wire \w[38][18] ;
 wire \w[38][19] ;
 wire \w[38][1] ;
 wire \w[38][20] ;
 wire \w[38][21] ;
 wire \w[38][22] ;
 wire \w[38][23] ;
 wire \w[38][24] ;
 wire \w[38][25] ;
 wire \w[38][26] ;
 wire \w[38][27] ;
 wire \w[38][28] ;
 wire \w[38][29] ;
 wire \w[38][2] ;
 wire \w[38][30] ;
 wire \w[38][31] ;
 wire \w[38][3] ;
 wire \w[38][4] ;
 wire \w[38][5] ;
 wire \w[38][6] ;
 wire \w[38][7] ;
 wire \w[38][8] ;
 wire \w[38][9] ;
 wire \w[39][0] ;
 wire \w[39][10] ;
 wire \w[39][11] ;
 wire \w[39][12] ;
 wire \w[39][13] ;
 wire \w[39][14] ;
 wire \w[39][15] ;
 wire \w[39][16] ;
 wire \w[39][17] ;
 wire \w[39][18] ;
 wire \w[39][19] ;
 wire \w[39][1] ;
 wire \w[39][20] ;
 wire \w[39][21] ;
 wire \w[39][22] ;
 wire \w[39][23] ;
 wire \w[39][24] ;
 wire \w[39][25] ;
 wire \w[39][26] ;
 wire \w[39][27] ;
 wire \w[39][28] ;
 wire \w[39][29] ;
 wire \w[39][2] ;
 wire \w[39][30] ;
 wire \w[39][31] ;
 wire \w[39][3] ;
 wire \w[39][4] ;
 wire \w[39][5] ;
 wire \w[39][6] ;
 wire \w[39][7] ;
 wire \w[39][8] ;
 wire \w[39][9] ;
 wire \w[3][0] ;
 wire \w[3][10] ;
 wire \w[3][11] ;
 wire \w[3][12] ;
 wire \w[3][13] ;
 wire \w[3][14] ;
 wire \w[3][15] ;
 wire \w[3][16] ;
 wire \w[3][17] ;
 wire \w[3][18] ;
 wire \w[3][19] ;
 wire \w[3][1] ;
 wire \w[3][20] ;
 wire \w[3][21] ;
 wire \w[3][22] ;
 wire \w[3][23] ;
 wire \w[3][24] ;
 wire \w[3][25] ;
 wire \w[3][26] ;
 wire \w[3][27] ;
 wire \w[3][28] ;
 wire \w[3][29] ;
 wire \w[3][2] ;
 wire \w[3][30] ;
 wire \w[3][31] ;
 wire \w[3][3] ;
 wire \w[3][4] ;
 wire \w[3][5] ;
 wire \w[3][6] ;
 wire \w[3][7] ;
 wire \w[3][8] ;
 wire \w[3][9] ;
 wire \w[40][0] ;
 wire \w[40][10] ;
 wire \w[40][11] ;
 wire \w[40][12] ;
 wire \w[40][13] ;
 wire \w[40][14] ;
 wire \w[40][15] ;
 wire \w[40][16] ;
 wire \w[40][17] ;
 wire \w[40][18] ;
 wire \w[40][19] ;
 wire \w[40][1] ;
 wire \w[40][20] ;
 wire \w[40][21] ;
 wire \w[40][22] ;
 wire \w[40][23] ;
 wire \w[40][24] ;
 wire \w[40][25] ;
 wire \w[40][26] ;
 wire \w[40][27] ;
 wire \w[40][28] ;
 wire \w[40][29] ;
 wire \w[40][2] ;
 wire \w[40][30] ;
 wire \w[40][31] ;
 wire \w[40][3] ;
 wire \w[40][4] ;
 wire \w[40][5] ;
 wire \w[40][6] ;
 wire \w[40][7] ;
 wire \w[40][8] ;
 wire \w[40][9] ;
 wire \w[41][0] ;
 wire \w[41][10] ;
 wire \w[41][11] ;
 wire \w[41][12] ;
 wire \w[41][13] ;
 wire \w[41][14] ;
 wire \w[41][15] ;
 wire \w[41][16] ;
 wire \w[41][17] ;
 wire \w[41][18] ;
 wire \w[41][19] ;
 wire \w[41][1] ;
 wire \w[41][20] ;
 wire \w[41][21] ;
 wire \w[41][22] ;
 wire \w[41][23] ;
 wire \w[41][24] ;
 wire \w[41][25] ;
 wire \w[41][26] ;
 wire \w[41][27] ;
 wire \w[41][28] ;
 wire \w[41][29] ;
 wire \w[41][2] ;
 wire \w[41][30] ;
 wire \w[41][31] ;
 wire \w[41][3] ;
 wire \w[41][4] ;
 wire \w[41][5] ;
 wire \w[41][6] ;
 wire \w[41][7] ;
 wire \w[41][8] ;
 wire \w[41][9] ;
 wire \w[42][0] ;
 wire \w[42][10] ;
 wire \w[42][11] ;
 wire \w[42][12] ;
 wire \w[42][13] ;
 wire \w[42][14] ;
 wire \w[42][15] ;
 wire \w[42][16] ;
 wire \w[42][17] ;
 wire \w[42][18] ;
 wire \w[42][19] ;
 wire \w[42][1] ;
 wire \w[42][20] ;
 wire \w[42][21] ;
 wire \w[42][22] ;
 wire \w[42][23] ;
 wire \w[42][24] ;
 wire \w[42][25] ;
 wire \w[42][26] ;
 wire \w[42][27] ;
 wire \w[42][28] ;
 wire \w[42][29] ;
 wire \w[42][2] ;
 wire \w[42][30] ;
 wire \w[42][31] ;
 wire \w[42][3] ;
 wire \w[42][4] ;
 wire \w[42][5] ;
 wire \w[42][6] ;
 wire \w[42][7] ;
 wire \w[42][8] ;
 wire \w[42][9] ;
 wire \w[43][0] ;
 wire \w[43][10] ;
 wire \w[43][11] ;
 wire \w[43][12] ;
 wire \w[43][13] ;
 wire \w[43][14] ;
 wire \w[43][15] ;
 wire \w[43][16] ;
 wire \w[43][17] ;
 wire \w[43][18] ;
 wire \w[43][19] ;
 wire \w[43][1] ;
 wire \w[43][20] ;
 wire \w[43][21] ;
 wire \w[43][22] ;
 wire \w[43][23] ;
 wire \w[43][24] ;
 wire \w[43][25] ;
 wire \w[43][26] ;
 wire \w[43][27] ;
 wire \w[43][28] ;
 wire \w[43][29] ;
 wire \w[43][2] ;
 wire \w[43][30] ;
 wire \w[43][31] ;
 wire \w[43][3] ;
 wire \w[43][4] ;
 wire \w[43][5] ;
 wire \w[43][6] ;
 wire \w[43][7] ;
 wire \w[43][8] ;
 wire \w[43][9] ;
 wire \w[44][0] ;
 wire \w[44][10] ;
 wire \w[44][11] ;
 wire \w[44][12] ;
 wire \w[44][13] ;
 wire \w[44][14] ;
 wire \w[44][15] ;
 wire \w[44][16] ;
 wire \w[44][17] ;
 wire \w[44][18] ;
 wire \w[44][19] ;
 wire \w[44][1] ;
 wire \w[44][20] ;
 wire \w[44][21] ;
 wire \w[44][22] ;
 wire \w[44][23] ;
 wire \w[44][24] ;
 wire \w[44][25] ;
 wire \w[44][26] ;
 wire \w[44][27] ;
 wire \w[44][28] ;
 wire \w[44][29] ;
 wire \w[44][2] ;
 wire \w[44][30] ;
 wire \w[44][31] ;
 wire \w[44][3] ;
 wire \w[44][4] ;
 wire \w[44][5] ;
 wire \w[44][6] ;
 wire \w[44][7] ;
 wire \w[44][8] ;
 wire \w[44][9] ;
 wire \w[45][0] ;
 wire \w[45][10] ;
 wire \w[45][11] ;
 wire \w[45][12] ;
 wire \w[45][13] ;
 wire \w[45][14] ;
 wire \w[45][15] ;
 wire \w[45][16] ;
 wire \w[45][17] ;
 wire \w[45][18] ;
 wire \w[45][19] ;
 wire \w[45][1] ;
 wire \w[45][20] ;
 wire \w[45][21] ;
 wire \w[45][22] ;
 wire \w[45][23] ;
 wire \w[45][24] ;
 wire \w[45][25] ;
 wire \w[45][26] ;
 wire \w[45][27] ;
 wire \w[45][28] ;
 wire \w[45][29] ;
 wire \w[45][2] ;
 wire \w[45][30] ;
 wire \w[45][31] ;
 wire \w[45][3] ;
 wire \w[45][4] ;
 wire \w[45][5] ;
 wire \w[45][6] ;
 wire \w[45][7] ;
 wire \w[45][8] ;
 wire \w[45][9] ;
 wire \w[46][0] ;
 wire \w[46][10] ;
 wire \w[46][11] ;
 wire \w[46][12] ;
 wire \w[46][13] ;
 wire \w[46][14] ;
 wire \w[46][15] ;
 wire \w[46][16] ;
 wire \w[46][17] ;
 wire \w[46][18] ;
 wire \w[46][19] ;
 wire \w[46][1] ;
 wire \w[46][20] ;
 wire \w[46][21] ;
 wire \w[46][22] ;
 wire \w[46][23] ;
 wire \w[46][24] ;
 wire \w[46][25] ;
 wire \w[46][26] ;
 wire \w[46][27] ;
 wire \w[46][28] ;
 wire \w[46][29] ;
 wire \w[46][2] ;
 wire \w[46][30] ;
 wire \w[46][31] ;
 wire \w[46][3] ;
 wire \w[46][4] ;
 wire \w[46][5] ;
 wire \w[46][6] ;
 wire \w[46][7] ;
 wire \w[46][8] ;
 wire \w[46][9] ;
 wire \w[47][0] ;
 wire \w[47][10] ;
 wire \w[47][11] ;
 wire \w[47][12] ;
 wire \w[47][13] ;
 wire \w[47][14] ;
 wire \w[47][15] ;
 wire \w[47][16] ;
 wire \w[47][17] ;
 wire \w[47][18] ;
 wire \w[47][19] ;
 wire \w[47][1] ;
 wire \w[47][20] ;
 wire \w[47][21] ;
 wire \w[47][22] ;
 wire \w[47][23] ;
 wire \w[47][24] ;
 wire \w[47][25] ;
 wire \w[47][26] ;
 wire \w[47][27] ;
 wire \w[47][28] ;
 wire \w[47][29] ;
 wire \w[47][2] ;
 wire \w[47][30] ;
 wire \w[47][31] ;
 wire \w[47][3] ;
 wire \w[47][4] ;
 wire \w[47][5] ;
 wire \w[47][6] ;
 wire \w[47][7] ;
 wire \w[47][8] ;
 wire \w[47][9] ;
 wire \w[48][0] ;
 wire \w[48][10] ;
 wire \w[48][11] ;
 wire \w[48][12] ;
 wire \w[48][13] ;
 wire \w[48][14] ;
 wire \w[48][15] ;
 wire \w[48][16] ;
 wire \w[48][17] ;
 wire \w[48][18] ;
 wire \w[48][19] ;
 wire \w[48][1] ;
 wire \w[48][20] ;
 wire \w[48][21] ;
 wire \w[48][22] ;
 wire \w[48][23] ;
 wire \w[48][24] ;
 wire \w[48][25] ;
 wire \w[48][26] ;
 wire \w[48][27] ;
 wire \w[48][28] ;
 wire \w[48][29] ;
 wire \w[48][2] ;
 wire \w[48][30] ;
 wire \w[48][31] ;
 wire \w[48][3] ;
 wire \w[48][4] ;
 wire \w[48][5] ;
 wire \w[48][6] ;
 wire \w[48][7] ;
 wire \w[48][8] ;
 wire \w[48][9] ;
 wire \w[49][0] ;
 wire \w[49][10] ;
 wire \w[49][11] ;
 wire \w[49][12] ;
 wire \w[49][13] ;
 wire \w[49][14] ;
 wire \w[49][15] ;
 wire \w[49][16] ;
 wire \w[49][17] ;
 wire \w[49][18] ;
 wire \w[49][19] ;
 wire \w[49][1] ;
 wire \w[49][20] ;
 wire \w[49][21] ;
 wire \w[49][22] ;
 wire \w[49][23] ;
 wire \w[49][24] ;
 wire \w[49][25] ;
 wire \w[49][26] ;
 wire \w[49][27] ;
 wire \w[49][28] ;
 wire \w[49][29] ;
 wire \w[49][2] ;
 wire \w[49][30] ;
 wire \w[49][31] ;
 wire \w[49][3] ;
 wire \w[49][4] ;
 wire \w[49][5] ;
 wire \w[49][6] ;
 wire \w[49][7] ;
 wire \w[49][8] ;
 wire \w[49][9] ;
 wire \w[4][0] ;
 wire \w[4][10] ;
 wire \w[4][11] ;
 wire \w[4][12] ;
 wire \w[4][13] ;
 wire \w[4][14] ;
 wire \w[4][15] ;
 wire \w[4][16] ;
 wire \w[4][17] ;
 wire \w[4][18] ;
 wire \w[4][19] ;
 wire \w[4][1] ;
 wire \w[4][20] ;
 wire \w[4][21] ;
 wire \w[4][22] ;
 wire \w[4][23] ;
 wire \w[4][24] ;
 wire \w[4][25] ;
 wire \w[4][26] ;
 wire \w[4][27] ;
 wire \w[4][28] ;
 wire \w[4][29] ;
 wire \w[4][2] ;
 wire \w[4][30] ;
 wire \w[4][31] ;
 wire \w[4][3] ;
 wire \w[4][4] ;
 wire \w[4][5] ;
 wire \w[4][6] ;
 wire \w[4][7] ;
 wire \w[4][8] ;
 wire \w[4][9] ;
 wire \w[50][0] ;
 wire \w[50][10] ;
 wire \w[50][11] ;
 wire \w[50][12] ;
 wire \w[50][13] ;
 wire \w[50][14] ;
 wire \w[50][15] ;
 wire \w[50][16] ;
 wire \w[50][17] ;
 wire \w[50][18] ;
 wire \w[50][19] ;
 wire \w[50][1] ;
 wire \w[50][20] ;
 wire \w[50][21] ;
 wire \w[50][22] ;
 wire \w[50][23] ;
 wire \w[50][24] ;
 wire \w[50][25] ;
 wire \w[50][26] ;
 wire \w[50][27] ;
 wire \w[50][28] ;
 wire \w[50][29] ;
 wire \w[50][2] ;
 wire \w[50][30] ;
 wire \w[50][31] ;
 wire \w[50][3] ;
 wire \w[50][4] ;
 wire \w[50][5] ;
 wire \w[50][6] ;
 wire \w[50][7] ;
 wire \w[50][8] ;
 wire \w[50][9] ;
 wire \w[51][0] ;
 wire \w[51][10] ;
 wire \w[51][11] ;
 wire \w[51][12] ;
 wire \w[51][13] ;
 wire \w[51][14] ;
 wire \w[51][15] ;
 wire \w[51][16] ;
 wire \w[51][17] ;
 wire \w[51][18] ;
 wire \w[51][19] ;
 wire \w[51][1] ;
 wire \w[51][20] ;
 wire \w[51][21] ;
 wire \w[51][22] ;
 wire \w[51][23] ;
 wire \w[51][24] ;
 wire \w[51][25] ;
 wire \w[51][26] ;
 wire \w[51][27] ;
 wire \w[51][28] ;
 wire \w[51][29] ;
 wire \w[51][2] ;
 wire \w[51][30] ;
 wire \w[51][31] ;
 wire \w[51][3] ;
 wire \w[51][4] ;
 wire \w[51][5] ;
 wire \w[51][6] ;
 wire \w[51][7] ;
 wire \w[51][8] ;
 wire \w[51][9] ;
 wire \w[52][0] ;
 wire \w[52][10] ;
 wire \w[52][11] ;
 wire \w[52][12] ;
 wire \w[52][13] ;
 wire \w[52][14] ;
 wire \w[52][15] ;
 wire \w[52][16] ;
 wire \w[52][17] ;
 wire \w[52][18] ;
 wire \w[52][19] ;
 wire \w[52][1] ;
 wire \w[52][20] ;
 wire \w[52][21] ;
 wire \w[52][22] ;
 wire \w[52][23] ;
 wire \w[52][24] ;
 wire \w[52][25] ;
 wire \w[52][26] ;
 wire \w[52][27] ;
 wire \w[52][28] ;
 wire \w[52][29] ;
 wire \w[52][2] ;
 wire \w[52][30] ;
 wire \w[52][31] ;
 wire \w[52][3] ;
 wire \w[52][4] ;
 wire \w[52][5] ;
 wire \w[52][6] ;
 wire \w[52][7] ;
 wire \w[52][8] ;
 wire \w[52][9] ;
 wire \w[53][0] ;
 wire \w[53][10] ;
 wire \w[53][11] ;
 wire \w[53][12] ;
 wire \w[53][13] ;
 wire \w[53][14] ;
 wire \w[53][15] ;
 wire \w[53][16] ;
 wire \w[53][17] ;
 wire \w[53][18] ;
 wire \w[53][19] ;
 wire \w[53][1] ;
 wire \w[53][20] ;
 wire \w[53][21] ;
 wire \w[53][22] ;
 wire \w[53][23] ;
 wire \w[53][24] ;
 wire \w[53][25] ;
 wire \w[53][26] ;
 wire \w[53][27] ;
 wire \w[53][28] ;
 wire \w[53][29] ;
 wire \w[53][2] ;
 wire \w[53][30] ;
 wire \w[53][31] ;
 wire \w[53][3] ;
 wire \w[53][4] ;
 wire \w[53][5] ;
 wire \w[53][6] ;
 wire \w[53][7] ;
 wire \w[53][8] ;
 wire \w[53][9] ;
 wire \w[54][0] ;
 wire \w[54][10] ;
 wire \w[54][11] ;
 wire \w[54][12] ;
 wire \w[54][13] ;
 wire \w[54][14] ;
 wire \w[54][15] ;
 wire \w[54][16] ;
 wire \w[54][17] ;
 wire \w[54][18] ;
 wire \w[54][19] ;
 wire \w[54][1] ;
 wire \w[54][20] ;
 wire \w[54][21] ;
 wire \w[54][22] ;
 wire \w[54][23] ;
 wire \w[54][24] ;
 wire \w[54][25] ;
 wire \w[54][26] ;
 wire \w[54][27] ;
 wire \w[54][28] ;
 wire \w[54][29] ;
 wire \w[54][2] ;
 wire \w[54][30] ;
 wire \w[54][31] ;
 wire \w[54][3] ;
 wire \w[54][4] ;
 wire \w[54][5] ;
 wire \w[54][6] ;
 wire \w[54][7] ;
 wire \w[54][8] ;
 wire \w[54][9] ;
 wire \w[55][0] ;
 wire \w[55][10] ;
 wire \w[55][11] ;
 wire \w[55][12] ;
 wire \w[55][13] ;
 wire \w[55][14] ;
 wire \w[55][15] ;
 wire \w[55][16] ;
 wire \w[55][17] ;
 wire \w[55][18] ;
 wire \w[55][19] ;
 wire \w[55][1] ;
 wire \w[55][20] ;
 wire \w[55][21] ;
 wire \w[55][22] ;
 wire \w[55][23] ;
 wire \w[55][24] ;
 wire \w[55][25] ;
 wire \w[55][26] ;
 wire \w[55][27] ;
 wire \w[55][28] ;
 wire \w[55][29] ;
 wire \w[55][2] ;
 wire \w[55][30] ;
 wire \w[55][31] ;
 wire \w[55][3] ;
 wire \w[55][4] ;
 wire \w[55][5] ;
 wire \w[55][6] ;
 wire \w[55][7] ;
 wire \w[55][8] ;
 wire \w[55][9] ;
 wire \w[56][0] ;
 wire \w[56][10] ;
 wire \w[56][11] ;
 wire \w[56][12] ;
 wire \w[56][13] ;
 wire \w[56][14] ;
 wire \w[56][15] ;
 wire \w[56][16] ;
 wire \w[56][17] ;
 wire \w[56][18] ;
 wire \w[56][19] ;
 wire \w[56][1] ;
 wire \w[56][20] ;
 wire \w[56][21] ;
 wire \w[56][22] ;
 wire \w[56][23] ;
 wire \w[56][24] ;
 wire \w[56][25] ;
 wire \w[56][26] ;
 wire \w[56][27] ;
 wire \w[56][28] ;
 wire \w[56][29] ;
 wire \w[56][2] ;
 wire \w[56][30] ;
 wire \w[56][31] ;
 wire \w[56][3] ;
 wire \w[56][4] ;
 wire \w[56][5] ;
 wire \w[56][6] ;
 wire \w[56][7] ;
 wire \w[56][8] ;
 wire \w[56][9] ;
 wire \w[57][0] ;
 wire \w[57][10] ;
 wire \w[57][11] ;
 wire \w[57][12] ;
 wire \w[57][13] ;
 wire \w[57][14] ;
 wire \w[57][15] ;
 wire \w[57][16] ;
 wire \w[57][17] ;
 wire \w[57][18] ;
 wire \w[57][19] ;
 wire \w[57][1] ;
 wire \w[57][20] ;
 wire \w[57][21] ;
 wire \w[57][22] ;
 wire \w[57][23] ;
 wire \w[57][24] ;
 wire \w[57][25] ;
 wire \w[57][26] ;
 wire \w[57][27] ;
 wire \w[57][28] ;
 wire \w[57][29] ;
 wire \w[57][2] ;
 wire \w[57][30] ;
 wire \w[57][31] ;
 wire \w[57][3] ;
 wire \w[57][4] ;
 wire \w[57][5] ;
 wire \w[57][6] ;
 wire \w[57][7] ;
 wire \w[57][8] ;
 wire \w[57][9] ;
 wire \w[58][0] ;
 wire \w[58][10] ;
 wire \w[58][11] ;
 wire \w[58][12] ;
 wire \w[58][13] ;
 wire \w[58][14] ;
 wire \w[58][15] ;
 wire \w[58][16] ;
 wire \w[58][17] ;
 wire \w[58][18] ;
 wire \w[58][19] ;
 wire \w[58][1] ;
 wire \w[58][20] ;
 wire \w[58][21] ;
 wire \w[58][22] ;
 wire \w[58][23] ;
 wire \w[58][24] ;
 wire \w[58][25] ;
 wire \w[58][26] ;
 wire \w[58][27] ;
 wire \w[58][28] ;
 wire \w[58][29] ;
 wire \w[58][2] ;
 wire \w[58][30] ;
 wire \w[58][31] ;
 wire \w[58][3] ;
 wire \w[58][4] ;
 wire \w[58][5] ;
 wire \w[58][6] ;
 wire \w[58][7] ;
 wire \w[58][8] ;
 wire \w[58][9] ;
 wire \w[59][0] ;
 wire \w[59][10] ;
 wire \w[59][11] ;
 wire \w[59][12] ;
 wire \w[59][13] ;
 wire \w[59][14] ;
 wire \w[59][15] ;
 wire \w[59][16] ;
 wire \w[59][17] ;
 wire \w[59][18] ;
 wire \w[59][19] ;
 wire \w[59][1] ;
 wire \w[59][20] ;
 wire \w[59][21] ;
 wire \w[59][22] ;
 wire \w[59][23] ;
 wire \w[59][24] ;
 wire \w[59][25] ;
 wire \w[59][26] ;
 wire \w[59][27] ;
 wire \w[59][28] ;
 wire \w[59][29] ;
 wire \w[59][2] ;
 wire \w[59][30] ;
 wire \w[59][31] ;
 wire \w[59][3] ;
 wire \w[59][4] ;
 wire \w[59][5] ;
 wire \w[59][6] ;
 wire \w[59][7] ;
 wire \w[59][8] ;
 wire \w[59][9] ;
 wire \w[5][0] ;
 wire \w[5][10] ;
 wire \w[5][11] ;
 wire \w[5][12] ;
 wire \w[5][13] ;
 wire \w[5][14] ;
 wire \w[5][15] ;
 wire \w[5][16] ;
 wire \w[5][17] ;
 wire \w[5][18] ;
 wire \w[5][19] ;
 wire \w[5][1] ;
 wire \w[5][20] ;
 wire \w[5][21] ;
 wire \w[5][22] ;
 wire \w[5][23] ;
 wire \w[5][24] ;
 wire \w[5][25] ;
 wire \w[5][26] ;
 wire \w[5][27] ;
 wire \w[5][28] ;
 wire \w[5][29] ;
 wire \w[5][2] ;
 wire \w[5][30] ;
 wire \w[5][31] ;
 wire \w[5][3] ;
 wire \w[5][4] ;
 wire \w[5][5] ;
 wire \w[5][6] ;
 wire \w[5][7] ;
 wire \w[5][8] ;
 wire \w[5][9] ;
 wire \w[60][0] ;
 wire \w[60][10] ;
 wire \w[60][11] ;
 wire \w[60][12] ;
 wire \w[60][13] ;
 wire \w[60][14] ;
 wire \w[60][15] ;
 wire \w[60][16] ;
 wire \w[60][17] ;
 wire \w[60][18] ;
 wire \w[60][19] ;
 wire \w[60][1] ;
 wire \w[60][20] ;
 wire \w[60][21] ;
 wire \w[60][22] ;
 wire \w[60][23] ;
 wire \w[60][24] ;
 wire \w[60][25] ;
 wire \w[60][26] ;
 wire \w[60][27] ;
 wire \w[60][28] ;
 wire \w[60][29] ;
 wire \w[60][2] ;
 wire \w[60][30] ;
 wire \w[60][31] ;
 wire \w[60][3] ;
 wire \w[60][4] ;
 wire \w[60][5] ;
 wire \w[60][6] ;
 wire \w[60][7] ;
 wire \w[60][8] ;
 wire \w[60][9] ;
 wire \w[61][0] ;
 wire \w[61][10] ;
 wire \w[61][11] ;
 wire \w[61][12] ;
 wire \w[61][13] ;
 wire \w[61][14] ;
 wire \w[61][15] ;
 wire \w[61][16] ;
 wire \w[61][17] ;
 wire \w[61][18] ;
 wire \w[61][19] ;
 wire \w[61][1] ;
 wire \w[61][20] ;
 wire \w[61][21] ;
 wire \w[61][22] ;
 wire \w[61][23] ;
 wire \w[61][24] ;
 wire \w[61][25] ;
 wire \w[61][26] ;
 wire \w[61][27] ;
 wire \w[61][28] ;
 wire \w[61][29] ;
 wire \w[61][2] ;
 wire \w[61][30] ;
 wire \w[61][31] ;
 wire \w[61][3] ;
 wire \w[61][4] ;
 wire \w[61][5] ;
 wire \w[61][6] ;
 wire \w[61][7] ;
 wire \w[61][8] ;
 wire \w[61][9] ;
 wire \w[62][0] ;
 wire \w[62][10] ;
 wire \w[62][11] ;
 wire \w[62][12] ;
 wire \w[62][13] ;
 wire \w[62][14] ;
 wire \w[62][15] ;
 wire \w[62][16] ;
 wire \w[62][17] ;
 wire \w[62][18] ;
 wire \w[62][19] ;
 wire \w[62][1] ;
 wire \w[62][20] ;
 wire \w[62][21] ;
 wire \w[62][22] ;
 wire \w[62][23] ;
 wire \w[62][24] ;
 wire \w[62][25] ;
 wire \w[62][26] ;
 wire \w[62][27] ;
 wire \w[62][28] ;
 wire \w[62][29] ;
 wire \w[62][2] ;
 wire \w[62][30] ;
 wire \w[62][31] ;
 wire \w[62][3] ;
 wire \w[62][4] ;
 wire \w[62][5] ;
 wire \w[62][6] ;
 wire \w[62][7] ;
 wire \w[62][8] ;
 wire \w[62][9] ;
 wire \w[63][0] ;
 wire \w[63][10] ;
 wire \w[63][11] ;
 wire \w[63][12] ;
 wire \w[63][13] ;
 wire \w[63][14] ;
 wire \w[63][15] ;
 wire \w[63][16] ;
 wire \w[63][17] ;
 wire \w[63][18] ;
 wire \w[63][19] ;
 wire \w[63][1] ;
 wire \w[63][20] ;
 wire \w[63][21] ;
 wire \w[63][22] ;
 wire \w[63][23] ;
 wire \w[63][24] ;
 wire \w[63][25] ;
 wire \w[63][26] ;
 wire \w[63][27] ;
 wire \w[63][28] ;
 wire \w[63][29] ;
 wire \w[63][2] ;
 wire \w[63][30] ;
 wire \w[63][31] ;
 wire \w[63][3] ;
 wire \w[63][4] ;
 wire \w[63][5] ;
 wire \w[63][6] ;
 wire \w[63][7] ;
 wire \w[63][8] ;
 wire \w[63][9] ;
 wire \w[6][0] ;
 wire \w[6][10] ;
 wire \w[6][11] ;
 wire \w[6][12] ;
 wire \w[6][13] ;
 wire \w[6][14] ;
 wire \w[6][15] ;
 wire \w[6][16] ;
 wire \w[6][17] ;
 wire \w[6][18] ;
 wire \w[6][19] ;
 wire \w[6][1] ;
 wire \w[6][20] ;
 wire \w[6][21] ;
 wire \w[6][22] ;
 wire \w[6][23] ;
 wire \w[6][24] ;
 wire \w[6][25] ;
 wire \w[6][26] ;
 wire \w[6][27] ;
 wire \w[6][28] ;
 wire \w[6][29] ;
 wire \w[6][2] ;
 wire \w[6][30] ;
 wire \w[6][31] ;
 wire \w[6][3] ;
 wire \w[6][4] ;
 wire \w[6][5] ;
 wire \w[6][6] ;
 wire \w[6][7] ;
 wire \w[6][8] ;
 wire \w[6][9] ;
 wire \w[7][0] ;
 wire \w[7][10] ;
 wire \w[7][11] ;
 wire \w[7][12] ;
 wire \w[7][13] ;
 wire \w[7][14] ;
 wire \w[7][15] ;
 wire \w[7][16] ;
 wire \w[7][17] ;
 wire \w[7][18] ;
 wire \w[7][19] ;
 wire \w[7][1] ;
 wire \w[7][20] ;
 wire \w[7][21] ;
 wire \w[7][22] ;
 wire \w[7][23] ;
 wire \w[7][24] ;
 wire \w[7][25] ;
 wire \w[7][26] ;
 wire \w[7][27] ;
 wire \w[7][28] ;
 wire \w[7][29] ;
 wire \w[7][2] ;
 wire \w[7][30] ;
 wire \w[7][31] ;
 wire \w[7][3] ;
 wire \w[7][4] ;
 wire \w[7][5] ;
 wire \w[7][6] ;
 wire \w[7][7] ;
 wire \w[7][8] ;
 wire \w[7][9] ;
 wire \w[8][0] ;
 wire \w[8][10] ;
 wire \w[8][11] ;
 wire \w[8][12] ;
 wire \w[8][13] ;
 wire \w[8][14] ;
 wire \w[8][15] ;
 wire \w[8][16] ;
 wire \w[8][17] ;
 wire \w[8][18] ;
 wire \w[8][19] ;
 wire \w[8][1] ;
 wire \w[8][20] ;
 wire \w[8][21] ;
 wire \w[8][22] ;
 wire \w[8][23] ;
 wire \w[8][24] ;
 wire \w[8][25] ;
 wire \w[8][26] ;
 wire \w[8][27] ;
 wire \w[8][28] ;
 wire \w[8][29] ;
 wire \w[8][2] ;
 wire \w[8][30] ;
 wire \w[8][31] ;
 wire \w[8][3] ;
 wire \w[8][4] ;
 wire \w[8][5] ;
 wire \w[8][6] ;
 wire \w[8][7] ;
 wire \w[8][8] ;
 wire \w[8][9] ;
 wire \w[9][0] ;
 wire \w[9][10] ;
 wire \w[9][11] ;
 wire \w[9][12] ;
 wire \w[9][13] ;
 wire \w[9][14] ;
 wire \w[9][15] ;
 wire \w[9][16] ;
 wire \w[9][17] ;
 wire \w[9][18] ;
 wire \w[9][19] ;
 wire \w[9][1] ;
 wire \w[9][20] ;
 wire \w[9][21] ;
 wire \w[9][22] ;
 wire \w[9][23] ;
 wire \w[9][24] ;
 wire \w[9][25] ;
 wire \w[9][26] ;
 wire \w[9][27] ;
 wire \w[9][28] ;
 wire \w[9][29] ;
 wire \w[9][2] ;
 wire \w[9][30] ;
 wire \w[9][31] ;
 wire \w[9][3] ;
 wire \w[9][4] ;
 wire \w[9][5] ;
 wire \w[9][6] ;
 wire \w[9][7] ;
 wire \w[9][8] ;
 wire \w[9][9] ;

 sky130_fd_sc_hd__mux4_2 _14209_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03883_));
 sky130_fd_sc_hd__mux4_2 _14210_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03884_));
 sky130_fd_sc_hd__mux4_2 _14211_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03885_));
 sky130_fd_sc_hd__mux4_2 _14212_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03886_));
 sky130_fd_sc_hd__mux4_2 _14213_ (.A0(_03883_),
    .A1(_03884_),
    .A2(_03885_),
    .A3(_03886_),
    .S0(net463),
    .S1(net459),
    .X(_03887_));
 sky130_fd_sc_hd__mux2i_4 _14214_ (.A0(_03882_),
    .A1(_03887_),
    .S(net458),
    .Y(_11944_));
 sky130_fd_sc_hd__mux4_2 _14215_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net426),
    .S1(net431),
    .X(_03888_));
 sky130_fd_sc_hd__mux4_2 _14216_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net426),
    .S1(net431),
    .X(_03889_));
 sky130_fd_sc_hd__mux4_2 _14217_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net426),
    .S1(net431),
    .X(_03890_));
 sky130_fd_sc_hd__mux4_2 _14218_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net426),
    .S1(net431),
    .X(_03891_));
 sky130_fd_sc_hd__mux4_2 _14219_ (.A0(_03888_),
    .A1(_03889_),
    .A2(_03890_),
    .A3(_03891_),
    .S0(net423),
    .S1(net421),
    .X(_03892_));
 sky130_fd_sc_hd__mux4_2 _14220_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net429),
    .S1(net432),
    .X(_03893_));
 sky130_fd_sc_hd__mux4_2 _14221_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net427),
    .S1(net432),
    .X(_03894_));
 sky130_fd_sc_hd__mux4_2 _14222_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net427),
    .S1(net432),
    .X(_03895_));
 sky130_fd_sc_hd__mux4_2 _14223_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net429),
    .S1(net432),
    .X(_03896_));
 sky130_fd_sc_hd__mux4_2 _14224_ (.A0(_03893_),
    .A1(_03894_),
    .A2(_03895_),
    .A3(_03896_),
    .S0(net422),
    .S1(net420),
    .X(_03897_));
 sky130_fd_sc_hd__mux2i_4 _14225_ (.A0(_03892_),
    .A1(_03897_),
    .S(net419),
    .Y(_03898_));
 sky130_fd_sc_hd__xnor2_1 _14226_ (.A(_03803_),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__xnor2_1 _14227_ (.A(_03389_),
    .B(_03899_),
    .Y(_11949_));
 sky130_fd_sc_hd__mux4_2 _14228_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net508),
    .S1(net513),
    .X(_03900_));
 sky130_fd_sc_hd__mux4_2 _14229_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net508),
    .S1(net513),
    .X(_03901_));
 sky130_fd_sc_hd__mux4_2 _14230_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net508),
    .S1(net513),
    .X(_03902_));
 sky130_fd_sc_hd__mux4_2 _14231_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net508),
    .S1(net513),
    .X(_03903_));
 sky130_fd_sc_hd__mux4_2 _14232_ (.A0(_03900_),
    .A1(_03901_),
    .A2(_03902_),
    .A3(_03903_),
    .S0(net502),
    .S1(net499),
    .X(_03904_));
 sky130_fd_sc_hd__mux4_2 _14233_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net509),
    .S1(net514),
    .X(_03905_));
 sky130_fd_sc_hd__mux4_2 _14234_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net509),
    .S1(net514),
    .X(_03906_));
 sky130_fd_sc_hd__mux4_2 _14235_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net509),
    .S1(net514),
    .X(_03907_));
 sky130_fd_sc_hd__mux4_2 _14236_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net509),
    .S1(net514),
    .X(_03908_));
 sky130_fd_sc_hd__mux4_2 _14237_ (.A0(_03905_),
    .A1(_03906_),
    .A2(_03907_),
    .A3(_03908_),
    .S0(net503),
    .S1(net500),
    .X(_03909_));
 sky130_fd_sc_hd__mux2i_4 _14238_ (.A0(_03904_),
    .A1(_03909_),
    .S(net497),
    .Y(_03910_));
 sky130_fd_sc_hd__xnor2_1 _14239_ (.A(_03264_),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__xnor2_2 _14240_ (.A(_02853_),
    .B(_03911_),
    .Y(_11948_));
 sky130_fd_sc_hd__mux4_2 _14241_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03912_));
 sky130_fd_sc_hd__mux4_2 _14242_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1464 ();
 sky130_fd_sc_hd__mux4_2 _14244_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03915_));
 sky130_fd_sc_hd__mux4_2 _14245_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03916_));
 sky130_fd_sc_hd__mux4_2 _14246_ (.A0(_03912_),
    .A1(_03913_),
    .A2(_03915_),
    .A3(_03916_),
    .S0(net386),
    .S1(net383),
    .X(_03917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1463 ();
 sky130_fd_sc_hd__mux4_2 _14248_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03919_));
 sky130_fd_sc_hd__mux4_2 _14249_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03920_));
 sky130_fd_sc_hd__mux4_2 _14250_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03921_));
 sky130_fd_sc_hd__mux4_2 _14251_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net389),
    .S1(net394),
    .X(_03922_));
 sky130_fd_sc_hd__mux4_2 _14252_ (.A0(_03919_),
    .A1(_03920_),
    .A2(_03921_),
    .A3(_03922_),
    .S0(net386),
    .S1(net383),
    .X(_03923_));
 sky130_fd_sc_hd__mux2i_4 _14253_ (.A0(_03917_),
    .A1(_03923_),
    .S(net381),
    .Y(_11947_));
 sky130_fd_sc_hd__mux4_2 _14254_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net471),
    .S1(net553),
    .X(_03924_));
 sky130_fd_sc_hd__mux4_2 _14255_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03925_));
 sky130_fd_sc_hd__mux4_2 _14256_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net471),
    .S1(net553),
    .X(_03926_));
 sky130_fd_sc_hd__mux4_2 _14257_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net471),
    .S1(net553),
    .X(_03927_));
 sky130_fd_sc_hd__mux4_2 _14258_ (.A0(_03924_),
    .A1(_03925_),
    .A2(_03926_),
    .A3(_03927_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_03928_));
 sky130_fd_sc_hd__mux4_2 _14259_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net471),
    .S1(net473),
    .X(_03929_));
 sky130_fd_sc_hd__mux4_2 _14260_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net471),
    .S1(\count16_2[1] ),
    .X(_03930_));
 sky130_fd_sc_hd__mux4_2 _14261_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net471),
    .S1(\count16_2[1] ),
    .X(_03931_));
 sky130_fd_sc_hd__mux4_2 _14262_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net471),
    .S1(\count16_2[1] ),
    .X(_03932_));
 sky130_fd_sc_hd__mux4_2 _14263_ (.A0(_03929_),
    .A1(_03930_),
    .A2(_03931_),
    .A3(_03932_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_03933_));
 sky130_fd_sc_hd__mux2i_4 _14264_ (.A0(_03928_),
    .A1(_03933_),
    .S(\count16_2[5] ),
    .Y(_11952_));
 sky130_fd_sc_hd__mux4_2 _14265_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03934_));
 sky130_fd_sc_hd__mux4_2 _14266_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03935_));
 sky130_fd_sc_hd__mux4_2 _14267_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03936_));
 sky130_fd_sc_hd__mux4_2 _14268_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03937_));
 sky130_fd_sc_hd__mux4_2 _14269_ (.A0(_03934_),
    .A1(_03935_),
    .A2(_03936_),
    .A3(_03937_),
    .S0(net549),
    .S1(net421),
    .X(_03938_));
 sky130_fd_sc_hd__mux4_2 _14270_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03939_));
 sky130_fd_sc_hd__mux4_2 _14271_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03940_));
 sky130_fd_sc_hd__mux4_2 _14272_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03941_));
 sky130_fd_sc_hd__mux4_2 _14273_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net424),
    .S1(net435),
    .X(_03942_));
 sky130_fd_sc_hd__mux4_2 _14274_ (.A0(_03939_),
    .A1(_03940_),
    .A2(_03941_),
    .A3(_03942_),
    .S0(net549),
    .S1(net548),
    .X(_03943_));
 sky130_fd_sc_hd__mux2i_4 _14275_ (.A0(_03938_),
    .A1(_03943_),
    .S(\count2_2[5] ),
    .Y(_03944_));
 sky130_fd_sc_hd__xnor2_1 _14276_ (.A(_03849_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__xnor2_1 _14277_ (.A(_03448_),
    .B(_03945_),
    .Y(_11957_));
 sky130_fd_sc_hd__mux4_2 _14278_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net505),
    .S1(net517),
    .X(_03946_));
 sky130_fd_sc_hd__mux4_2 _14279_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net505),
    .S1(net517),
    .X(_03947_));
 sky130_fd_sc_hd__mux4_2 _14280_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net505),
    .S1(net517),
    .X(_03948_));
 sky130_fd_sc_hd__mux4_2 _14281_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net505),
    .S1(net517),
    .X(_03949_));
 sky130_fd_sc_hd__mux4_2 _14282_ (.A0(_03946_),
    .A1(_03947_),
    .A2(_03948_),
    .A3(_03949_),
    .S0(net504),
    .S1(net501),
    .X(_03950_));
 sky130_fd_sc_hd__mux4_2 _14283_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03951_));
 sky130_fd_sc_hd__mux4_2 _14284_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03952_));
 sky130_fd_sc_hd__mux4_2 _14285_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03953_));
 sky130_fd_sc_hd__mux4_2 _14286_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03954_));
 sky130_fd_sc_hd__mux4_2 _14287_ (.A0(_03951_),
    .A1(_03952_),
    .A2(_03953_),
    .A3(_03954_),
    .S0(net504),
    .S1(net501),
    .X(_03955_));
 sky130_fd_sc_hd__mux2i_4 _14288_ (.A0(_03950_),
    .A1(_03955_),
    .S(\count15_2[5] ),
    .Y(_03956_));
 sky130_fd_sc_hd__xnor2_1 _14289_ (.A(_03333_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__xnor2_1 _14290_ (.A(net1140),
    .B(_03957_),
    .Y(_11956_));
 sky130_fd_sc_hd__mux4_2 _14291_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net389),
    .S1(net394),
    .X(_03958_));
 sky130_fd_sc_hd__mux4_2 _14292_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net393),
    .S1(net394),
    .X(_03959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1462 ();
 sky130_fd_sc_hd__mux4_2 _14294_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net393),
    .S1(net394),
    .X(_03961_));
 sky130_fd_sc_hd__mux4_2 _14295_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net393),
    .S1(net394),
    .X(_03962_));
 sky130_fd_sc_hd__mux4_2 _14296_ (.A0(_03958_),
    .A1(_03959_),
    .A2(_03961_),
    .A3(_03962_),
    .S0(net386),
    .S1(net383),
    .X(_03963_));
 sky130_fd_sc_hd__mux4_2 _14297_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net393),
    .S1(net544),
    .X(_03964_));
 sky130_fd_sc_hd__mux4_2 _14298_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net393),
    .S1(net544),
    .X(_03965_));
 sky130_fd_sc_hd__mux4_2 _14299_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net393),
    .S1(net544),
    .X(_03966_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1461 ();
 sky130_fd_sc_hd__mux4_2 _14301_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net393),
    .S1(net544),
    .X(_03968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1460 ();
 sky130_fd_sc_hd__mux4_2 _14303_ (.A0(_03964_),
    .A1(_03965_),
    .A2(_03966_),
    .A3(_03968_),
    .S0(net385),
    .S1(\count7_2[4] ),
    .X(_03970_));
 sky130_fd_sc_hd__mux2i_4 _14304_ (.A0(_03963_),
    .A1(_03970_),
    .S(net381),
    .Y(_11955_));
 sky130_fd_sc_hd__mux4_2 _14305_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net465),
    .S1(net476),
    .X(_03971_));
 sky130_fd_sc_hd__mux4_2 _14306_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net465),
    .S1(net476),
    .X(_03972_));
 sky130_fd_sc_hd__mux4_2 _14307_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net465),
    .S1(net476),
    .X(_03973_));
 sky130_fd_sc_hd__mux4_2 _14308_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net465),
    .S1(net476),
    .X(_03974_));
 sky130_fd_sc_hd__mux4_2 _14309_ (.A0(_03971_),
    .A1(_03972_),
    .A2(_03973_),
    .A3(_03974_),
    .S0(net462),
    .S1(net460),
    .X(_03975_));
 sky130_fd_sc_hd__mux4_2 _14310_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net469),
    .S1(net473),
    .X(_03976_));
 sky130_fd_sc_hd__mux4_2 _14311_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net469),
    .S1(net473),
    .X(_03977_));
 sky130_fd_sc_hd__mux4_2 _14312_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net469),
    .S1(net473),
    .X(_03978_));
 sky130_fd_sc_hd__mux4_2 _14313_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net469),
    .S1(net473),
    .X(_03979_));
 sky130_fd_sc_hd__mux4_2 _14314_ (.A0(_03976_),
    .A1(_03977_),
    .A2(_03978_),
    .A3(_03979_),
    .S0(net463),
    .S1(net459),
    .X(_03980_));
 sky130_fd_sc_hd__mux2i_4 _14315_ (.A0(_03975_),
    .A1(_03980_),
    .S(net457),
    .Y(_11960_));
 sky130_fd_sc_hd__mux4_2 _14316_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net426),
    .S1(net431),
    .X(_03981_));
 sky130_fd_sc_hd__mux4_2 _14317_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net426),
    .S1(net431),
    .X(_03982_));
 sky130_fd_sc_hd__mux4_2 _14318_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net426),
    .S1(net431),
    .X(_03983_));
 sky130_fd_sc_hd__mux4_2 _14319_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net426),
    .S1(net431),
    .X(_03984_));
 sky130_fd_sc_hd__mux4_2 _14320_ (.A0(_03981_),
    .A1(_03982_),
    .A2(_03983_),
    .A3(_03984_),
    .S0(net423),
    .S1(net421),
    .X(_03985_));
 sky130_fd_sc_hd__mux4_2 _14321_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net429),
    .S1(net432),
    .X(_03986_));
 sky130_fd_sc_hd__mux4_2 _14322_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net429),
    .S1(net432),
    .X(_03987_));
 sky130_fd_sc_hd__mux4_2 _14323_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net429),
    .S1(net432),
    .X(_03988_));
 sky130_fd_sc_hd__mux4_2 _14324_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net429),
    .S1(net432),
    .X(_03989_));
 sky130_fd_sc_hd__mux4_2 _14325_ (.A0(_03986_),
    .A1(_03987_),
    .A2(_03988_),
    .A3(_03989_),
    .S0(net422),
    .S1(net421),
    .X(_03990_));
 sky130_fd_sc_hd__mux2i_4 _14326_ (.A0(_03985_),
    .A1(_03990_),
    .S(net419),
    .Y(_03991_));
 sky130_fd_sc_hd__xnor2_1 _14327_ (.A(_03898_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__xnor2_1 _14328_ (.A(_03507_),
    .B(_03992_),
    .Y(_11965_));
 sky130_fd_sc_hd__xnor2_1 _14329_ (.A(_03109_),
    .B(_03413_),
    .Y(_03993_));
 sky130_fd_sc_hd__xnor2_1 _14330_ (.A(_02824_),
    .B(_03993_),
    .Y(_11964_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1459 ();
 sky130_fd_sc_hd__mux4_2 _14332_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net387),
    .S1(net544),
    .X(_03995_));
 sky130_fd_sc_hd__mux4_2 _14333_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net387),
    .S1(net544),
    .X(_03996_));
 sky130_fd_sc_hd__mux4_2 _14334_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net387),
    .S1(net544),
    .X(_03997_));
 sky130_fd_sc_hd__mux4_2 _14335_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net387),
    .S1(net544),
    .X(_03998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1458 ();
 sky130_fd_sc_hd__mux4_2 _14337_ (.A0(_03995_),
    .A1(_03996_),
    .A2(_03997_),
    .A3(_03998_),
    .S0(net385),
    .S1(net382),
    .X(_04000_));
 sky130_fd_sc_hd__mux4_2 _14338_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net387),
    .S1(net544),
    .X(_04001_));
 sky130_fd_sc_hd__mux4_2 _14339_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net387),
    .S1(net544),
    .X(_04002_));
 sky130_fd_sc_hd__mux4_2 _14340_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net387),
    .S1(net544),
    .X(_04003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1457 ();
 sky130_fd_sc_hd__mux4_2 _14342_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net388),
    .S1(net544),
    .X(_04005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1456 ();
 sky130_fd_sc_hd__mux4_2 _14344_ (.A0(_04001_),
    .A1(_04002_),
    .A2(_04003_),
    .A3(_04005_),
    .S0(net385),
    .S1(net382),
    .X(_04007_));
 sky130_fd_sc_hd__mux2i_4 _14345_ (.A0(_04000_),
    .A1(_04007_),
    .S(net381),
    .Y(_11963_));
 sky130_fd_sc_hd__mux4_2 _14346_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net467),
    .S1(net475),
    .X(_04008_));
 sky130_fd_sc_hd__mux4_2 _14347_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net467),
    .S1(net475),
    .X(_04009_));
 sky130_fd_sc_hd__mux4_2 _14348_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net467),
    .S1(net475),
    .X(_04010_));
 sky130_fd_sc_hd__mux4_2 _14349_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net467),
    .S1(net475),
    .X(_04011_));
 sky130_fd_sc_hd__mux4_2 _14350_ (.A0(_04008_),
    .A1(_04009_),
    .A2(_04010_),
    .A3(_04011_),
    .S0(net462),
    .S1(net460),
    .X(_04012_));
 sky130_fd_sc_hd__mux4_2 _14351_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net467),
    .S1(net476),
    .X(_04013_));
 sky130_fd_sc_hd__mux4_2 _14352_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net467),
    .S1(net476),
    .X(_04014_));
 sky130_fd_sc_hd__mux4_2 _14353_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net467),
    .S1(net476),
    .X(_04015_));
 sky130_fd_sc_hd__mux4_2 _14354_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net467),
    .S1(net476),
    .X(_04016_));
 sky130_fd_sc_hd__mux4_2 _14355_ (.A0(_04013_),
    .A1(_04014_),
    .A2(_04015_),
    .A3(_04016_),
    .S0(net462),
    .S1(net460),
    .X(_04017_));
 sky130_fd_sc_hd__mux2i_4 _14356_ (.A0(_04012_),
    .A1(_04017_),
    .S(net458),
    .Y(_11968_));
 sky130_fd_sc_hd__mux4_2 _14357_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04018_));
 sky130_fd_sc_hd__mux4_2 _14358_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04019_));
 sky130_fd_sc_hd__mux4_2 _14359_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04020_));
 sky130_fd_sc_hd__mux4_2 _14360_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04021_));
 sky130_fd_sc_hd__mux4_2 _14361_ (.A0(_04018_),
    .A1(_04019_),
    .A2(_04020_),
    .A3(_04021_),
    .S0(net549),
    .S1(net548),
    .X(_04022_));
 sky130_fd_sc_hd__mux4_2 _14362_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04023_));
 sky130_fd_sc_hd__mux4_2 _14363_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04024_));
 sky130_fd_sc_hd__mux4_2 _14364_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04025_));
 sky130_fd_sc_hd__mux4_2 _14365_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net424),
    .S1(net435),
    .X(_04026_));
 sky130_fd_sc_hd__mux4_2 _14366_ (.A0(_04023_),
    .A1(_04024_),
    .A2(_04025_),
    .A3(_04026_),
    .S0(net549),
    .S1(net548),
    .X(_04027_));
 sky130_fd_sc_hd__mux2i_4 _14367_ (.A0(_04022_),
    .A1(_04027_),
    .S(\count2_2[5] ),
    .Y(_04028_));
 sky130_fd_sc_hd__xnor2_1 _14368_ (.A(_03944_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__xnor2_1 _14369_ (.A(_03567_),
    .B(_04029_),
    .Y(_11973_));
 sky130_fd_sc_hd__xnor2_1 _14370_ (.A(_03181_),
    .B(_03471_),
    .Y(_04030_));
 sky130_fd_sc_hd__xnor2_1 _14371_ (.A(_02976_),
    .B(_04030_),
    .Y(_11972_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1455 ();
 sky130_fd_sc_hd__mux4_2 _14373_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04032_));
 sky130_fd_sc_hd__mux4_2 _14374_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04033_));
 sky130_fd_sc_hd__mux4_2 _14375_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1454 ();
 sky130_fd_sc_hd__mux4_2 _14377_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1453 ();
 sky130_fd_sc_hd__mux4_2 _14379_ (.A0(_04032_),
    .A1(_04033_),
    .A2(_04034_),
    .A3(_04036_),
    .S0(net384),
    .S1(net542),
    .X(_04038_));
 sky130_fd_sc_hd__mux4_2 _14380_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04039_));
 sky130_fd_sc_hd__mux4_2 _14381_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04040_));
 sky130_fd_sc_hd__mux4_2 _14382_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04041_));
 sky130_fd_sc_hd__mux4_2 _14383_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net391),
    .S1(net397),
    .X(_04042_));
 sky130_fd_sc_hd__mux4_2 _14384_ (.A0(_04039_),
    .A1(_04040_),
    .A2(_04041_),
    .A3(_04042_),
    .S0(net384),
    .S1(net542),
    .X(_04043_));
 sky130_fd_sc_hd__mux2i_4 _14385_ (.A0(_04038_),
    .A1(_04043_),
    .S(net380),
    .Y(_11971_));
 sky130_fd_sc_hd__mux4_2 _14386_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net470),
    .S1(net474),
    .X(_04044_));
 sky130_fd_sc_hd__mux4_2 _14387_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net470),
    .S1(net474),
    .X(_04045_));
 sky130_fd_sc_hd__mux4_2 _14388_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net470),
    .S1(net474),
    .X(_04046_));
 sky130_fd_sc_hd__mux4_2 _14389_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net470),
    .S1(net474),
    .X(_04047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1452 ();
 sky130_fd_sc_hd__mux4_2 _14391_ (.A0(_04044_),
    .A1(_04045_),
    .A2(_04046_),
    .A3(_04047_),
    .S0(\count16_2[3] ),
    .S1(net459),
    .X(_04049_));
 sky130_fd_sc_hd__mux4_2 _14392_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net466),
    .S1(net474),
    .X(_04050_));
 sky130_fd_sc_hd__mux4_2 _14393_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net466),
    .S1(net474),
    .X(_04051_));
 sky130_fd_sc_hd__mux4_2 _14394_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net466),
    .S1(net474),
    .X(_04052_));
 sky130_fd_sc_hd__mux4_2 _14395_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net466),
    .S1(net474),
    .X(_04053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1451 ();
 sky130_fd_sc_hd__mux4_2 _14397_ (.A0(_04050_),
    .A1(_04051_),
    .A2(_04052_),
    .A3(_04053_),
    .S0(net463),
    .S1(net459),
    .X(_04055_));
 sky130_fd_sc_hd__mux2i_4 _14398_ (.A0(_04049_),
    .A1(_04055_),
    .S(net458),
    .Y(_11976_));
 sky130_fd_sc_hd__mux4_2 _14399_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_04056_));
 sky130_fd_sc_hd__mux4_2 _14400_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_04057_));
 sky130_fd_sc_hd__mux4_2 _14401_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_04058_));
 sky130_fd_sc_hd__mux4_2 _14402_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_04059_));
 sky130_fd_sc_hd__mux4_2 _14403_ (.A0(_04056_),
    .A1(_04057_),
    .A2(_04058_),
    .A3(_04059_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_04060_));
 sky130_fd_sc_hd__mux4_2 _14404_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(\count2_2[2] ),
    .S1(net433),
    .X(_04061_));
 sky130_fd_sc_hd__mux4_2 _14405_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(\count2_2[2] ),
    .S1(net433),
    .X(_04062_));
 sky130_fd_sc_hd__mux4_2 _14406_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_04063_));
 sky130_fd_sc_hd__mux4_2 _14407_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(\count2_2[2] ),
    .S1(net435),
    .X(_04064_));
 sky130_fd_sc_hd__mux4_2 _14408_ (.A0(_04061_),
    .A1(_04062_),
    .A2(_04063_),
    .A3(_04064_),
    .S0(net423),
    .S1(net548),
    .X(_04065_));
 sky130_fd_sc_hd__mux2i_4 _14409_ (.A0(_04060_),
    .A1(_04065_),
    .S(net419),
    .Y(_04066_));
 sky130_fd_sc_hd__xnor2_1 _14410_ (.A(_03991_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__xnor2_1 _14411_ (.A(_03633_),
    .B(_04067_),
    .Y(_11981_));
 sky130_fd_sc_hd__xnor2_1 _14412_ (.A(_03264_),
    .B(_03530_),
    .Y(_04068_));
 sky130_fd_sc_hd__xnor2_1 _14413_ (.A(_03098_),
    .B(_04068_),
    .Y(_11980_));
 sky130_fd_sc_hd__mux4_2 _14414_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net387),
    .S1(net396),
    .X(_04069_));
 sky130_fd_sc_hd__mux4_2 _14415_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net387),
    .S1(net396),
    .X(_04070_));
 sky130_fd_sc_hd__mux4_2 _14416_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net387),
    .S1(net396),
    .X(_04071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1450 ();
 sky130_fd_sc_hd__mux4_2 _14418_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net387),
    .S1(net396),
    .X(_04073_));
 sky130_fd_sc_hd__mux4_2 _14419_ (.A0(_04069_),
    .A1(_04070_),
    .A2(_04071_),
    .A3(_04073_),
    .S0(net385),
    .S1(net382),
    .X(_04074_));
 sky130_fd_sc_hd__mux4_2 _14420_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net390),
    .S1(net395),
    .X(_04075_));
 sky130_fd_sc_hd__mux4_2 _14421_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net392),
    .S1(net396),
    .X(_04076_));
 sky130_fd_sc_hd__mux4_2 _14422_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net392),
    .S1(net396),
    .X(_04077_));
 sky130_fd_sc_hd__mux4_2 _14423_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net392),
    .S1(net396),
    .X(_04078_));
 sky130_fd_sc_hd__mux4_2 _14424_ (.A0(_04075_),
    .A1(_04076_),
    .A2(_04077_),
    .A3(_04078_),
    .S0(net384),
    .S1(net542),
    .X(_04079_));
 sky130_fd_sc_hd__mux2i_4 _14425_ (.A0(_04074_),
    .A1(_04079_),
    .S(net380),
    .Y(_11979_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1449 ();
 sky130_fd_sc_hd__mux4_2 _14427_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net466),
    .S1(net474),
    .X(_04081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1448 ();
 sky130_fd_sc_hd__mux4_2 _14429_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net466),
    .S1(net474),
    .X(_04083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1447 ();
 sky130_fd_sc_hd__mux4_2 _14431_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net466),
    .S1(net474),
    .X(_04085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1446 ();
 sky130_fd_sc_hd__mux4_2 _14433_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net466),
    .S1(net474),
    .X(_04087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1445 ();
 sky130_fd_sc_hd__mux4_2 _14435_ (.A0(_04081_),
    .A1(_04083_),
    .A2(_04085_),
    .A3(_04087_),
    .S0(net462),
    .S1(net460),
    .X(_04089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1444 ();
 sky130_fd_sc_hd__mux4_2 _14437_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net469),
    .S1(net473),
    .X(_04091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1443 ();
 sky130_fd_sc_hd__mux4_2 _14439_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net469),
    .S1(net473),
    .X(_04093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1442 ();
 sky130_fd_sc_hd__mux4_2 _14441_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net469),
    .S1(net473),
    .X(_04095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1441 ();
 sky130_fd_sc_hd__mux4_2 _14443_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net469),
    .S1(net473),
    .X(_04097_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1440 ();
 sky130_fd_sc_hd__mux4_2 _14445_ (.A0(_04091_),
    .A1(_04093_),
    .A2(_04095_),
    .A3(_04097_),
    .S0(net463),
    .S1(net459),
    .X(_04099_));
 sky130_fd_sc_hd__mux2i_4 _14446_ (.A0(_04089_),
    .A1(_04099_),
    .S(net457),
    .Y(_11984_));
 sky130_fd_sc_hd__mux4_2 _14447_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net425),
    .S1(net436),
    .X(_04100_));
 sky130_fd_sc_hd__mux4_2 _14448_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net425),
    .S1(net436),
    .X(_04101_));
 sky130_fd_sc_hd__mux4_2 _14449_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net425),
    .S1(net436),
    .X(_04102_));
 sky130_fd_sc_hd__mux4_2 _14450_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net425),
    .S1(net436),
    .X(_04103_));
 sky130_fd_sc_hd__mux4_2 _14451_ (.A0(_04100_),
    .A1(_04101_),
    .A2(_04102_),
    .A3(_04103_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_04104_));
 sky130_fd_sc_hd__mux4_2 _14452_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net430),
    .S1(net433),
    .X(_04105_));
 sky130_fd_sc_hd__mux4_2 _14453_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net430),
    .S1(net433),
    .X(_04106_));
 sky130_fd_sc_hd__mux4_2 _14454_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net430),
    .S1(net433),
    .X(_04107_));
 sky130_fd_sc_hd__mux4_2 _14455_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net430),
    .S1(net433),
    .X(_04108_));
 sky130_fd_sc_hd__mux4_2 _14456_ (.A0(_04105_),
    .A1(_04106_),
    .A2(_04107_),
    .A3(_04108_),
    .S0(net423),
    .S1(\count2_2[4] ),
    .X(_04109_));
 sky130_fd_sc_hd__mux2i_4 _14457_ (.A0(_04104_),
    .A1(_04109_),
    .S(net419),
    .Y(_04110_));
 sky130_fd_sc_hd__xnor2_1 _14458_ (.A(_04028_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__xnor2_1 _14459_ (.A(_03697_),
    .B(_04111_),
    .Y(_11989_));
 sky130_fd_sc_hd__xnor2_1 _14460_ (.A(_03333_),
    .B(_03590_),
    .Y(_04112_));
 sky130_fd_sc_hd__xnor2_2 _14461_ (.A(_03194_),
    .B(_04112_),
    .Y(_11988_));
 sky130_fd_sc_hd__mux4_2 _14462_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net390),
    .S1(net395),
    .X(_04113_));
 sky130_fd_sc_hd__mux4_2 _14463_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net390),
    .S1(net395),
    .X(_04114_));
 sky130_fd_sc_hd__mux4_2 _14464_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net390),
    .S1(net395),
    .X(_04115_));
 sky130_fd_sc_hd__mux4_2 _14465_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net390),
    .S1(net395),
    .X(_04116_));
 sky130_fd_sc_hd__mux4_2 _14466_ (.A0(_04113_),
    .A1(_04114_),
    .A2(_04115_),
    .A3(_04116_),
    .S0(net384),
    .S1(net542),
    .X(_04117_));
 sky130_fd_sc_hd__mux4_2 _14467_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net391),
    .S1(net397),
    .X(_04118_));
 sky130_fd_sc_hd__mux4_2 _14468_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net391),
    .S1(net397),
    .X(_04119_));
 sky130_fd_sc_hd__mux4_2 _14469_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net391),
    .S1(net397),
    .X(_04120_));
 sky130_fd_sc_hd__mux4_2 _14470_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net391),
    .S1(net397),
    .X(_04121_));
 sky130_fd_sc_hd__mux4_2 _14471_ (.A0(_04118_),
    .A1(_04119_),
    .A2(_04120_),
    .A3(_04121_),
    .S0(net384),
    .S1(net542),
    .X(_04122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1439 ();
 sky130_fd_sc_hd__mux2i_4 _14473_ (.A0(_04117_),
    .A1(_04122_),
    .S(net380),
    .Y(_11987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1438 ();
 sky130_fd_sc_hd__mux4_2 _14475_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1437 ();
 sky130_fd_sc_hd__mux4_2 _14477_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1436 ();
 sky130_fd_sc_hd__mux4_2 _14479_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04129_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1435 ();
 sky130_fd_sc_hd__mux4_2 _14481_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04131_));
 sky130_fd_sc_hd__mux4_2 _14482_ (.A0(_04125_),
    .A1(_04127_),
    .A2(_04129_),
    .A3(_04131_),
    .S0(\count16_2[3] ),
    .S1(net461),
    .X(_04132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1434 ();
 sky130_fd_sc_hd__mux4_2 _14484_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1433 ();
 sky130_fd_sc_hd__mux4_2 _14486_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04136_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1432 ();
 sky130_fd_sc_hd__mux4_2 _14488_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1431 ();
 sky130_fd_sc_hd__mux4_2 _14490_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net472),
    .S1(net477),
    .X(_04140_));
 sky130_fd_sc_hd__mux4_2 _14491_ (.A0(_04134_),
    .A1(_04136_),
    .A2(_04138_),
    .A3(_04140_),
    .S0(\count16_2[3] ),
    .S1(net461),
    .X(_04141_));
 sky130_fd_sc_hd__mux2i_4 _14492_ (.A0(_04132_),
    .A1(_04141_),
    .S(net458),
    .Y(_11992_));
 sky130_fd_sc_hd__mux4_2 _14493_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net427),
    .S1(net432),
    .X(_04142_));
 sky130_fd_sc_hd__mux4_2 _14494_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net427),
    .S1(net432),
    .X(_04143_));
 sky130_fd_sc_hd__mux4_2 _14495_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net427),
    .S1(net432),
    .X(_04144_));
 sky130_fd_sc_hd__mux4_2 _14496_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net427),
    .S1(net432),
    .X(_04145_));
 sky130_fd_sc_hd__mux4_2 _14497_ (.A0(_04142_),
    .A1(_04143_),
    .A2(_04144_),
    .A3(_04145_),
    .S0(net423),
    .S1(net421),
    .X(_04146_));
 sky130_fd_sc_hd__mux4_2 _14498_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net429),
    .S1(net433),
    .X(_04147_));
 sky130_fd_sc_hd__mux4_2 _14499_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net429),
    .S1(net433),
    .X(_04148_));
 sky130_fd_sc_hd__mux4_2 _14500_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net429),
    .S1(net433),
    .X(_04149_));
 sky130_fd_sc_hd__mux4_2 _14501_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net429),
    .S1(net433),
    .X(_04150_));
 sky130_fd_sc_hd__mux4_2 _14502_ (.A0(_04147_),
    .A1(_04148_),
    .A2(_04149_),
    .A3(_04150_),
    .S0(net422),
    .S1(net420),
    .X(_04151_));
 sky130_fd_sc_hd__mux2i_2 _14503_ (.A0(_04146_),
    .A1(_04151_),
    .S(net418),
    .Y(_04152_));
 sky130_fd_sc_hd__xnor2_1 _14504_ (.A(_04066_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__xnor2_1 _14505_ (.A(_03743_),
    .B(_04153_),
    .Y(_11997_));
 sky130_fd_sc_hd__xnor2_1 _14506_ (.A(_03413_),
    .B(_03645_),
    .Y(_04154_));
 sky130_fd_sc_hd__xnor2_2 _14507_ (.A(_02882_),
    .B(_04154_),
    .Y(_11996_));
 sky130_fd_sc_hd__mux4_2 _14508_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net387),
    .S1(net398),
    .X(_04155_));
 sky130_fd_sc_hd__mux4_2 _14509_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net387),
    .S1(net398),
    .X(_04156_));
 sky130_fd_sc_hd__mux4_2 _14510_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net387),
    .S1(net398),
    .X(_04157_));
 sky130_fd_sc_hd__mux4_2 _14511_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net387),
    .S1(net398),
    .X(_04158_));
 sky130_fd_sc_hd__mux4_2 _14512_ (.A0(_04155_),
    .A1(_04156_),
    .A2(_04157_),
    .A3(_04158_),
    .S0(net385),
    .S1(net382),
    .X(_04159_));
 sky130_fd_sc_hd__mux4_2 _14513_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net392),
    .S1(net396),
    .X(_04160_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1430 ();
 sky130_fd_sc_hd__mux4_2 _14515_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net392),
    .S1(net396),
    .X(_04162_));
 sky130_fd_sc_hd__mux4_2 _14516_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net392),
    .S1(net396),
    .X(_04163_));
 sky130_fd_sc_hd__mux4_2 _14517_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net392),
    .S1(net396),
    .X(_04164_));
 sky130_fd_sc_hd__mux4_2 _14518_ (.A0(_04160_),
    .A1(_04162_),
    .A2(_04163_),
    .A3(_04164_),
    .S0(net385),
    .S1(net382),
    .X(_04165_));
 sky130_fd_sc_hd__mux2i_4 _14519_ (.A0(_04159_),
    .A1(_04165_),
    .S(net380),
    .Y(_11995_));
 sky130_fd_sc_hd__mux4_2 _14520_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04166_));
 sky130_fd_sc_hd__mux4_2 _14521_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04167_));
 sky130_fd_sc_hd__mux4_2 _14522_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04168_));
 sky130_fd_sc_hd__mux4_2 _14523_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04169_));
 sky130_fd_sc_hd__mux4_2 _14524_ (.A0(_04166_),
    .A1(_04167_),
    .A2(_04168_),
    .A3(_04169_),
    .S0(\count16_2[3] ),
    .S1(net459),
    .X(_04170_));
 sky130_fd_sc_hd__mux4_2 _14525_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04171_));
 sky130_fd_sc_hd__mux4_2 _14526_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04172_));
 sky130_fd_sc_hd__mux4_2 _14527_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04173_));
 sky130_fd_sc_hd__mux4_2 _14528_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net470),
    .S1(net473),
    .X(_04174_));
 sky130_fd_sc_hd__mux4_2 _14529_ (.A0(_04171_),
    .A1(_04172_),
    .A2(_04173_),
    .A3(_04174_),
    .S0(\count16_2[3] ),
    .S1(net459),
    .X(_04175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1429 ();
 sky130_fd_sc_hd__mux2i_4 _14531_ (.A0(_04170_),
    .A1(_04175_),
    .S(net457),
    .Y(_12000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1428 ();
 sky130_fd_sc_hd__mux4_2 _14533_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net430),
    .S1(net434),
    .X(_04178_));
 sky130_fd_sc_hd__mux4_2 _14534_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net430),
    .S1(net434),
    .X(_04179_));
 sky130_fd_sc_hd__mux4_2 _14535_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net430),
    .S1(net434),
    .X(_04180_));
 sky130_fd_sc_hd__mux4_2 _14536_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net430),
    .S1(net434),
    .X(_04181_));
 sky130_fd_sc_hd__mux4_2 _14537_ (.A0(_04178_),
    .A1(_04179_),
    .A2(_04180_),
    .A3(_04181_),
    .S0(net422),
    .S1(net420),
    .X(_04182_));
 sky130_fd_sc_hd__mux4_2 _14538_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net430),
    .S1(net434),
    .X(_04183_));
 sky130_fd_sc_hd__mux4_2 _14539_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net430),
    .S1(net434),
    .X(_04184_));
 sky130_fd_sc_hd__mux4_2 _14540_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net430),
    .S1(net434),
    .X(_04185_));
 sky130_fd_sc_hd__mux4_2 _14541_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_04186_));
 sky130_fd_sc_hd__mux4_2 _14542_ (.A0(_04183_),
    .A1(_04184_),
    .A2(_04185_),
    .A3(_04186_),
    .S0(net423),
    .S1(net420),
    .X(_04187_));
 sky130_fd_sc_hd__mux2i_4 _14543_ (.A0(_04182_),
    .A1(_04187_),
    .S(net418),
    .Y(_04188_));
 sky130_fd_sc_hd__xnor2_1 _14544_ (.A(_04110_),
    .B(_04188_),
    .Y(_12005_));
 sky130_fd_sc_hd__xnor2_1 _14545_ (.A(_03471_),
    .B(_03709_),
    .Y(_04189_));
 sky130_fd_sc_hd__xnor2_1 _14546_ (.A(net1133),
    .B(_04189_),
    .Y(_12004_));
 sky130_fd_sc_hd__mux4_2 _14547_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net390),
    .S1(net395),
    .X(_04190_));
 sky130_fd_sc_hd__mux4_2 _14548_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net390),
    .S1(net395),
    .X(_04191_));
 sky130_fd_sc_hd__mux4_2 _14549_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net390),
    .S1(net395),
    .X(_04192_));
 sky130_fd_sc_hd__mux4_2 _14550_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net390),
    .S1(net395),
    .X(_04193_));
 sky130_fd_sc_hd__mux4_2 _14551_ (.A0(_04190_),
    .A1(_04191_),
    .A2(_04192_),
    .A3(_04193_),
    .S0(net384),
    .S1(net542),
    .X(_04194_));
 sky130_fd_sc_hd__mux4_2 _14552_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net391),
    .S1(net397),
    .X(_04195_));
 sky130_fd_sc_hd__mux4_2 _14553_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net391),
    .S1(net397),
    .X(_04196_));
 sky130_fd_sc_hd__mux4_2 _14554_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net391),
    .S1(net397),
    .X(_04197_));
 sky130_fd_sc_hd__mux4_2 _14555_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net391),
    .S1(net397),
    .X(_04198_));
 sky130_fd_sc_hd__mux4_2 _14556_ (.A0(_04195_),
    .A1(_04196_),
    .A2(_04197_),
    .A3(_04198_),
    .S0(net384),
    .S1(net542),
    .X(_04199_));
 sky130_fd_sc_hd__mux2i_4 _14557_ (.A0(_04194_),
    .A1(_04199_),
    .S(net380),
    .Y(_12003_));
 sky130_fd_sc_hd__mux4_2 _14558_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net470),
    .S1(net474),
    .X(_04200_));
 sky130_fd_sc_hd__mux4_2 _14559_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net470),
    .S1(net474),
    .X(_04201_));
 sky130_fd_sc_hd__mux4_2 _14560_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net470),
    .S1(net474),
    .X(_04202_));
 sky130_fd_sc_hd__mux4_2 _14561_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net470),
    .S1(net474),
    .X(_04203_));
 sky130_fd_sc_hd__mux4_2 _14562_ (.A0(_04200_),
    .A1(_04201_),
    .A2(_04202_),
    .A3(_04203_),
    .S0(\count16_2[3] ),
    .S1(net459),
    .X(_04204_));
 sky130_fd_sc_hd__mux4_2 _14563_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net466),
    .S1(net474),
    .X(_04205_));
 sky130_fd_sc_hd__mux4_2 _14564_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net466),
    .S1(net474),
    .X(_04206_));
 sky130_fd_sc_hd__mux4_2 _14565_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net466),
    .S1(net474),
    .X(_04207_));
 sky130_fd_sc_hd__mux4_2 _14566_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net466),
    .S1(net474),
    .X(_04208_));
 sky130_fd_sc_hd__mux4_2 _14567_ (.A0(_04205_),
    .A1(_04206_),
    .A2(_04207_),
    .A3(_04208_),
    .S0(net463),
    .S1(net459),
    .X(_04209_));
 sky130_fd_sc_hd__mux2i_4 _14568_ (.A0(_04204_),
    .A1(_04209_),
    .S(net458),
    .Y(_12008_));
 sky130_fd_sc_hd__xnor2_1 _14569_ (.A(_02738_),
    .B(_04152_),
    .Y(_12013_));
 sky130_fd_sc_hd__xnor2_1 _14570_ (.A(_03530_),
    .B(_03755_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_2 _14571_ (.A(net1130),
    .B(_04210_),
    .Y(_12012_));
 sky130_fd_sc_hd__mux4_2 _14572_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04211_));
 sky130_fd_sc_hd__mux4_2 _14573_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04212_));
 sky130_fd_sc_hd__mux4_2 _14574_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04213_));
 sky130_fd_sc_hd__mux4_2 _14575_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04214_));
 sky130_fd_sc_hd__mux4_2 _14576_ (.A0(_04211_),
    .A1(_04212_),
    .A2(_04213_),
    .A3(_04214_),
    .S0(net386),
    .S1(net383),
    .X(_04215_));
 sky130_fd_sc_hd__mux4_2 _14577_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04216_));
 sky130_fd_sc_hd__mux4_2 _14578_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04217_));
 sky130_fd_sc_hd__mux4_2 _14579_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04218_));
 sky130_fd_sc_hd__mux4_2 _14580_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net388),
    .S1(net398),
    .X(_04219_));
 sky130_fd_sc_hd__mux4_2 _14581_ (.A0(_04216_),
    .A1(_04217_),
    .A2(_04218_),
    .A3(_04219_),
    .S0(net385),
    .S1(\count7_2[4] ),
    .X(_04220_));
 sky130_fd_sc_hd__mux2i_4 _14582_ (.A0(_04215_),
    .A1(_04220_),
    .S(net381),
    .Y(_12011_));
 sky130_fd_sc_hd__mux4_2 _14583_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net471),
    .S1(net476),
    .X(_04221_));
 sky130_fd_sc_hd__mux4_2 _14584_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net471),
    .S1(net476),
    .X(_04222_));
 sky130_fd_sc_hd__mux4_2 _14585_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net471),
    .S1(net476),
    .X(_04223_));
 sky130_fd_sc_hd__mux4_2 _14586_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net471),
    .S1(net476),
    .X(_04224_));
 sky130_fd_sc_hd__mux4_2 _14587_ (.A0(_04221_),
    .A1(_04222_),
    .A2(_04223_),
    .A3(_04224_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_04225_));
 sky130_fd_sc_hd__mux4_2 _14588_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net469),
    .S1(net473),
    .X(_04226_));
 sky130_fd_sc_hd__mux4_2 _14589_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net469),
    .S1(net473),
    .X(_04227_));
 sky130_fd_sc_hd__mux4_2 _14590_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net469),
    .S1(net473),
    .X(_04228_));
 sky130_fd_sc_hd__mux4_2 _14591_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net469),
    .S1(net473),
    .X(_04229_));
 sky130_fd_sc_hd__mux4_2 _14592_ (.A0(_04226_),
    .A1(_04227_),
    .A2(_04228_),
    .A3(_04229_),
    .S0(net463),
    .S1(net460),
    .X(_04230_));
 sky130_fd_sc_hd__mux2i_4 _14593_ (.A0(_04225_),
    .A1(_04230_),
    .S(net458),
    .Y(_12016_));
 sky130_fd_sc_hd__xnor2_1 _14594_ (.A(_02938_),
    .B(_04188_),
    .Y(_12021_));
 sky130_fd_sc_hd__xnor2_1 _14595_ (.A(_03590_),
    .B(_03815_),
    .Y(_04231_));
 sky130_fd_sc_hd__xnor2_1 _14596_ (.A(_03205_),
    .B(_04231_),
    .Y(_12020_));
 sky130_fd_sc_hd__mux4_2 _14597_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net387),
    .S1(net396),
    .X(_04232_));
 sky130_fd_sc_hd__mux4_2 _14598_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net387),
    .S1(net396),
    .X(_04233_));
 sky130_fd_sc_hd__mux4_2 _14599_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net387),
    .S1(net396),
    .X(_04234_));
 sky130_fd_sc_hd__mux4_2 _14600_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net387),
    .S1(net396),
    .X(_04235_));
 sky130_fd_sc_hd__mux4_2 _14601_ (.A0(_04232_),
    .A1(_04233_),
    .A2(_04234_),
    .A3(_04235_),
    .S0(net385),
    .S1(net382),
    .X(_04236_));
 sky130_fd_sc_hd__mux4_2 _14602_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net392),
    .S1(net396),
    .X(_04237_));
 sky130_fd_sc_hd__mux4_2 _14603_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net392),
    .S1(net396),
    .X(_04238_));
 sky130_fd_sc_hd__mux4_2 _14604_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net392),
    .S1(net396),
    .X(_04239_));
 sky130_fd_sc_hd__mux4_2 _14605_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net392),
    .S1(net396),
    .X(_04240_));
 sky130_fd_sc_hd__mux4_2 _14606_ (.A0(_04237_),
    .A1(_04238_),
    .A2(_04239_),
    .A3(_04240_),
    .S0(net385),
    .S1(net382),
    .X(_04241_));
 sky130_fd_sc_hd__mux2i_4 _14607_ (.A0(_04236_),
    .A1(_04241_),
    .S(net380),
    .Y(_12019_));
 sky130_fd_sc_hd__mux4_2 _14608_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net471),
    .S1(net476),
    .X(_04242_));
 sky130_fd_sc_hd__mux4_2 _14609_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net471),
    .S1(net476),
    .X(_04243_));
 sky130_fd_sc_hd__mux4_2 _14610_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net471),
    .S1(net476),
    .X(_04244_));
 sky130_fd_sc_hd__mux4_2 _14611_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net471),
    .S1(net476),
    .X(_04245_));
 sky130_fd_sc_hd__mux4_2 _14612_ (.A0(_04242_),
    .A1(_04243_),
    .A2(_04244_),
    .A3(_04245_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_04246_));
 sky130_fd_sc_hd__mux4_2 _14613_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net468),
    .S1(net476),
    .X(_04247_));
 sky130_fd_sc_hd__mux4_2 _14614_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net468),
    .S1(net476),
    .X(_04248_));
 sky130_fd_sc_hd__mux4_2 _14615_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net468),
    .S1(net476),
    .X(_04249_));
 sky130_fd_sc_hd__mux4_2 _14616_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net468),
    .S1(\count16_2[1] ),
    .X(_04250_));
 sky130_fd_sc_hd__mux4_2 _14617_ (.A0(_04247_),
    .A1(_04248_),
    .A2(_04249_),
    .A3(_04250_),
    .S0(net464),
    .S1(net461),
    .X(_04251_));
 sky130_fd_sc_hd__mux2i_4 _14618_ (.A0(_04246_),
    .A1(_04251_),
    .S(\count16_2[5] ),
    .Y(_12024_));
 sky130_fd_sc_hd__xnor2_1 _14619_ (.A(_02738_),
    .B(_03075_),
    .Y(_12029_));
 sky130_fd_sc_hd__xnor2_1 _14620_ (.A(_03645_),
    .B(_03864_),
    .Y(_04252_));
 sky130_fd_sc_hd__xnor2_2 _14621_ (.A(_03275_),
    .B(_04252_),
    .Y(_12028_));
 sky130_fd_sc_hd__mux4_2 _14622_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04253_));
 sky130_fd_sc_hd__mux4_2 _14623_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04254_));
 sky130_fd_sc_hd__mux4_2 _14624_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04255_));
 sky130_fd_sc_hd__mux4_2 _14625_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04256_));
 sky130_fd_sc_hd__mux4_2 _14626_ (.A0(_04253_),
    .A1(_04254_),
    .A2(_04255_),
    .A3(_04256_),
    .S0(net385),
    .S1(net382),
    .X(_04257_));
 sky130_fd_sc_hd__mux4_2 _14627_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04258_));
 sky130_fd_sc_hd__mux4_2 _14628_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04259_));
 sky130_fd_sc_hd__mux4_2 _14629_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04260_));
 sky130_fd_sc_hd__mux4_2 _14630_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net387),
    .S1(net396),
    .X(_04261_));
 sky130_fd_sc_hd__mux4_2 _14631_ (.A0(_04258_),
    .A1(_04259_),
    .A2(_04260_),
    .A3(_04261_),
    .S0(net385),
    .S1(net382),
    .X(_04262_));
 sky130_fd_sc_hd__mux2i_4 _14632_ (.A0(_04257_),
    .A1(_04262_),
    .S(net380),
    .Y(_12027_));
 sky130_fd_sc_hd__mux4_2 _14633_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net466),
    .S1(net474),
    .X(_04263_));
 sky130_fd_sc_hd__mux4_2 _14634_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net466),
    .S1(net474),
    .X(_04264_));
 sky130_fd_sc_hd__mux4_2 _14635_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net466),
    .S1(net474),
    .X(_04265_));
 sky130_fd_sc_hd__mux4_2 _14636_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net466),
    .S1(net474),
    .X(_04266_));
 sky130_fd_sc_hd__mux4_2 _14637_ (.A0(_04263_),
    .A1(_04264_),
    .A2(_04265_),
    .A3(_04266_),
    .S0(net462),
    .S1(net460),
    .X(_04267_));
 sky130_fd_sc_hd__mux4_2 _14638_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net469),
    .S1(net474),
    .X(_04268_));
 sky130_fd_sc_hd__mux4_2 _14639_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net469),
    .S1(net474),
    .X(_04269_));
 sky130_fd_sc_hd__mux4_2 _14640_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net469),
    .S1(net474),
    .X(_04270_));
 sky130_fd_sc_hd__mux4_2 _14641_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net469),
    .S1(net474),
    .X(_04271_));
 sky130_fd_sc_hd__mux4_2 _14642_ (.A0(_04268_),
    .A1(_04269_),
    .A2(_04270_),
    .A3(_04271_),
    .S0(net463),
    .S1(net459),
    .X(_04272_));
 sky130_fd_sc_hd__mux2i_4 _14643_ (.A0(_04267_),
    .A1(_04272_),
    .S(net457),
    .Y(_12032_));
 sky130_fd_sc_hd__xnor2_1 _14644_ (.A(_02938_),
    .B(_03157_),
    .Y(_12037_));
 sky130_fd_sc_hd__xnor2_1 _14645_ (.A(_03709_),
    .B(_03910_),
    .Y(_04273_));
 sky130_fd_sc_hd__xnor2_2 _14646_ (.A(_03344_),
    .B(_04273_),
    .Y(_12036_));
 sky130_fd_sc_hd__mux4_2 _14647_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net387),
    .S1(net396),
    .X(_04274_));
 sky130_fd_sc_hd__mux4_2 _14648_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net387),
    .S1(net396),
    .X(_04275_));
 sky130_fd_sc_hd__mux4_2 _14649_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net387),
    .S1(net396),
    .X(_04276_));
 sky130_fd_sc_hd__mux4_2 _14650_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net387),
    .S1(net396),
    .X(_04277_));
 sky130_fd_sc_hd__mux4_2 _14651_ (.A0(_04274_),
    .A1(_04275_),
    .A2(_04276_),
    .A3(_04277_),
    .S0(net385),
    .S1(net382),
    .X(_04278_));
 sky130_fd_sc_hd__mux4_2 _14652_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net392),
    .S1(net396),
    .X(_04279_));
 sky130_fd_sc_hd__mux4_2 _14653_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net392),
    .S1(net396),
    .X(_04280_));
 sky130_fd_sc_hd__mux4_2 _14654_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net392),
    .S1(net396),
    .X(_04281_));
 sky130_fd_sc_hd__mux4_2 _14655_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net392),
    .S1(net396),
    .X(_04282_));
 sky130_fd_sc_hd__mux4_2 _14656_ (.A0(_04279_),
    .A1(_04280_),
    .A2(_04281_),
    .A3(_04282_),
    .S0(net385),
    .S1(net382),
    .X(_04283_));
 sky130_fd_sc_hd__mux2i_4 _14657_ (.A0(_04278_),
    .A1(_04283_),
    .S(net380),
    .Y(_12035_));
 sky130_fd_sc_hd__mux4_2 _14658_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net471),
    .S1(net553),
    .X(_04284_));
 sky130_fd_sc_hd__mux4_2 _14659_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net471),
    .S1(net553),
    .X(_04285_));
 sky130_fd_sc_hd__mux4_2 _14660_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net471),
    .S1(net553),
    .X(_04286_));
 sky130_fd_sc_hd__mux4_2 _14661_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net471),
    .S1(net553),
    .X(_04287_));
 sky130_fd_sc_hd__mux4_2 _14662_ (.A0(_04284_),
    .A1(_04285_),
    .A2(_04286_),
    .A3(_04287_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_04288_));
 sky130_fd_sc_hd__mux4_2 _14663_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net469),
    .S1(net473),
    .X(_04289_));
 sky130_fd_sc_hd__mux4_2 _14664_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net469),
    .S1(net473),
    .X(_04290_));
 sky130_fd_sc_hd__mux4_2 _14665_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net471),
    .S1(net473),
    .X(_04291_));
 sky130_fd_sc_hd__mux4_2 _14666_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net469),
    .S1(net473),
    .X(_04292_));
 sky130_fd_sc_hd__mux4_2 _14667_ (.A0(_04289_),
    .A1(_04290_),
    .A2(_04291_),
    .A3(_04292_),
    .S0(net463),
    .S1(net461),
    .X(_04293_));
 sky130_fd_sc_hd__mux2i_2 _14668_ (.A0(_04288_),
    .A1(_04293_),
    .S(net458),
    .Y(_12040_));
 sky130_fd_sc_hd__xnor2_1 _14669_ (.A(_03075_),
    .B(_03239_),
    .Y(_12045_));
 sky130_fd_sc_hd__xnor2_1 _14670_ (.A(_03755_),
    .B(_03956_),
    .Y(_04294_));
 sky130_fd_sc_hd__xnor2_2 _14671_ (.A(_03402_),
    .B(_04294_),
    .Y(_12044_));
 sky130_fd_sc_hd__mux4_2 _14672_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04295_));
 sky130_fd_sc_hd__mux4_2 _14673_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04296_));
 sky130_fd_sc_hd__mux4_2 _14674_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04297_));
 sky130_fd_sc_hd__mux4_2 _14675_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04298_));
 sky130_fd_sc_hd__mux4_2 _14676_ (.A0(_04295_),
    .A1(_04296_),
    .A2(_04297_),
    .A3(_04298_),
    .S0(net386),
    .S1(net383),
    .X(_04299_));
 sky130_fd_sc_hd__mux4_2 _14677_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04300_));
 sky130_fd_sc_hd__mux4_2 _14678_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04301_));
 sky130_fd_sc_hd__mux4_2 _14679_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04302_));
 sky130_fd_sc_hd__mux4_2 _14680_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net389),
    .S1(net398),
    .X(_04303_));
 sky130_fd_sc_hd__mux4_2 _14681_ (.A0(_04300_),
    .A1(_04301_),
    .A2(_04302_),
    .A3(_04303_),
    .S0(net386),
    .S1(net383),
    .X(_04304_));
 sky130_fd_sc_hd__mux2i_4 _14682_ (.A0(_04299_),
    .A1(_04304_),
    .S(net381),
    .Y(_12043_));
 sky130_fd_sc_hd__mux4_2 _14683_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net465),
    .S1(net475),
    .X(_04305_));
 sky130_fd_sc_hd__mux4_2 _14684_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net465),
    .S1(net475),
    .X(_04306_));
 sky130_fd_sc_hd__mux4_2 _14685_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net465),
    .S1(net475),
    .X(_04307_));
 sky130_fd_sc_hd__mux4_2 _14686_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net465),
    .S1(net475),
    .X(_04308_));
 sky130_fd_sc_hd__mux4_2 _14687_ (.A0(_04305_),
    .A1(_04306_),
    .A2(_04307_),
    .A3(_04308_),
    .S0(net462),
    .S1(net460),
    .X(_04309_));
 sky130_fd_sc_hd__mux4_2 _14688_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net467),
    .S1(net473),
    .X(_04310_));
 sky130_fd_sc_hd__mux4_2 _14689_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net467),
    .S1(net473),
    .X(_04311_));
 sky130_fd_sc_hd__mux4_2 _14690_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net467),
    .S1(net473),
    .X(_04312_));
 sky130_fd_sc_hd__mux4_2 _14691_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net469),
    .S1(net473),
    .X(_04313_));
 sky130_fd_sc_hd__mux4_2 _14692_ (.A0(_04310_),
    .A1(_04311_),
    .A2(_04312_),
    .A3(_04313_),
    .S0(net463),
    .S1(net460),
    .X(_04314_));
 sky130_fd_sc_hd__mux2i_4 _14693_ (.A0(_04309_),
    .A1(_04314_),
    .S(net458),
    .Y(_12048_));
 sky130_fd_sc_hd__xnor2_1 _14694_ (.A(_03157_),
    .B(_03309_),
    .Y(_12053_));
 sky130_fd_sc_hd__xnor2_1 _14695_ (.A(_03460_),
    .B(_03815_),
    .Y(_04315_));
 sky130_fd_sc_hd__xnor2_1 _14696_ (.A(_02824_),
    .B(_04315_),
    .Y(_12052_));
 sky130_fd_sc_hd__mux4_2 _14697_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net388),
    .S1(net398),
    .X(_04316_));
 sky130_fd_sc_hd__mux4_2 _14698_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net388),
    .S1(net398),
    .X(_04317_));
 sky130_fd_sc_hd__mux4_2 _14699_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net388),
    .S1(net398),
    .X(_04318_));
 sky130_fd_sc_hd__mux4_2 _14700_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net388),
    .S1(net398),
    .X(_04319_));
 sky130_fd_sc_hd__mux4_2 _14701_ (.A0(_04316_),
    .A1(_04317_),
    .A2(_04318_),
    .A3(_04319_),
    .S0(net386),
    .S1(net382),
    .X(_04320_));
 sky130_fd_sc_hd__mux4_2 _14702_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net391),
    .S1(net397),
    .X(_04321_));
 sky130_fd_sc_hd__mux4_2 _14703_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net392),
    .S1(net396),
    .X(_04322_));
 sky130_fd_sc_hd__mux4_2 _14704_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net392),
    .S1(net396),
    .X(_04323_));
 sky130_fd_sc_hd__mux4_2 _14705_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net392),
    .S1(net397),
    .X(_04324_));
 sky130_fd_sc_hd__mux4_2 _14706_ (.A0(_04321_),
    .A1(_04322_),
    .A2(_04323_),
    .A3(_04324_),
    .S0(net385),
    .S1(net382),
    .X(_04325_));
 sky130_fd_sc_hd__mux2i_4 _14707_ (.A0(_04320_),
    .A1(_04325_),
    .S(net380),
    .Y(_12051_));
 sky130_fd_sc_hd__mux4_2 _14708_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net471),
    .S1(net476),
    .X(_04326_));
 sky130_fd_sc_hd__mux4_2 _14709_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net471),
    .S1(net476),
    .X(_04327_));
 sky130_fd_sc_hd__mux4_2 _14710_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net471),
    .S1(net476),
    .X(_04328_));
 sky130_fd_sc_hd__mux4_2 _14711_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net471),
    .S1(net476),
    .X(_04329_));
 sky130_fd_sc_hd__mux4_2 _14712_ (.A0(_04326_),
    .A1(_04327_),
    .A2(_04328_),
    .A3(_04329_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_04330_));
 sky130_fd_sc_hd__mux4_2 _14713_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net468),
    .S1(\count16_2[1] ),
    .X(_04331_));
 sky130_fd_sc_hd__mux4_2 _14714_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net468),
    .S1(net476),
    .X(_04332_));
 sky130_fd_sc_hd__mux4_2 _14715_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net468),
    .S1(net476),
    .X(_04333_));
 sky130_fd_sc_hd__mux4_2 _14716_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net468),
    .S1(net476),
    .X(_04334_));
 sky130_fd_sc_hd__mux4_2 _14717_ (.A0(_04331_),
    .A1(_04332_),
    .A2(_04333_),
    .A3(_04334_),
    .S0(net464),
    .S1(net461),
    .X(_04335_));
 sky130_fd_sc_hd__mux2i_4 _14718_ (.A0(_04330_),
    .A1(_04335_),
    .S(\count16_2[5] ),
    .Y(_12056_));
 sky130_fd_sc_hd__xnor2_1 _14719_ (.A(_03239_),
    .B(_03378_),
    .Y(_12061_));
 sky130_fd_sc_hd__xnor2_1 _14720_ (.A(_02976_),
    .B(_03519_),
    .Y(_12060_));
 sky130_fd_sc_hd__mux4_2 _14721_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net543),
    .S1(net394),
    .X(_04336_));
 sky130_fd_sc_hd__mux4_2 _14722_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net543),
    .S1(net394),
    .X(_04337_));
 sky130_fd_sc_hd__mux4_2 _14723_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net543),
    .S1(net394),
    .X(_04338_));
 sky130_fd_sc_hd__mux4_2 _14724_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net543),
    .S1(net394),
    .X(_04339_));
 sky130_fd_sc_hd__mux4_2 _14725_ (.A0(_04336_),
    .A1(_04337_),
    .A2(_04338_),
    .A3(_04339_),
    .S0(net386),
    .S1(net383),
    .X(_04340_));
 sky130_fd_sc_hd__mux4_2 _14726_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net393),
    .S1(net394),
    .X(_04341_));
 sky130_fd_sc_hd__mux4_2 _14727_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net393),
    .S1(net394),
    .X(_04342_));
 sky130_fd_sc_hd__mux4_2 _14728_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net393),
    .S1(net394),
    .X(_04343_));
 sky130_fd_sc_hd__mux4_2 _14729_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net393),
    .S1(net394),
    .X(_04344_));
 sky130_fd_sc_hd__mux4_2 _14730_ (.A0(_04341_),
    .A1(_04342_),
    .A2(_04343_),
    .A3(_04344_),
    .S0(net386),
    .S1(net383),
    .X(_04345_));
 sky130_fd_sc_hd__mux2i_4 _14731_ (.A0(_04340_),
    .A1(_04345_),
    .S(\count7_2[5] ),
    .Y(_12059_));
 sky130_fd_sc_hd__mux4_2 _14732_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net471),
    .S1(net476),
    .X(_04346_));
 sky130_fd_sc_hd__mux4_2 _14733_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net471),
    .S1(net476),
    .X(_04347_));
 sky130_fd_sc_hd__mux4_2 _14734_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net471),
    .S1(net476),
    .X(_04348_));
 sky130_fd_sc_hd__mux4_2 _14735_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net471),
    .S1(net476),
    .X(_04349_));
 sky130_fd_sc_hd__mux4_2 _14736_ (.A0(_04346_),
    .A1(_04347_),
    .A2(_04348_),
    .A3(_04349_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_04350_));
 sky130_fd_sc_hd__mux4_2 _14737_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net469),
    .S1(\count16_2[1] ),
    .X(_04351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1427 ();
 sky130_fd_sc_hd__mux4_2 _14739_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net468),
    .S1(\count16_2[1] ),
    .X(_04353_));
 sky130_fd_sc_hd__mux4_2 _14740_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net468),
    .S1(\count16_2[1] ),
    .X(_04354_));
 sky130_fd_sc_hd__mux4_2 _14741_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net468),
    .S1(\count16_2[1] ),
    .X(_04355_));
 sky130_fd_sc_hd__mux4_2 _14742_ (.A0(_04351_),
    .A1(_04353_),
    .A2(_04354_),
    .A3(_04355_),
    .S0(net464),
    .S1(net461),
    .X(_04356_));
 sky130_fd_sc_hd__mux2i_4 _14743_ (.A0(_04350_),
    .A1(_04356_),
    .S(\count16_2[5] ),
    .Y(_12064_));
 sky130_fd_sc_hd__xnor2_1 _14744_ (.A(_02788_),
    .B(_03309_),
    .Y(_12069_));
 sky130_fd_sc_hd__xnor2_1 _14745_ (.A(_03098_),
    .B(_03579_),
    .Y(_12068_));
 sky130_fd_sc_hd__mux4_2 _14746_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net543),
    .S1(net394),
    .X(_04357_));
 sky130_fd_sc_hd__mux4_2 _14747_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net543),
    .S1(net394),
    .X(_04358_));
 sky130_fd_sc_hd__mux4_2 _14748_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net543),
    .S1(net394),
    .X(_04359_));
 sky130_fd_sc_hd__mux4_2 _14749_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net543),
    .S1(net394),
    .X(_04360_));
 sky130_fd_sc_hd__mux4_2 _14750_ (.A0(_04357_),
    .A1(_04358_),
    .A2(_04359_),
    .A3(_04360_),
    .S0(\count7_2[3] ),
    .S1(net383),
    .X(_04361_));
 sky130_fd_sc_hd__mux4_2 _14751_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net393),
    .S1(net394),
    .X(_04362_));
 sky130_fd_sc_hd__mux4_2 _14752_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net393),
    .S1(net394),
    .X(_04363_));
 sky130_fd_sc_hd__mux4_2 _14753_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net393),
    .S1(net394),
    .X(_04364_));
 sky130_fd_sc_hd__mux4_2 _14754_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net393),
    .S1(net394),
    .X(_04365_));
 sky130_fd_sc_hd__mux4_2 _14755_ (.A0(_04362_),
    .A1(_04363_),
    .A2(_04364_),
    .A3(_04365_),
    .S0(net386),
    .S1(net383),
    .X(_04366_));
 sky130_fd_sc_hd__mux2i_4 _14756_ (.A0(_04361_),
    .A1(_04366_),
    .S(\count7_2[5] ),
    .Y(_12067_));
 sky130_fd_sc_hd__mux4_2 _14757_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_04367_));
 sky130_fd_sc_hd__mux4_2 _14758_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_04368_));
 sky130_fd_sc_hd__mux4_2 _14759_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_04369_));
 sky130_fd_sc_hd__mux4_2 _14760_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_04370_));
 sky130_fd_sc_hd__mux4_2 _14761_ (.A0(_04367_),
    .A1(_04368_),
    .A2(_04369_),
    .A3(_04370_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_04371_));
 sky130_fd_sc_hd__mux4_2 _14762_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net472),
    .S1(net477),
    .X(_04372_));
 sky130_fd_sc_hd__mux4_2 _14763_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net472),
    .S1(net477),
    .X(_04373_));
 sky130_fd_sc_hd__mux4_2 _14764_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net472),
    .S1(net477),
    .X(_04374_));
 sky130_fd_sc_hd__mux4_2 _14765_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net472),
    .S1(net477),
    .X(_04375_));
 sky130_fd_sc_hd__mux4_2 _14766_ (.A0(_04372_),
    .A1(_04373_),
    .A2(_04374_),
    .A3(_04375_),
    .S0(\count16_2[3] ),
    .S1(net461),
    .X(_04376_));
 sky130_fd_sc_hd__mux2i_1 _14767_ (.A0(_04371_),
    .A1(_04376_),
    .S(net458),
    .Y(_12072_));
 sky130_fd_sc_hd__a21o_1 _14768_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_12922_),
    .B1(\hash.CA2.b_dash[0] ),
    .X(_04377_));
 sky130_fd_sc_hd__o21ai_2 _14769_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_12922_),
    .B1(_04377_),
    .Y(_12077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1424 ();
 sky130_fd_sc_hd__xnor2_4 _14773_ (.A(\hash.CA2.S1.X[6] ),
    .B(\hash.CA2.S1.X[25] ),
    .Y(_04381_));
 sky130_fd_sc_hd__xnor2_4 _14774_ (.A(\hash.CA2.S1.X[11] ),
    .B(_04381_),
    .Y(_13230_));
 sky130_fd_sc_hd__a21o_1 _14775_ (.A1(_12956_),
    .A2(_12953_),
    .B1(_12955_),
    .X(_04382_));
 sky130_fd_sc_hd__a21oi_1 _14776_ (.A1(_12958_),
    .A2(_04382_),
    .B1(_12957_),
    .Y(_04383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1423 ();
 sky130_fd_sc_hd__nand2_1 _14778_ (.A(_12962_),
    .B(_12964_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _14779_ (.A(_12962_),
    .B(_12963_),
    .Y(_04386_));
 sky130_fd_sc_hd__o21ai_1 _14780_ (.A1(_04383_),
    .A2(_04385_),
    .B1(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1422 ();
 sky130_fd_sc_hd__nand3_1 _14782_ (.A(_12946_),
    .B(_12950_),
    .C(_12952_),
    .Y(_04389_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1421 ();
 sky130_fd_sc_hd__nor2_1 _14784_ (.A(_12948_),
    .B(_12947_),
    .Y(_04391_));
 sky130_fd_sc_hd__a21o_1 _14785_ (.A1(_12952_),
    .A2(_12945_),
    .B1(_12951_),
    .X(_04392_));
 sky130_fd_sc_hd__a21oi_2 _14786_ (.A1(_12950_),
    .A2(_04392_),
    .B1(_12949_),
    .Y(_04393_));
 sky130_fd_sc_hd__o21a_4 _14787_ (.A1(_04389_),
    .A2(_04391_),
    .B1(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1420 ();
 sky130_fd_sc_hd__or2_4 _14789_ (.A(_12930_),
    .B(_12929_),
    .X(_04396_));
 sky130_fd_sc_hd__a21o_4 _14790_ (.A1(_12928_),
    .A2(_04396_),
    .B1(_12927_),
    .X(_04397_));
 sky130_fd_sc_hd__a211oi_4 _14791_ (.A1(_12924_),
    .A2(_12081_),
    .B1(_12923_),
    .C1(_12935_),
    .Y(_04398_));
 sky130_fd_sc_hd__o211ai_1 _14792_ (.A1(_12936_),
    .A2(_12935_),
    .B1(_12932_),
    .C1(_12934_),
    .Y(_04399_));
 sky130_fd_sc_hd__a21oi_2 _14793_ (.A1(_12932_),
    .A2(_12933_),
    .B1(_12931_),
    .Y(_04400_));
 sky130_fd_sc_hd__nor2_1 _14794_ (.A(_12927_),
    .B(_12929_),
    .Y(_04401_));
 sky130_fd_sc_hd__o211ai_1 _14795_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04400_),
    .C1(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__clkinv_1 _14796_ (.A(_12944_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_4 _14797_ (.A(_12938_),
    .B(_12942_),
    .Y(_04404_));
 sky130_fd_sc_hd__nor2_1 _14798_ (.A(_04403_),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__and4_4 _14799_ (.A(_12940_),
    .B(_04397_),
    .C(_04402_),
    .D(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__nand2_1 _14800_ (.A(_12944_),
    .B(_12939_),
    .Y(_04407_));
 sky130_fd_sc_hd__a21oi_2 _14801_ (.A1(_12942_),
    .A2(_12937_),
    .B1(_12941_),
    .Y(_04408_));
 sky130_fd_sc_hd__o22ai_2 _14802_ (.A1(_04404_),
    .A2(_04407_),
    .B1(_04408_),
    .B2(_04403_),
    .Y(_04409_));
 sky130_fd_sc_hd__nor2_1 _14803_ (.A(_12943_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nor4bb_4 _14804_ (.A(_12947_),
    .B(_04406_),
    .C_N(_04410_),
    .D_N(_04393_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand3_1 _14805_ (.A(_12954_),
    .B(_12956_),
    .C(_12958_),
    .Y(_04412_));
 sky130_fd_sc_hd__or4_4 _14806_ (.A(_04411_),
    .B(_04385_),
    .C(_04412_),
    .D(_04394_),
    .X(_04413_));
 sky130_fd_sc_hd__nand2b_1 _14807_ (.A_N(_04387_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__o21ai_2 _14808_ (.A1(_12961_),
    .A2(_04414_),
    .B1(_12960_),
    .Y(_04415_));
 sky130_fd_sc_hd__nor2_2 _14809_ (.A(_12966_),
    .B(_12959_),
    .Y(_04416_));
 sky130_fd_sc_hd__nor3_2 _14810_ (.A(_12959_),
    .B(_12961_),
    .C(_04387_),
    .Y(_04417_));
 sky130_fd_sc_hd__o21ai_2 _14811_ (.A1(_12960_),
    .A2(_12959_),
    .B1(_12966_),
    .Y(_04418_));
 sky130_fd_sc_hd__a21oi_4 _14812_ (.A1(_04417_),
    .A2(_04413_),
    .B1(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__a21oi_4 _14813_ (.A1(_04415_),
    .A2(_04416_),
    .B1(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__xor2_4 _14814_ (.A(_12924_),
    .B(net1097),
    .X(_04421_));
 sky130_fd_sc_hd__o31a_1 _14815_ (.A1(_12932_),
    .A2(_12929_),
    .A3(_12931_),
    .B1(_04396_),
    .X(_04422_));
 sky130_fd_sc_hd__a211oi_1 _14816_ (.A1(_12080_),
    .A2(_12926_),
    .B1(_12923_),
    .C1(_12925_),
    .Y(_04423_));
 sky130_fd_sc_hd__o211ai_1 _14817_ (.A1(_12924_),
    .A2(_12923_),
    .B1(_12936_),
    .C1(_12934_),
    .Y(_04424_));
 sky130_fd_sc_hd__a21oi_1 _14818_ (.A1(_12934_),
    .A2(_12935_),
    .B1(_12933_),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_1 _14819_ (.A(_12929_),
    .B(_12931_),
    .Y(_04426_));
 sky130_fd_sc_hd__o211ai_1 _14820_ (.A1(_04424_),
    .A2(_04423_),
    .B1(_04425_),
    .C1(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_4 _14821_ (.A(_04422_),
    .B(net1099),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_1 _14822_ (.A(_12928_),
    .B(_12940_),
    .Y(_04429_));
 sky130_fd_sc_hd__nor2_1 _14823_ (.A(_04404_),
    .B(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__nand2_1 _14824_ (.A(_12944_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__a21oi_2 _14825_ (.A1(_12940_),
    .A2(_12927_),
    .B1(_12939_),
    .Y(_04432_));
 sky130_fd_sc_hd__o21ai_4 _14826_ (.A1(_04404_),
    .A2(_04432_),
    .B1(_04408_),
    .Y(_04433_));
 sky130_fd_sc_hd__a21oi_1 _14827_ (.A1(_12944_),
    .A2(_04433_),
    .B1(_12943_),
    .Y(_04434_));
 sky130_fd_sc_hd__o21ai_2 _14828_ (.A1(_04428_),
    .A2(_04431_),
    .B1(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__a21oi_4 _14829_ (.A1(_12948_),
    .A2(_04435_),
    .B1(_12947_),
    .Y(_04436_));
 sky130_fd_sc_hd__xnor2_4 _14830_ (.A(_12946_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1419 ();
 sky130_fd_sc_hd__xor2_1 _14832_ (.A(_04421_),
    .B(_04437_),
    .X(_04439_));
 sky130_fd_sc_hd__xnor2_2 _14833_ (.A(_04420_),
    .B(_04439_),
    .Y(_12075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1418 ();
 sky130_fd_sc_hd__nor2_4 _14835_ (.A(net349),
    .B(_13235_),
    .Y(_00658_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1417 ();
 sky130_fd_sc_hd__a21o_1 _14837_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_12082_),
    .B1(\hash.CA2.b_dash[1] ),
    .X(_04442_));
 sky130_fd_sc_hd__o21ai_2 _14838_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_12082_),
    .B1(_04442_),
    .Y(_12089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1414 ();
 sky130_fd_sc_hd__xnor2_2 _14842_ (.A(\hash.CA2.S1.X[7] ),
    .B(\hash.CA2.S1.X[26] ),
    .Y(_04446_));
 sky130_fd_sc_hd__xnor2_2 _14843_ (.A(\hash.CA2.S1.X[12] ),
    .B(_04446_),
    .Y(_13237_));
 sky130_fd_sc_hd__inv_1 _14844_ (.A(net1049),
    .Y(_12085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1413 ();
 sky130_fd_sc_hd__mux2_1 _14846_ (.A0(\hash.CA2.f_dash[1] ),
    .A1(\hash.CA2.e_dash[1] ),
    .S(\hash.CA2.S1.X[1] ),
    .X(_13236_));
 sky130_fd_sc_hd__inv_1 _14847_ (.A(_13236_),
    .Y(_12084_));
 sky130_fd_sc_hd__a21o_1 _14848_ (.A1(_12954_),
    .A2(_12949_),
    .B1(_12953_),
    .X(_04448_));
 sky130_fd_sc_hd__a21o_1 _14849_ (.A1(_12956_),
    .A2(_04448_),
    .B1(_12955_),
    .X(_04449_));
 sky130_fd_sc_hd__a21o_4 _14850_ (.A1(_12958_),
    .A2(_04449_),
    .B1(_12957_),
    .X(_04450_));
 sky130_fd_sc_hd__a21o_1 _14851_ (.A1(_12948_),
    .A2(_12943_),
    .B1(_12947_),
    .X(_04451_));
 sky130_fd_sc_hd__a21o_1 _14852_ (.A1(_12946_),
    .A2(_04451_),
    .B1(_12945_),
    .X(_04452_));
 sky130_fd_sc_hd__a21o_4 _14853_ (.A1(_12952_),
    .A2(_04452_),
    .B1(_12951_),
    .X(_04453_));
 sky130_fd_sc_hd__inv_1 _14854_ (.A(_12964_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand4_1 _14855_ (.A(_12950_),
    .B(_12954_),
    .C(_12956_),
    .D(_12958_),
    .Y(_04455_));
 sky130_fd_sc_hd__nor2_2 _14856_ (.A(_04454_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__a22oi_2 _14857_ (.A1(_12964_),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__and3_4 _14858_ (.A(_04422_),
    .B(_04427_),
    .C(_04430_),
    .X(_04458_));
 sky130_fd_sc_hd__nand4_1 _14859_ (.A(_12946_),
    .B(_12944_),
    .C(_12948_),
    .D(_12952_),
    .Y(_04459_));
 sky130_fd_sc_hd__inv_1 _14860_ (.A(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__o211ai_1 _14861_ (.A1(_04458_),
    .A2(_04433_),
    .B1(_04460_),
    .C1(_04456_),
    .Y(_04461_));
 sky130_fd_sc_hd__nor3_1 _14862_ (.A(_12959_),
    .B(_12961_),
    .C(_12963_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand3_2 _14863_ (.A(_04457_),
    .B(net1091),
    .C(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__o21ai_1 _14864_ (.A1(_12962_),
    .A2(_12961_),
    .B1(_12960_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2b_2 _14865_ (.A_N(_12959_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__a31oi_2 _14866_ (.A1(_12966_),
    .A2(_04463_),
    .A3(_04465_),
    .B1(_12965_),
    .Y(_04466_));
 sky130_fd_sc_hd__xnor2_4 _14867_ (.A(_12970_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__a21o_1 _14868_ (.A1(_12080_),
    .A2(_12926_),
    .B1(_12925_),
    .X(_04468_));
 sky130_fd_sc_hd__a21oi_2 _14869_ (.A1(_12924_),
    .A2(_04468_),
    .B1(_12923_),
    .Y(_04469_));
 sky130_fd_sc_hd__xnor2_4 _14870_ (.A(_12936_),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__inv_1 _14871_ (.A(_12948_),
    .Y(_04471_));
 sky130_fd_sc_hd__nor3_4 _14872_ (.A(_12943_),
    .B(_04406_),
    .C(_04409_),
    .Y(_04472_));
 sky130_fd_sc_hd__o21bai_1 _14873_ (.A1(_04471_),
    .A2(_04472_),
    .B1_N(_12947_),
    .Y(_04473_));
 sky130_fd_sc_hd__a21o_4 _14874_ (.A1(_12946_),
    .A2(_04473_),
    .B1(_12945_),
    .X(_04474_));
 sky130_fd_sc_hd__xnor2_4 _14875_ (.A(_04474_),
    .B(_12952_),
    .Y(_04475_));
 sky130_fd_sc_hd__xnor2_1 _14876_ (.A(_04470_),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__xnor2_1 _14877_ (.A(_04467_),
    .B(_04476_),
    .Y(_12088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1412 ();
 sky130_fd_sc_hd__or2_0 _14879_ (.A(net349),
    .B(_13241_),
    .X(\hash.CA1.S0.X[1] ));
 sky130_fd_sc_hd__inv_1 _14880_ (.A(\hash.CA1.S0.X[1] ),
    .Y(_13543_));
 sky130_fd_sc_hd__a21o_1 _14881_ (.A1(\hash.CA2.a_dash[2] ),
    .A2(_04421_),
    .B1(\hash.CA2.b_dash[2] ),
    .X(_04478_));
 sky130_fd_sc_hd__o21ai_2 _14882_ (.A1(\hash.CA2.a_dash[2] ),
    .A2(_04421_),
    .B1(_04478_),
    .Y(_12098_));
 sky130_fd_sc_hd__xnor2_2 _14883_ (.A(net1083),
    .B(_13245_),
    .Y(_13246_));
 sky130_fd_sc_hd__inv_4 _14884_ (.A(_13246_),
    .Y(_12097_));
 sky130_fd_sc_hd__o21a_1 _14885_ (.A1(_12965_),
    .A2(_04419_),
    .B1(_12970_),
    .X(_04479_));
 sky130_fd_sc_hd__nor2_4 _14886_ (.A(_12969_),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__xor2_4 _14887_ (.A(_12968_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__o21a_4 _14888_ (.A1(_04433_),
    .A2(_04458_),
    .B1(_04460_),
    .X(_04482_));
 sky130_fd_sc_hd__nor2_4 _14889_ (.A(_04453_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__xnor2_4 _14890_ (.A(_12950_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__a21o_1 _14891_ (.A1(_12924_),
    .A2(_12081_),
    .B1(_12923_),
    .X(_04485_));
 sky130_fd_sc_hd__a21oi_2 _14892_ (.A1(_12936_),
    .A2(_04485_),
    .B1(_12935_),
    .Y(_04486_));
 sky130_fd_sc_hd__xnor2_4 _14893_ (.A(_12934_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__xnor2_1 _14894_ (.A(_04484_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__xnor2_2 _14895_ (.A(_04481_),
    .B(_04488_),
    .Y(_12096_));
 sky130_fd_sc_hd__maj3_1 _14896_ (.A(\hash.CA2.b_dash[3] ),
    .B(\hash.CA2.a_dash[3] ),
    .C(_04470_),
    .X(_04489_));
 sky130_fd_sc_hd__clkinv_1 _14897_ (.A(_04489_),
    .Y(_12112_));
 sky130_fd_sc_hd__a21o_1 _14898_ (.A1(_13231_),
    .A2(_13239_),
    .B1(_13238_),
    .X(_04490_));
 sky130_fd_sc_hd__a21oi_1 _14899_ (.A1(_13245_),
    .A2(_04490_),
    .B1(_13244_),
    .Y(_04491_));
 sky130_fd_sc_hd__xnor2_2 _14900_ (.A(_13252_),
    .B(_04491_),
    .Y(_13253_));
 sky130_fd_sc_hd__inv_4 _14901_ (.A(_13253_),
    .Y(_12111_));
 sky130_fd_sc_hd__clkinv_2 _14902_ (.A(_12972_),
    .Y(_04492_));
 sky130_fd_sc_hd__o21ai_0 _14903_ (.A1(_12966_),
    .A2(_12965_),
    .B1(_12970_),
    .Y(_04493_));
 sky130_fd_sc_hd__nor2_1 _14904_ (.A(_12967_),
    .B(_12969_),
    .Y(_04494_));
 sky130_fd_sc_hd__nor2_1 _14905_ (.A(_12968_),
    .B(_12967_),
    .Y(_04495_));
 sky130_fd_sc_hd__a21oi_2 _14906_ (.A1(_04493_),
    .A2(_04494_),
    .B1(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__a2111o_2 _14907_ (.A1(_04463_),
    .A2(_04465_),
    .B1(_12965_),
    .C1(_12967_),
    .D1(_12969_),
    .X(_04497_));
 sky130_fd_sc_hd__nand2_4 _14908_ (.A(_04496_),
    .B(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__xnor2_4 _14909_ (.A(_04492_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__o21ai_2 _14910_ (.A1(_04423_),
    .A2(_04424_),
    .B1(_04425_),
    .Y(_04500_));
 sky130_fd_sc_hd__xor2_4 _14911_ (.A(_12932_),
    .B(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__or2_4 _14912_ (.A(_04394_),
    .B(_04411_),
    .X(_04502_));
 sky130_fd_sc_hd__xnor2_4 _14913_ (.A(_12954_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__xnor2_1 _14914_ (.A(_04501_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__xnor2_1 _14915_ (.A(_04499_),
    .B(_04504_),
    .Y(_12110_));
 sky130_fd_sc_hd__maj3_1 _14916_ (.A(\hash.CA2.b_dash[4] ),
    .B(\hash.CA2.a_dash[4] ),
    .C(_04487_),
    .X(_04505_));
 sky130_fd_sc_hd__inv_1 _14917_ (.A(_04505_),
    .Y(_12121_));
 sky130_fd_sc_hd__clkinv_1 _14918_ (.A(_13251_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2b_2 _14919_ (.A(_12086_),
    .B_N(_13245_),
    .Y(_04507_));
 sky130_fd_sc_hd__o21ai_2 _14920_ (.A1(_13244_),
    .A2(_04507_),
    .B1(_13252_),
    .Y(_04508_));
 sky130_fd_sc_hd__a21boi_2 _14921_ (.A1(_04508_),
    .A2(_04506_),
    .B1_N(_13259_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _14922_ (.A(_04506_),
    .B(_04508_),
    .Y(_04510_));
 sky130_fd_sc_hd__nor2_2 _14923_ (.A(_13259_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_4 _14924_ (.A(net1057),
    .B(_04511_),
    .Y(_13260_));
 sky130_fd_sc_hd__clkinv_2 _14925_ (.A(_13260_),
    .Y(_12120_));
 sky130_fd_sc_hd__o2111ai_4 _14926_ (.A1(_04419_),
    .A2(_12965_),
    .B1(_12968_),
    .C1(_12970_),
    .D1(_12972_),
    .Y(_04512_));
 sky130_fd_sc_hd__a21o_1 _14927_ (.A1(_12968_),
    .A2(_12969_),
    .B1(_12967_),
    .X(_04513_));
 sky130_fd_sc_hd__nand2_1 _14928_ (.A(_12972_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__nand2_1 _14929_ (.A(_04512_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__nor2_2 _14930_ (.A(_12971_),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__xnor2_4 _14931_ (.A(_12976_),
    .B(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__o21ai_0 _14932_ (.A1(_04389_),
    .A2(_04436_),
    .B1(_04393_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21oi_2 _14933_ (.A1(_12954_),
    .A2(_04518_),
    .B1(_12953_),
    .Y(_04519_));
 sky130_fd_sc_hd__xnor2_4 _14934_ (.A(_12956_),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__o21ai_2 _14935_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04400_),
    .Y(_04521_));
 sky130_fd_sc_hd__xor2_4 _14936_ (.A(_12930_),
    .B(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__xor2_1 _14937_ (.A(_04520_),
    .B(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__xnor2_2 _14938_ (.A(_04517_),
    .B(_04523_),
    .Y(_12119_));
 sky130_fd_sc_hd__maj3_1 _14939_ (.A(\hash.CA2.b_dash[5] ),
    .B(\hash.CA2.a_dash[5] ),
    .C(_04501_),
    .X(_04524_));
 sky130_fd_sc_hd__inv_1 _14940_ (.A(_04524_),
    .Y(_12130_));
 sky130_fd_sc_hd__a211oi_2 _14941_ (.A1(_13239_),
    .A2(net1055),
    .B1(_13238_),
    .C1(_13244_),
    .Y(_04525_));
 sky130_fd_sc_hd__o211ai_1 _14942_ (.A1(_13245_),
    .A2(_13244_),
    .B1(_13259_),
    .C1(_13252_),
    .Y(_04526_));
 sky130_fd_sc_hd__a21oi_1 _14943_ (.A1(_13259_),
    .A2(_13251_),
    .B1(_13258_),
    .Y(_04527_));
 sky130_fd_sc_hd__o21ai_2 _14944_ (.A1(_04526_),
    .A2(_04525_),
    .B1(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__xor2_2 _14945_ (.A(_13266_),
    .B(_04528_),
    .X(_13267_));
 sky130_fd_sc_hd__clkinv_2 _14946_ (.A(_13267_),
    .Y(_12129_));
 sky130_fd_sc_hd__nor2_1 _14947_ (.A(_04492_),
    .B(_04498_),
    .Y(_04529_));
 sky130_fd_sc_hd__o21ai_2 _14948_ (.A1(_12971_),
    .A2(_04529_),
    .B1(_12976_),
    .Y(_04530_));
 sky130_fd_sc_hd__nor2_2 _14949_ (.A(_12974_),
    .B(_12975_),
    .Y(_04531_));
 sky130_fd_sc_hd__and3_1 _14950_ (.A(_12974_),
    .B(_12972_),
    .C(_12976_),
    .X(_04532_));
 sky130_fd_sc_hd__nand3_2 _14951_ (.A(_04496_),
    .B(_04497_),
    .C(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__nand2_2 _14952_ (.A(_12974_),
    .B(_12975_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand3_2 _14953_ (.A(_12974_),
    .B(_12976_),
    .C(_12971_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand3_2 _14954_ (.A(_04533_),
    .B(_04534_),
    .C(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__a21oi_4 _14955_ (.A1(_04530_),
    .A2(_04531_),
    .B1(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__nor2_1 _14956_ (.A(_04394_),
    .B(_04411_),
    .Y(_04538_));
 sky130_fd_sc_hd__a21o_1 _14957_ (.A1(_12954_),
    .A2(_04538_),
    .B1(_12953_),
    .X(_04539_));
 sky130_fd_sc_hd__a21oi_2 _14958_ (.A1(_12956_),
    .A2(_04539_),
    .B1(_12955_),
    .Y(_04540_));
 sky130_fd_sc_hd__xnor2_4 _14959_ (.A(_12958_),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__xnor2_4 _14960_ (.A(_12928_),
    .B(_04428_),
    .Y(_04542_));
 sky130_fd_sc_hd__inv_4 _14961_ (.A(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__xnor2_1 _14962_ (.A(_04541_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__xnor2_1 _14963_ (.A(_04537_),
    .B(_04544_),
    .Y(_12128_));
 sky130_fd_sc_hd__maj3_1 _14964_ (.A(\hash.CA2.b_dash[6] ),
    .B(\hash.CA2.a_dash[6] ),
    .C(_04522_),
    .X(_04545_));
 sky130_fd_sc_hd__inv_1 _14965_ (.A(_04545_),
    .Y(_12139_));
 sky130_fd_sc_hd__o21a_1 _14966_ (.A1(_04509_),
    .A2(_13258_),
    .B1(_13266_),
    .X(_04546_));
 sky130_fd_sc_hd__or2_1 _14967_ (.A(_13265_),
    .B(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__xor2_2 _14968_ (.A(_04547_),
    .B(_13273_),
    .X(_13274_));
 sky130_fd_sc_hd__clkinvlp_2 _14969_ (.A(_13274_),
    .Y(_12138_));
 sky130_fd_sc_hd__nor3_1 _14970_ (.A(_12971_),
    .B(_12973_),
    .C(_12975_),
    .Y(_04548_));
 sky130_fd_sc_hd__nand3_2 _14971_ (.A(_04514_),
    .B(_04512_),
    .C(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__nor3_1 _14972_ (.A(_12976_),
    .B(_12973_),
    .C(_12975_),
    .Y(_04550_));
 sky130_fd_sc_hd__nor2_1 _14973_ (.A(_12974_),
    .B(_12973_),
    .Y(_04551_));
 sky130_fd_sc_hd__nor2_2 _14974_ (.A(_04550_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_4 _14975_ (.A(net1090),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__xnor2_4 _14976_ (.A(_12978_),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__nor2_1 _14977_ (.A(_04455_),
    .B(_04483_),
    .Y(_04555_));
 sky130_fd_sc_hd__a22o_1 _14978_ (.A1(_12964_),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_04456_),
    .X(_04556_));
 sky130_fd_sc_hd__and2_4 _14979_ (.A(_04482_),
    .B(_04456_),
    .X(_04557_));
 sky130_fd_sc_hd__nor2_1 _14980_ (.A(_04556_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__o31a_1 _14981_ (.A1(_12964_),
    .A2(_04450_),
    .A3(_04555_),
    .B1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1411 ();
 sky130_fd_sc_hd__nand2_2 _14983_ (.A(_04397_),
    .B(net1089),
    .Y(_04561_));
 sky130_fd_sc_hd__xnor2_4 _14984_ (.A(_12940_),
    .B(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__xor2_1 _14985_ (.A(_04559_),
    .B(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__xnor2_2 _14986_ (.A(_04554_),
    .B(_04563_),
    .Y(_12137_));
 sky130_fd_sc_hd__maj3_1 _14987_ (.A(\hash.CA2.b_dash[7] ),
    .B(\hash.CA2.a_dash[7] ),
    .C(_04542_),
    .X(_04564_));
 sky130_fd_sc_hd__inv_1 _14988_ (.A(_04564_),
    .Y(_12148_));
 sky130_fd_sc_hd__clkinv_1 _14989_ (.A(_13272_),
    .Y(_04565_));
 sky130_fd_sc_hd__o21ai_0 _14990_ (.A1(_13266_),
    .A2(_13265_),
    .B1(_13273_),
    .Y(_04566_));
 sky130_fd_sc_hd__nand2_1 _14991_ (.A(_04565_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__o31ai_1 _14992_ (.A1(_13265_),
    .A2(_13272_),
    .A3(_04528_),
    .B1(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__xnor2_1 _14993_ (.A(_13280_),
    .B(_04568_),
    .Y(_13281_));
 sky130_fd_sc_hd__clkinvlp_4 _14994_ (.A(_13281_),
    .Y(_12147_));
 sky130_fd_sc_hd__o21ai_2 _14995_ (.A1(_12973_),
    .A2(_04536_),
    .B1(_12978_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_2 _14996_ (.A(_12980_),
    .B(_12977_),
    .Y(_04570_));
 sky130_fd_sc_hd__nor2_2 _14997_ (.A(_12973_),
    .B(_12977_),
    .Y(_04571_));
 sky130_fd_sc_hd__o21ai_2 _14998_ (.A1(_12978_),
    .A2(_12977_),
    .B1(_12980_),
    .Y(_04572_));
 sky130_fd_sc_hd__a41oi_4 _14999_ (.A1(_04533_),
    .A2(_04534_),
    .A3(_04535_),
    .A4(_04571_),
    .B1(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__a21o_4 _15000_ (.A1(_04569_),
    .A2(_04570_),
    .B1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__o21ai_0 _15001_ (.A1(_04502_),
    .A2(_04412_),
    .B1(_04383_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21o_4 _15002_ (.A1(_12964_),
    .A2(_04575_),
    .B1(_12963_),
    .X(_04576_));
 sky130_fd_sc_hd__xor2_4 _15003_ (.A(_12962_),
    .B(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__a21o_1 _15004_ (.A1(_12940_),
    .A2(_12927_),
    .B1(_12939_),
    .X(_04578_));
 sky130_fd_sc_hd__a41oi_2 _15005_ (.A1(_12928_),
    .A2(_12940_),
    .A3(_04422_),
    .A4(_04427_),
    .B1(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__xnor2_4 _15006_ (.A(_12938_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__xnor2_1 _15007_ (.A(_04577_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__xnor2_1 _15008_ (.A(_04574_),
    .B(_04581_),
    .Y(_12146_));
 sky130_fd_sc_hd__maj3_1 _15009_ (.A(\hash.CA2.b_dash[8] ),
    .B(\hash.CA2.a_dash[8] ),
    .C(_04562_),
    .X(_04582_));
 sky130_fd_sc_hd__inv_1 _15010_ (.A(_04582_),
    .Y(_12157_));
 sky130_fd_sc_hd__o21ai_2 _15011_ (.A1(_13265_),
    .A2(_04546_),
    .B1(_13273_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _15012_ (.A(_04565_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__a21o_1 _15013_ (.A1(_13280_),
    .A2(_04584_),
    .B1(_13279_),
    .X(_04585_));
 sky130_fd_sc_hd__xor2_2 _15014_ (.A(_13287_),
    .B(_04585_),
    .X(_13288_));
 sky130_fd_sc_hd__clkinv_2 _15015_ (.A(net1051),
    .Y(_12156_));
 sky130_fd_sc_hd__a31o_4 _15016_ (.A1(_04549_),
    .A2(_12978_),
    .A3(_04552_),
    .B1(_12977_),
    .X(_04586_));
 sky130_fd_sc_hd__a21oi_4 _15017_ (.A1(_12980_),
    .A2(_04586_),
    .B1(_12979_),
    .Y(_04587_));
 sky130_fd_sc_hd__xor2_4 _15018_ (.A(_04587_),
    .B(_12982_),
    .X(_04588_));
 sky130_fd_sc_hd__clkinv_1 _15019_ (.A(_12960_),
    .Y(_04589_));
 sky130_fd_sc_hd__nor3_1 _15020_ (.A(_04589_),
    .B(_12961_),
    .C(_12963_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_2 _15021_ (.A(_04558_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2b_4 _15022_ (.A(_12960_),
    .B_N(_12962_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_2 _15023_ (.A1(_04556_),
    .A2(_04557_),
    .B1(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__nor3_1 _15024_ (.A(_04589_),
    .B(_12962_),
    .C(_12961_),
    .Y(_04594_));
 sky130_fd_sc_hd__a221oi_2 _15025_ (.A1(_04589_),
    .A2(_12961_),
    .B1(_12963_),
    .B2(_04592_),
    .C1(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand3_4 _15026_ (.A(_04591_),
    .B(_04593_),
    .C(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__a31o_1 _15027_ (.A1(_12940_),
    .A2(_04397_),
    .A3(_04402_),
    .B1(_12939_),
    .X(_04597_));
 sky130_fd_sc_hd__a21oi_2 _15028_ (.A1(_12938_),
    .A2(_04597_),
    .B1(_12937_),
    .Y(_04598_));
 sky130_fd_sc_hd__xnor2_4 _15029_ (.A(_12942_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__xnor2_1 _15030_ (.A(_04596_),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__xnor2_2 _15031_ (.A(_04588_),
    .B(_04600_),
    .Y(_12155_));
 sky130_fd_sc_hd__maj3_1 _15032_ (.A(\hash.CA2.b_dash[9] ),
    .B(\hash.CA2.a_dash[9] ),
    .C(_04580_),
    .X(_04601_));
 sky130_fd_sc_hd__inv_1 _15033_ (.A(_04601_),
    .Y(_12166_));
 sky130_fd_sc_hd__nor2b_1 _15034_ (.A(_04568_),
    .B_N(_13280_),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_0 _15035_ (.A1(_13279_),
    .A2(_04602_),
    .B1(_13287_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand2b_2 _15036_ (.A_N(_13286_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__xor2_2 _15037_ (.A(_13294_),
    .B(_04604_),
    .X(_13295_));
 sky130_fd_sc_hd__inv_2 _15038_ (.A(_13295_),
    .Y(_12165_));
 sky130_fd_sc_hd__xor2_1 _15039_ (.A(\hash.CA2.p1[31] ),
    .B(\hash.CA2.p3[31] ),
    .X(_04605_));
 sky130_fd_sc_hd__or3_1 _15040_ (.A(_12979_),
    .B(_12981_),
    .C(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__nand2_1 _15041_ (.A(_12982_),
    .B(_04605_),
    .Y(_04607_));
 sky130_fd_sc_hd__mux2i_1 _15042_ (.A0(_04606_),
    .A1(_04607_),
    .S(_04573_),
    .Y(_04608_));
 sky130_fd_sc_hd__and2_0 _15043_ (.A(_12982_),
    .B(_12979_),
    .X(_04609_));
 sky130_fd_sc_hd__o21ai_0 _15044_ (.A1(_12981_),
    .A2(_04609_),
    .B1(_04605_),
    .Y(_04610_));
 sky130_fd_sc_hd__o31ai_2 _15045_ (.A1(_12982_),
    .A2(_12981_),
    .A3(_04605_),
    .B1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nor2_4 _15046_ (.A(_04611_),
    .B(_04608_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_2 _15047_ (.A(_04433_),
    .B(_04458_),
    .Y(_04613_));
 sky130_fd_sc_hd__xnor2_4 _15048_ (.A(_12944_),
    .B(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__xor2_1 _15049_ (.A(_04420_),
    .B(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__xnor2_1 _15050_ (.A(_04612_),
    .B(_04615_),
    .Y(_12164_));
 sky130_fd_sc_hd__maj3_1 _15051_ (.A(\hash.CA2.b_dash[10] ),
    .B(\hash.CA2.a_dash[10] ),
    .C(_04599_),
    .X(_04616_));
 sky130_fd_sc_hd__inv_1 _15052_ (.A(_04616_),
    .Y(_12175_));
 sky130_fd_sc_hd__and3_1 _15053_ (.A(_13280_),
    .B(_13287_),
    .C(_13294_),
    .X(_04617_));
 sky130_fd_sc_hd__a21boi_2 _15054_ (.A1(_04565_),
    .A2(_04583_),
    .B1_N(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__a21oi_1 _15055_ (.A1(_13287_),
    .A2(_13279_),
    .B1(_13286_),
    .Y(_04619_));
 sky130_fd_sc_hd__nor2b_2 _15056_ (.A(_04619_),
    .B_N(_13294_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _15057_ (.A(_13293_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__nand2b_1 _15058_ (.A_N(_04618_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__xor2_1 _15059_ (.A(_13301_),
    .B(_04622_),
    .X(_13302_));
 sky130_fd_sc_hd__clkinvlp_2 _15060_ (.A(_13302_),
    .Y(_12174_));
 sky130_fd_sc_hd__xnor2_2 _15061_ (.A(_12948_),
    .B(_04472_),
    .Y(_04623_));
 sky130_fd_sc_hd__xnor2_1 _15062_ (.A(_12922_),
    .B(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__xor2_1 _15063_ (.A(_04467_),
    .B(_04624_),
    .X(_12173_));
 sky130_fd_sc_hd__maj3_1 _15064_ (.A(\hash.CA2.b_dash[11] ),
    .B(\hash.CA2.a_dash[11] ),
    .C(_04614_),
    .X(_04625_));
 sky130_fd_sc_hd__inv_1 _15065_ (.A(_04625_),
    .Y(_12184_));
 sky130_fd_sc_hd__o311ai_2 _15066_ (.A1(_04528_),
    .A2(_13272_),
    .A3(_13265_),
    .B1(_04567_),
    .C1(_04617_),
    .Y(_04626_));
 sky130_fd_sc_hd__a21boi_2 _15067_ (.A1(_04626_),
    .A2(_04621_),
    .B1_N(_13301_),
    .Y(_04627_));
 sky130_fd_sc_hd__nor2_1 _15068_ (.A(_13300_),
    .B(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__xnor2_2 _15069_ (.A(_13308_),
    .B(_04628_),
    .Y(_13309_));
 sky130_fd_sc_hd__clkinv_4 _15070_ (.A(_13309_),
    .Y(_12183_));
 sky130_fd_sc_hd__xnor2_1 _15071_ (.A(_12082_),
    .B(_04437_),
    .Y(_04629_));
 sky130_fd_sc_hd__xnor2_1 _15072_ (.A(net1114),
    .B(_04629_),
    .Y(_12182_));
 sky130_fd_sc_hd__maj3_1 _15073_ (.A(\hash.CA2.b_dash[12] ),
    .B(\hash.CA2.a_dash[12] ),
    .C(_04623_),
    .X(_04630_));
 sky130_fd_sc_hd__inv_1 _15074_ (.A(_04630_),
    .Y(_12193_));
 sky130_fd_sc_hd__or3_1 _15075_ (.A(_13293_),
    .B(_13300_),
    .C(_13307_),
    .X(_04631_));
 sky130_fd_sc_hd__nor3_1 _15076_ (.A(_13301_),
    .B(_13300_),
    .C(_13307_),
    .Y(_04632_));
 sky130_fd_sc_hd__nor2_1 _15077_ (.A(_13308_),
    .B(_13307_),
    .Y(_04633_));
 sky130_fd_sc_hd__nor2_1 _15078_ (.A(_04632_),
    .B(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__o31ai_4 _15079_ (.A1(_04620_),
    .A2(_04631_),
    .A3(_04618_),
    .B1(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__xnor2_2 _15080_ (.A(_13315_),
    .B(net1103),
    .Y(_13316_));
 sky130_fd_sc_hd__clkinvlp_4 _15081_ (.A(net1104),
    .Y(_12192_));
 sky130_fd_sc_hd__xor2_1 _15082_ (.A(_12952_),
    .B(_04474_),
    .X(_04636_));
 sky130_fd_sc_hd__xnor2_1 _15083_ (.A(_04421_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__xnor2_1 _15084_ (.A(_04499_),
    .B(_04637_),
    .Y(_12191_));
 sky130_fd_sc_hd__nor2_4 _15085_ (.A(\hash.CA2.a_dash[13] ),
    .B(_04437_),
    .Y(_04638_));
 sky130_fd_sc_hd__a21oi_1 _15086_ (.A1(\hash.CA2.a_dash[13] ),
    .A2(_04437_),
    .B1(\hash.CA2.b_dash[13] ),
    .Y(_04639_));
 sky130_fd_sc_hd__nor2_1 _15087_ (.A(_04638_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__inv_1 _15088_ (.A(_04640_),
    .Y(_12202_));
 sky130_fd_sc_hd__clkinv_1 _15089_ (.A(_13322_),
    .Y(_04641_));
 sky130_fd_sc_hd__o21ai_1 _15090_ (.A1(_13300_),
    .A2(_04627_),
    .B1(_13308_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand2b_1 _15091_ (.A_N(_13307_),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__a21o_1 _15092_ (.A1(_13315_),
    .A2(_04643_),
    .B1(_13314_),
    .X(_04644_));
 sky130_fd_sc_hd__xnor2_2 _15093_ (.A(_04641_),
    .B(_04644_),
    .Y(_13323_));
 sky130_fd_sc_hd__inv_4 _15094_ (.A(_13323_),
    .Y(_12201_));
 sky130_fd_sc_hd__xor2_1 _15095_ (.A(_04470_),
    .B(_04484_),
    .X(_04645_));
 sky130_fd_sc_hd__xnor2_1 _15096_ (.A(_04517_),
    .B(_04645_),
    .Y(_12200_));
 sky130_fd_sc_hd__nor2_1 _15097_ (.A(\hash.CA2.a_dash[14] ),
    .B(_04636_),
    .Y(_04646_));
 sky130_fd_sc_hd__a21oi_1 _15098_ (.A1(\hash.CA2.a_dash[14] ),
    .A2(_04636_),
    .B1(\hash.CA2.b_dash[14] ),
    .Y(_04647_));
 sky130_fd_sc_hd__nor2_1 _15099_ (.A(_04646_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__clkinv_1 _15100_ (.A(_04648_),
    .Y(_12211_));
 sky130_fd_sc_hd__inv_1 _15101_ (.A(_13315_),
    .Y(_04649_));
 sky130_fd_sc_hd__nor2_1 _15102_ (.A(_04649_),
    .B(_04641_),
    .Y(_04650_));
 sky130_fd_sc_hd__nand2_1 _15103_ (.A(_13329_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__and3_1 _15104_ (.A(_13322_),
    .B(_13329_),
    .C(_13314_),
    .X(_04652_));
 sky130_fd_sc_hd__a21oi_1 _15105_ (.A1(_13329_),
    .A2(_13321_),
    .B1(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__o21ai_4 _15106_ (.A1(_04635_),
    .A2(_04651_),
    .B1(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__o21bai_1 _15107_ (.A1(_04649_),
    .A2(_04635_),
    .B1_N(_13314_),
    .Y(_04655_));
 sky130_fd_sc_hd__a211oi_2 _15108_ (.A1(_13322_),
    .A2(_04655_),
    .B1(_13321_),
    .C1(_13329_),
    .Y(_04656_));
 sky130_fd_sc_hd__nor2_2 _15109_ (.A(net1074),
    .B(_04656_),
    .Y(_13330_));
 sky130_fd_sc_hd__clkinv_2 _15110_ (.A(net1067),
    .Y(_12210_));
 sky130_fd_sc_hd__xor2_1 _15111_ (.A(_04487_),
    .B(_04503_),
    .X(_04657_));
 sky130_fd_sc_hd__xnor2_1 _15112_ (.A(_04537_),
    .B(_04657_),
    .Y(_12209_));
 sky130_fd_sc_hd__maj3_1 _15113_ (.A(\hash.CA2.b_dash[15] ),
    .B(\hash.CA2.a_dash[15] ),
    .C(_04484_),
    .X(_04658_));
 sky130_fd_sc_hd__inv_1 _15114_ (.A(_04658_),
    .Y(_12220_));
 sky130_fd_sc_hd__a211oi_2 _15115_ (.A1(_04644_),
    .A2(_13322_),
    .B1(_13328_),
    .C1(_13321_),
    .Y(_04659_));
 sky130_fd_sc_hd__nor2_1 _15116_ (.A(_13329_),
    .B(_13328_),
    .Y(_04660_));
 sky130_fd_sc_hd__nor2_2 _15117_ (.A(_04659_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__xor2_1 _15118_ (.A(_13336_),
    .B(_04661_),
    .X(_13337_));
 sky130_fd_sc_hd__clkinvlp_2 _15119_ (.A(_13337_),
    .Y(_12219_));
 sky130_fd_sc_hd__xor2_2 _15120_ (.A(_12978_),
    .B(_04553_),
    .X(_04662_));
 sky130_fd_sc_hd__xnor2_1 _15121_ (.A(_04501_),
    .B(_04520_),
    .Y(_04663_));
 sky130_fd_sc_hd__xnor2_1 _15122_ (.A(_04662_),
    .B(_04663_),
    .Y(_12218_));
 sky130_fd_sc_hd__maj3_1 _15123_ (.A(\hash.CA2.b_dash[16] ),
    .B(\hash.CA2.a_dash[16] ),
    .C(_04503_),
    .X(_04664_));
 sky130_fd_sc_hd__inv_1 _15124_ (.A(_04664_),
    .Y(_12229_));
 sky130_fd_sc_hd__o21ai_1 _15125_ (.A1(_13328_),
    .A2(net1074),
    .B1(_13336_),
    .Y(_04665_));
 sky130_fd_sc_hd__nand2b_2 _15126_ (.A_N(_13335_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__xor2_4 _15127_ (.A(_13343_),
    .B(_04666_),
    .X(_13344_));
 sky130_fd_sc_hd__inv_2 _15128_ (.A(_13344_),
    .Y(_12228_));
 sky130_fd_sc_hd__xnor2_1 _15129_ (.A(_04522_),
    .B(_04541_),
    .Y(_04667_));
 sky130_fd_sc_hd__xnor2_1 _15130_ (.A(_04574_),
    .B(_04667_),
    .Y(_12227_));
 sky130_fd_sc_hd__maj3_1 _15131_ (.A(\hash.CA2.b_dash[17] ),
    .B(\hash.CA2.a_dash[17] ),
    .C(_04520_),
    .X(_04668_));
 sky130_fd_sc_hd__inv_1 _15132_ (.A(_04668_),
    .Y(_12238_));
 sky130_fd_sc_hd__a21o_1 _15133_ (.A1(_13336_),
    .A2(_04661_),
    .B1(_13335_),
    .X(_04669_));
 sky130_fd_sc_hd__a21o_1 _15134_ (.A1(_13343_),
    .A2(_04669_),
    .B1(_13342_),
    .X(_04670_));
 sky130_fd_sc_hd__xor2_2 _15135_ (.A(_13350_),
    .B(_04670_),
    .X(_13351_));
 sky130_fd_sc_hd__inv_2 _15136_ (.A(_13351_),
    .Y(_12237_));
 sky130_fd_sc_hd__xnor2_1 _15137_ (.A(_04542_),
    .B(_04559_),
    .Y(_04671_));
 sky130_fd_sc_hd__xnor2_1 _15138_ (.A(net1113),
    .B(_04671_),
    .Y(_12236_));
 sky130_fd_sc_hd__nor2_2 _15139_ (.A(\hash.CA2.a_dash[18] ),
    .B(_04541_),
    .Y(_04672_));
 sky130_fd_sc_hd__a21oi_1 _15140_ (.A1(\hash.CA2.a_dash[18] ),
    .A2(_04541_),
    .B1(\hash.CA2.b_dash[18] ),
    .Y(_04673_));
 sky130_fd_sc_hd__nor2_1 _15141_ (.A(_04672_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__inv_2 _15142_ (.A(_04674_),
    .Y(_12247_));
 sky130_fd_sc_hd__a21o_1 _15143_ (.A1(_13336_),
    .A2(_13328_),
    .B1(_13335_),
    .X(_04675_));
 sky130_fd_sc_hd__a21o_1 _15144_ (.A1(_13343_),
    .A2(_04675_),
    .B1(_13342_),
    .X(_04676_));
 sky130_fd_sc_hd__a21oi_1 _15145_ (.A1(_13350_),
    .A2(_04676_),
    .B1(_13349_),
    .Y(_04677_));
 sky130_fd_sc_hd__and3_4 _15146_ (.A(_13336_),
    .B(_13343_),
    .C(_13350_),
    .X(_04678_));
 sky130_fd_sc_hd__nand2_1 _15147_ (.A(net1074),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__nand2_1 _15148_ (.A(_04677_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__xor2_1 _15149_ (.A(_13357_),
    .B(_04680_),
    .X(_13358_));
 sky130_fd_sc_hd__inv_2 _15150_ (.A(_13358_),
    .Y(_12246_));
 sky130_fd_sc_hd__xnor2_2 _15151_ (.A(_12962_),
    .B(_04576_),
    .Y(_04681_));
 sky130_fd_sc_hd__xnor2_1 _15152_ (.A(_04562_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__xnor2_1 _15153_ (.A(_04612_),
    .B(_04682_),
    .Y(_12245_));
 sky130_fd_sc_hd__maj3_1 _15154_ (.A(\hash.CA2.b_dash[19] ),
    .B(\hash.CA2.a_dash[19] ),
    .C(_04559_),
    .X(_04683_));
 sky130_fd_sc_hd__inv_1 _15155_ (.A(_04683_),
    .Y(_12256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1410 ();
 sky130_fd_sc_hd__a21o_1 _15157_ (.A1(_13343_),
    .A2(_13335_),
    .B1(_13342_),
    .X(_04685_));
 sky130_fd_sc_hd__a21o_1 _15158_ (.A1(_13350_),
    .A2(_04685_),
    .B1(_13349_),
    .X(_04686_));
 sky130_fd_sc_hd__a21o_1 _15159_ (.A1(_13357_),
    .A2(_04686_),
    .B1(_13356_),
    .X(_04687_));
 sky130_fd_sc_hd__a31oi_2 _15160_ (.A1(_13357_),
    .A2(_04678_),
    .A3(_04661_),
    .B1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__xnor2_1 _15161_ (.A(_13364_),
    .B(_04688_),
    .Y(_13365_));
 sky130_fd_sc_hd__clkinvlp_2 _15162_ (.A(_13365_),
    .Y(_12255_));
 sky130_fd_sc_hd__xnor2_1 _15163_ (.A(_12922_),
    .B(_04580_),
    .Y(_04689_));
 sky130_fd_sc_hd__xor2_1 _15164_ (.A(_04596_),
    .B(_04689_),
    .X(_12254_));
 sky130_fd_sc_hd__maj3_1 _15165_ (.A(\hash.CA2.b_dash[20] ),
    .B(\hash.CA2.a_dash[20] ),
    .C(_04577_),
    .X(_04690_));
 sky130_fd_sc_hd__inv_1 _15166_ (.A(_04690_),
    .Y(_12265_));
 sky130_fd_sc_hd__nand2_1 _15167_ (.A(_13357_),
    .B(_13364_),
    .Y(_04691_));
 sky130_fd_sc_hd__nand2_1 _15168_ (.A(_13364_),
    .B(_13356_),
    .Y(_04692_));
 sky130_fd_sc_hd__o21ai_0 _15169_ (.A1(_04677_),
    .A2(_04691_),
    .B1(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__a41oi_2 _15170_ (.A1(_13357_),
    .A2(_04654_),
    .A3(_13364_),
    .A4(_04678_),
    .B1(_04693_),
    .Y(_04694_));
 sky130_fd_sc_hd__nor2b_1 _15171_ (.A(_13363_),
    .B_N(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__xnor2_1 _15172_ (.A(_13371_),
    .B(_04695_),
    .Y(_13372_));
 sky130_fd_sc_hd__inv_2 _15173_ (.A(_13372_),
    .Y(_12264_));
 sky130_fd_sc_hd__xnor2_1 _15174_ (.A(_12082_),
    .B(_04599_),
    .Y(_04696_));
 sky130_fd_sc_hd__xor2_1 _15175_ (.A(_04420_),
    .B(_04696_),
    .X(_12263_));
 sky130_fd_sc_hd__nor2_2 _15176_ (.A(\hash.CA2.a_dash[21] ),
    .B(_04596_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21oi_1 _15177_ (.A1(\hash.CA2.a_dash[21] ),
    .A2(_04596_),
    .B1(\hash.CA2.b_dash[21] ),
    .Y(_04698_));
 sky130_fd_sc_hd__nor2_1 _15178_ (.A(_04697_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__inv_1 _15179_ (.A(_04699_),
    .Y(_12274_));
 sky130_fd_sc_hd__inv_1 _15180_ (.A(_13364_),
    .Y(_04700_));
 sky130_fd_sc_hd__o21bai_1 _15181_ (.A1(_04700_),
    .A2(_04688_),
    .B1_N(_13363_),
    .Y(_04701_));
 sky130_fd_sc_hd__a21oi_2 _15182_ (.A1(_04701_),
    .A2(_13371_),
    .B1(_13370_),
    .Y(_04702_));
 sky130_fd_sc_hd__xnor2_2 _15183_ (.A(_13378_),
    .B(_04702_),
    .Y(_13379_));
 sky130_fd_sc_hd__inv_4 _15184_ (.A(net1078),
    .Y(_12273_));
 sky130_fd_sc_hd__xor2_1 _15185_ (.A(_04421_),
    .B(_04614_),
    .X(_04703_));
 sky130_fd_sc_hd__xnor2_1 _15186_ (.A(_04467_),
    .B(_04703_),
    .Y(_12272_));
 sky130_fd_sc_hd__nand2_2 _15187_ (.A(\hash.CA2.a_dash[22] ),
    .B(_04420_),
    .Y(_04704_));
 sky130_fd_sc_hd__o21ai_0 _15188_ (.A1(\hash.CA2.a_dash[22] ),
    .A2(_04420_),
    .B1(\hash.CA2.b_dash[22] ),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_1 _15189_ (.A(_04704_),
    .B(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__inv_1 _15190_ (.A(_04706_),
    .Y(_12283_));
 sky130_fd_sc_hd__nor3_1 _15191_ (.A(_13363_),
    .B(_13370_),
    .C(_13377_),
    .Y(_04707_));
 sky130_fd_sc_hd__or2_0 _15192_ (.A(_13371_),
    .B(_13370_),
    .X(_04708_));
 sky130_fd_sc_hd__a21oi_1 _15193_ (.A1(_13378_),
    .A2(_04708_),
    .B1(_13377_),
    .Y(_04709_));
 sky130_fd_sc_hd__a21oi_2 _15194_ (.A1(_04694_),
    .A2(_04707_),
    .B1(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__xor2_2 _15195_ (.A(_13385_),
    .B(net1068),
    .X(_13386_));
 sky130_fd_sc_hd__clkinv_2 _15196_ (.A(_13386_),
    .Y(_12282_));
 sky130_fd_sc_hd__xnor2_1 _15197_ (.A(_04470_),
    .B(_04623_),
    .Y(_04711_));
 sky130_fd_sc_hd__xnor2_1 _15198_ (.A(_04481_),
    .B(_04711_),
    .Y(_12281_));
 sky130_fd_sc_hd__maj3_1 _15199_ (.A(\hash.CA2.b_dash[23] ),
    .B(\hash.CA2.a_dash[23] ),
    .C(_04467_),
    .X(_04712_));
 sky130_fd_sc_hd__inv_1 _15200_ (.A(_04712_),
    .Y(_12292_));
 sky130_fd_sc_hd__a211o_1 _15201_ (.A1(_13364_),
    .A2(_04687_),
    .B1(_13370_),
    .C1(_13363_),
    .X(_04713_));
 sky130_fd_sc_hd__and3_1 _15202_ (.A(_13378_),
    .B(_13385_),
    .C(_04708_),
    .X(_04714_));
 sky130_fd_sc_hd__a221oi_1 _15203_ (.A1(_13385_),
    .A2(_13377_),
    .B1(_04713_),
    .B2(_04714_),
    .C1(_13384_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand4_1 _15204_ (.A(_13364_),
    .B(_13371_),
    .C(_13378_),
    .D(_13385_),
    .Y(_04716_));
 sky130_fd_sc_hd__nor2_1 _15205_ (.A(_04660_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__and3_4 _15206_ (.A(_13357_),
    .B(_04678_),
    .C(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__o2111ai_1 _15207_ (.A1(_13300_),
    .A2(_04627_),
    .B1(_04650_),
    .C1(_04718_),
    .D1(_13308_),
    .Y(_04719_));
 sky130_fd_sc_hd__a21oi_1 _15208_ (.A1(_13315_),
    .A2(_13307_),
    .B1(_13314_),
    .Y(_04720_));
 sky130_fd_sc_hd__nor2_1 _15209_ (.A(_04641_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__o31ai_1 _15210_ (.A1(_13321_),
    .A2(_13328_),
    .A3(_04721_),
    .B1(_04718_),
    .Y(_04722_));
 sky130_fd_sc_hd__and3_4 _15211_ (.A(_04715_),
    .B(_04719_),
    .C(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__xnor2_2 _15212_ (.A(_13392_),
    .B(_04723_),
    .Y(_13393_));
 sky130_fd_sc_hd__clkinvlp_4 _15213_ (.A(_13393_),
    .Y(_12291_));
 sky130_fd_sc_hd__xnor2_1 _15214_ (.A(_04437_),
    .B(_04487_),
    .Y(_04724_));
 sky130_fd_sc_hd__xnor2_1 _15215_ (.A(_04499_),
    .B(_04724_),
    .Y(_12290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1409 ();
 sky130_fd_sc_hd__xnor2_2 _15217_ (.A(_12968_),
    .B(_04480_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_2 _15218_ (.A(\hash.CA2.a_dash[24] ),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__o21ai_0 _15219_ (.A1(\hash.CA2.a_dash[24] ),
    .A2(_04726_),
    .B1(\hash.CA2.b_dash[24] ),
    .Y(_04728_));
 sky130_fd_sc_hd__nand2_1 _15220_ (.A(_04727_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__inv_1 _15221_ (.A(_04729_),
    .Y(_12301_));
 sky130_fd_sc_hd__a21o_1 _15222_ (.A1(_13385_),
    .A2(_04710_),
    .B1(_13384_),
    .X(_04730_));
 sky130_fd_sc_hd__a21oi_1 _15223_ (.A1(_13392_),
    .A2(_04730_),
    .B1(_13391_),
    .Y(_04731_));
 sky130_fd_sc_hd__xnor2_1 _15224_ (.A(_13399_),
    .B(_04731_),
    .Y(_13400_));
 sky130_fd_sc_hd__clkinv_2 _15225_ (.A(_13400_),
    .Y(_12300_));
 sky130_fd_sc_hd__xnor2_1 _15226_ (.A(net1092),
    .B(_04501_),
    .Y(_04732_));
 sky130_fd_sc_hd__xnor2_1 _15227_ (.A(_04517_),
    .B(_04732_),
    .Y(_12299_));
 sky130_fd_sc_hd__inv_8 _15228_ (.A(\hash.CA2.b_dash[25] ),
    .Y(_04733_));
 sky130_fd_sc_hd__inv_2 _15229_ (.A(\hash.CA2.a_dash[25] ),
    .Y(_04734_));
 sky130_fd_sc_hd__maj3_1 _15230_ (.A(_04733_),
    .B(_04734_),
    .C(_04499_),
    .X(_12310_));
 sky130_fd_sc_hd__a21o_1 _15231_ (.A1(_13399_),
    .A2(_13391_),
    .B1(_13398_),
    .X(_04735_));
 sky130_fd_sc_hd__nand2_1 _15232_ (.A(_13392_),
    .B(_13399_),
    .Y(_04736_));
 sky130_fd_sc_hd__nor2_1 _15233_ (.A(_04723_),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__nor2_1 _15234_ (.A(_04735_),
    .B(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__xnor2_2 _15235_ (.A(_13406_),
    .B(_04738_),
    .Y(_13407_));
 sky130_fd_sc_hd__inv_4 _15236_ (.A(_13407_),
    .Y(_12309_));
 sky130_fd_sc_hd__xor2_1 _15237_ (.A(_04484_),
    .B(_04522_),
    .X(_04739_));
 sky130_fd_sc_hd__xnor2_1 _15238_ (.A(_04537_),
    .B(_04739_),
    .Y(_12308_));
 sky130_fd_sc_hd__maj3_1 _15239_ (.A(\hash.CA2.b_dash[26] ),
    .B(\hash.CA2.a_dash[26] ),
    .C(_04517_),
    .X(_04740_));
 sky130_fd_sc_hd__inv_1 _15240_ (.A(_04740_),
    .Y(_12319_));
 sky130_fd_sc_hd__nand2_1 _15241_ (.A(_13385_),
    .B(_13406_),
    .Y(_04741_));
 sky130_fd_sc_hd__nor2_1 _15242_ (.A(_04736_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_1 _15243_ (.A(_13406_),
    .B(_13384_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _15244_ (.A(_13406_),
    .B(_04735_),
    .Y(_04744_));
 sky130_fd_sc_hd__o21ai_0 _15245_ (.A1(_04736_),
    .A2(_04743_),
    .B1(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__a211o_4 _15246_ (.A1(_04742_),
    .A2(net1084),
    .B1(_04745_),
    .C1(_13405_),
    .X(_04746_));
 sky130_fd_sc_hd__xor2_4 _15247_ (.A(_04746_),
    .B(_13413_),
    .X(_13414_));
 sky130_fd_sc_hd__clkinv_4 _15248_ (.A(net1082),
    .Y(_12318_));
 sky130_fd_sc_hd__xnor2_1 _15249_ (.A(_04503_),
    .B(_04542_),
    .Y(_04747_));
 sky130_fd_sc_hd__xnor2_1 _15250_ (.A(_04662_),
    .B(_04747_),
    .Y(_12317_));
 sky130_fd_sc_hd__maj3_1 _15251_ (.A(\hash.CA2.b_dash[27] ),
    .B(\hash.CA2.a_dash[27] ),
    .C(_04537_),
    .X(_04748_));
 sky130_fd_sc_hd__inv_1 _15252_ (.A(_04748_),
    .Y(_12328_));
 sky130_fd_sc_hd__nand4_1 _15253_ (.A(_13392_),
    .B(_13399_),
    .C(_13406_),
    .D(_13413_),
    .Y(_04749_));
 sky130_fd_sc_hd__inv_1 _15254_ (.A(_04744_),
    .Y(_04750_));
 sky130_fd_sc_hd__o21ai_0 _15255_ (.A1(_13405_),
    .A2(_04750_),
    .B1(_13413_),
    .Y(_04751_));
 sky130_fd_sc_hd__o21ai_1 _15256_ (.A1(_04723_),
    .A2(_04749_),
    .B1(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nor2_1 _15257_ (.A(_13412_),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__xnor2_1 _15258_ (.A(_13420_),
    .B(_04753_),
    .Y(_13421_));
 sky130_fd_sc_hd__clkinv_2 _15259_ (.A(_13421_),
    .Y(_12327_));
 sky130_fd_sc_hd__a21oi_4 _15260_ (.A1(_04569_),
    .A2(_04570_),
    .B1(_04573_),
    .Y(_04754_));
 sky130_fd_sc_hd__xor2_1 _15261_ (.A(_04520_),
    .B(_04562_),
    .X(_04755_));
 sky130_fd_sc_hd__xnor2_1 _15262_ (.A(_04754_),
    .B(_04755_),
    .Y(_12326_));
 sky130_fd_sc_hd__nand2_1 _15263_ (.A(\hash.CA2.a_dash[28] ),
    .B(_04554_),
    .Y(_04756_));
 sky130_fd_sc_hd__o21ai_0 _15264_ (.A1(\hash.CA2.a_dash[28] ),
    .A2(_04554_),
    .B1(\hash.CA2.b_dash[28] ),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _15265_ (.A(_04756_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__inv_1 _15266_ (.A(_04758_),
    .Y(_12337_));
 sky130_fd_sc_hd__a21o_1 _15267_ (.A1(_13413_),
    .A2(_04746_),
    .B1(_13412_),
    .X(_04759_));
 sky130_fd_sc_hd__a21oi_2 _15268_ (.A1(_13420_),
    .A2(_04759_),
    .B1(_13419_),
    .Y(_04760_));
 sky130_fd_sc_hd__xor2_2 _15269_ (.A(_13427_),
    .B(_04760_),
    .X(_12336_));
 sky130_fd_sc_hd__xnor2_1 _15270_ (.A(_04541_),
    .B(_04580_),
    .Y(_04761_));
 sky130_fd_sc_hd__xnor2_1 _15271_ (.A(net1113),
    .B(_04761_),
    .Y(_12335_));
 sky130_fd_sc_hd__nor2_2 _15272_ (.A(\hash.CA2.a_dash[29] ),
    .B(_04754_),
    .Y(_04762_));
 sky130_fd_sc_hd__a21oi_1 _15273_ (.A1(\hash.CA2.a_dash[29] ),
    .A2(_04754_),
    .B1(\hash.CA2.b_dash[29] ),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2_1 _15274_ (.A(_04762_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__inv_1 _15275_ (.A(_04764_),
    .Y(_12346_));
 sky130_fd_sc_hd__inv_1 _15276_ (.A(_13420_),
    .Y(_04765_));
 sky130_fd_sc_hd__o21bai_1 _15277_ (.A1(_04765_),
    .A2(_04753_),
    .B1_N(_13419_),
    .Y(_04766_));
 sky130_fd_sc_hd__a21oi_1 _15278_ (.A1(_13427_),
    .A2(_04766_),
    .B1(_13426_),
    .Y(_04767_));
 sky130_fd_sc_hd__xnor2_2 _15279_ (.A(_13434_),
    .B(_04767_),
    .Y(_13435_));
 sky130_fd_sc_hd__inv_4 _15280_ (.A(_13435_),
    .Y(_12345_));
 sky130_fd_sc_hd__xor2_1 _15281_ (.A(_04559_),
    .B(_04599_),
    .X(_04768_));
 sky130_fd_sc_hd__xnor2_1 _15282_ (.A(_04612_),
    .B(_04768_),
    .Y(_12344_));
 sky130_fd_sc_hd__inv_2 _15283_ (.A(\hash.CA2.a_dash[30] ),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_1 _15284_ (.A(_04769_),
    .B(_04588_),
    .Y(_04770_));
 sky130_fd_sc_hd__nor2_1 _15285_ (.A(_04769_),
    .B(_04588_),
    .Y(_04771_));
 sky130_fd_sc_hd__a21oi_2 _15286_ (.A1(\hash.CA2.b_dash[30] ),
    .A2(_04770_),
    .B1(_04771_),
    .Y(_12355_));
 sky130_fd_sc_hd__nand2_1 _15287_ (.A(_13413_),
    .B(_04746_),
    .Y(_04772_));
 sky130_fd_sc_hd__a21oi_1 _15288_ (.A1(_13427_),
    .A2(_13419_),
    .B1(_13426_),
    .Y(_04773_));
 sky130_fd_sc_hd__nor2b_2 _15289_ (.A(_04773_),
    .B_N(_13434_),
    .Y(_04774_));
 sky130_fd_sc_hd__nor3_2 _15290_ (.A(_13412_),
    .B(_13433_),
    .C(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__a311o_1 _15291_ (.A1(_13420_),
    .A2(_13427_),
    .A3(_13434_),
    .B1(_13433_),
    .C1(_04774_),
    .X(_04776_));
 sky130_fd_sc_hd__a21boi_2 _15292_ (.A1(_04772_),
    .A2(_04775_),
    .B1_N(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__xnor2_2 _15293_ (.A(_13441_),
    .B(_04777_),
    .Y(_12354_));
 sky130_fd_sc_hd__xnor2_1 _15294_ (.A(_12922_),
    .B(_04614_),
    .Y(_04778_));
 sky130_fd_sc_hd__xnor2_1 _15295_ (.A(_04681_),
    .B(_04778_),
    .Y(_12353_));
 sky130_fd_sc_hd__nor2_4 _15296_ (.A(net353),
    .B(_13445_),
    .Y(_00781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1408 ();
 sky130_fd_sc_hd__or2_0 _15298_ (.A(\hash.reset ),
    .B(\hash.CA2.S1.X[2] ),
    .X(\hash.CA1.f[2] ));
 sky130_fd_sc_hd__clkinvlp_2 _15299_ (.A(\hash.CA1.f[2] ),
    .Y(_00813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1404 ();
 sky130_fd_sc_hd__nor2_4 _15304_ (.A(net355),
    .B(\hash.CA2.S1.X[3] ),
    .Y(_13851_));
 sky130_fd_sc_hd__nor2b_4 _15305_ (.A(net1043),
    .B_N(_13528_),
    .Y(_04784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1403 ();
 sky130_fd_sc_hd__nand2_8 _15307_ (.A(_09735_),
    .B(_04784_),
    .Y(_04786_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1400 ();
 sky130_fd_sc_hd__mux2i_4 _15311_ (.A0(_12986_),
    .A1(\w[62][0] ),
    .S(net362),
    .Y(_04790_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1398 ();
 sky130_fd_sc_hd__nand2_1 _15314_ (.A(net245),
    .B(_04786_),
    .Y(_04793_));
 sky130_fd_sc_hd__o21ai_0 _15315_ (.A1(_04786_),
    .A2(_04790_),
    .B1(_04793_),
    .Y(_00129_));
 sky130_fd_sc_hd__mux2i_4 _15316_ (.A0(_12989_),
    .A1(\w[62][1] ),
    .S(net362),
    .Y(_04794_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1397 ();
 sky130_fd_sc_hd__nand2_1 _15318_ (.A(net234),
    .B(_04786_),
    .Y(_04796_));
 sky130_fd_sc_hd__o21ai_0 _15319_ (.A1(_04786_),
    .A2(_04794_),
    .B1(_04796_),
    .Y(_00140_));
 sky130_fd_sc_hd__clkinv_16 _15320_ (.A(net364),
    .Y(_04797_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1395 ();
 sky130_fd_sc_hd__nand2_4 _15323_ (.A(_11602_),
    .B(net348),
    .Y(_04800_));
 sky130_fd_sc_hd__o21ai_4 _15324_ (.A1(\w[62][2] ),
    .A2(net348),
    .B1(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1394 ();
 sky130_fd_sc_hd__nand2_1 _15326_ (.A(net222),
    .B(_04786_),
    .Y(_04803_));
 sky130_fd_sc_hd__o21ai_0 _15327_ (.A1(_04786_),
    .A2(_04801_),
    .B1(_04803_),
    .Y(_00151_));
 sky130_fd_sc_hd__nor2b_1 _15328_ (.A(_12997_),
    .B_N(_11601_),
    .Y(_04804_));
 sky130_fd_sc_hd__nor2b_2 _15329_ (.A(_11601_),
    .B_N(_12997_),
    .Y(_04805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1393 ();
 sky130_fd_sc_hd__o21ai_2 _15331_ (.A1(_04804_),
    .A2(_04805_),
    .B1(net348),
    .Y(_04807_));
 sky130_fd_sc_hd__o21ai_4 _15332_ (.A1(\w[62][3] ),
    .A2(net348),
    .B1(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1392 ();
 sky130_fd_sc_hd__nand2_1 _15334_ (.A(net211),
    .B(_04786_),
    .Y(_04810_));
 sky130_fd_sc_hd__o21ai_0 _15335_ (.A1(_04786_),
    .A2(_04808_),
    .B1(_04810_),
    .Y(_00154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1391 ();
 sky130_fd_sc_hd__clkinv_1 _15337_ (.A(_13001_),
    .Y(_04812_));
 sky130_fd_sc_hd__a21o_1 _15338_ (.A1(_12988_),
    .A2(_12993_),
    .B1(_12992_),
    .X(_04813_));
 sky130_fd_sc_hd__a21oi_2 _15339_ (.A1(_12997_),
    .A2(_04813_),
    .B1(_12996_),
    .Y(_04814_));
 sky130_fd_sc_hd__xnor2_2 _15340_ (.A(_04812_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_4 _15341_ (.A(net348),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21ai_4 _15342_ (.A1(\w[62][4] ),
    .A2(net348),
    .B1(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1390 ();
 sky130_fd_sc_hd__nand2_1 _15344_ (.A(net200),
    .B(_04786_),
    .Y(_04819_));
 sky130_fd_sc_hd__o21ai_0 _15345_ (.A1(_04786_),
    .A2(_04817_),
    .B1(_04819_),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_2 _15346_ (.A(_13000_),
    .Y(_04820_));
 sky130_fd_sc_hd__o21ai_2 _15347_ (.A1(_12996_),
    .A2(_04805_),
    .B1(_13001_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21boi_4 _15348_ (.A1(_04820_),
    .A2(_04821_),
    .B1_N(_13005_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand2_1 _15349_ (.A(_04820_),
    .B(_04821_),
    .Y(_04823_));
 sky130_fd_sc_hd__nor2_1 _15350_ (.A(_13005_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__o21ai_4 _15351_ (.A1(_04822_),
    .A2(_04824_),
    .B1(net348),
    .Y(_04825_));
 sky130_fd_sc_hd__o21ai_4 _15352_ (.A1(\w[62][5] ),
    .A2(net348),
    .B1(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1389 ();
 sky130_fd_sc_hd__nand2_1 _15354_ (.A(net189),
    .B(_04786_),
    .Y(_04828_));
 sky130_fd_sc_hd__o21ai_0 _15355_ (.A1(_04786_),
    .A2(_04826_),
    .B1(_04828_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _15356_ (.A(_13009_),
    .Y(_04829_));
 sky130_fd_sc_hd__o21ai_1 _15357_ (.A1(_04812_),
    .A2(_04814_),
    .B1(_04820_),
    .Y(_04830_));
 sky130_fd_sc_hd__a21oi_2 _15358_ (.A1(_13005_),
    .A2(_04830_),
    .B1(_13004_),
    .Y(_04831_));
 sky130_fd_sc_hd__xnor2_1 _15359_ (.A(_04829_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__nand2_2 _15360_ (.A(net348),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__o21ai_4 _15361_ (.A1(\w[62][6] ),
    .A2(net348),
    .B1(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1388 ();
 sky130_fd_sc_hd__nand2_1 _15363_ (.A(net178),
    .B(_04786_),
    .Y(_04836_));
 sky130_fd_sc_hd__o21ai_0 _15364_ (.A1(_04786_),
    .A2(_04834_),
    .B1(_04836_),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_4 _15365_ (.A(_13008_),
    .Y(_04837_));
 sky130_fd_sc_hd__o21ai_2 _15366_ (.A1(_13004_),
    .A2(_04822_),
    .B1(_13009_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21boi_4 _15367_ (.A1(_04837_),
    .A2(_04838_),
    .B1_N(_13013_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand2_1 _15368_ (.A(_04837_),
    .B(_04838_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_1 _15369_ (.A(_13013_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__o21ai_4 _15370_ (.A1(_04839_),
    .A2(_04841_),
    .B1(net348),
    .Y(_04842_));
 sky130_fd_sc_hd__o21ai_4 _15371_ (.A1(\w[62][7] ),
    .A2(net348),
    .B1(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1387 ();
 sky130_fd_sc_hd__nand2_1 _15373_ (.A(net167),
    .B(_04786_),
    .Y(_04845_));
 sky130_fd_sc_hd__o21ai_0 _15374_ (.A1(_04786_),
    .A2(_04843_),
    .B1(_04845_),
    .Y(_00158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1385 ();
 sky130_fd_sc_hd__o21ai_4 _15377_ (.A1(_04829_),
    .A2(_04831_),
    .B1(_04837_),
    .Y(_04848_));
 sky130_fd_sc_hd__a21oi_4 _15378_ (.A1(_13013_),
    .A2(_04848_),
    .B1(_13012_),
    .Y(_04849_));
 sky130_fd_sc_hd__xor2_4 _15379_ (.A(_13017_),
    .B(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__nor2_4 _15380_ (.A(net362),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__a21oi_4 _15381_ (.A1(\w[62][8] ),
    .A2(net361),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1384 ();
 sky130_fd_sc_hd__nand2_1 _15383_ (.A(net156),
    .B(_04786_),
    .Y(_04854_));
 sky130_fd_sc_hd__o21ai_0 _15384_ (.A1(_04786_),
    .A2(_04852_),
    .B1(_04854_),
    .Y(_00159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1383 ();
 sky130_fd_sc_hd__o21ai_2 _15386_ (.A1(_13012_),
    .A2(_04839_),
    .B1(_13017_),
    .Y(_04856_));
 sky130_fd_sc_hd__nand2b_4 _15387_ (.A_N(_13016_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__xnor2_4 _15388_ (.A(_13021_),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__nor2_4 _15389_ (.A(net362),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__a21oi_4 _15390_ (.A1(\w[62][9] ),
    .A2(net362),
    .B1(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1382 ();
 sky130_fd_sc_hd__nand2_1 _15392_ (.A(net145),
    .B(_04786_),
    .Y(_04862_));
 sky130_fd_sc_hd__o21ai_0 _15393_ (.A1(_04786_),
    .A2(_04860_),
    .B1(_04862_),
    .Y(_00160_));
 sky130_fd_sc_hd__clkinv_1 _15394_ (.A(_13020_),
    .Y(_04863_));
 sky130_fd_sc_hd__a211o_4 _15395_ (.A1(_13013_),
    .A2(_04848_),
    .B1(_13016_),
    .C1(_13012_),
    .X(_04864_));
 sky130_fd_sc_hd__o21a_4 _15396_ (.A1(_13017_),
    .A2(_13016_),
    .B1(_13021_),
    .X(_04865_));
 sky130_fd_sc_hd__nand2_2 _15397_ (.A(_04864_),
    .B(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__inv_1 _15398_ (.A(_13025_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21oi_2 _15399_ (.A1(_04863_),
    .A2(_04866_),
    .B1(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__and3_4 _15400_ (.A(_04867_),
    .B(_04863_),
    .C(_04866_),
    .X(_04869_));
 sky130_fd_sc_hd__nor3_4 _15401_ (.A(net363),
    .B(_04868_),
    .C(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__a21oi_4 _15402_ (.A1(\w[62][10] ),
    .A2(net362),
    .B1(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1380 ();
 sky130_fd_sc_hd__nand2_1 _15405_ (.A(net134),
    .B(_04786_),
    .Y(_04874_));
 sky130_fd_sc_hd__o21ai_0 _15406_ (.A1(_04786_),
    .A2(_04871_),
    .B1(_04874_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _15407_ (.A(_13021_),
    .B(_13016_),
    .Y(_04875_));
 sky130_fd_sc_hd__nand2_1 _15408_ (.A(_04863_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21oi_2 _15409_ (.A1(_13025_),
    .A2(_04876_),
    .B1(_13024_),
    .Y(_04877_));
 sky130_fd_sc_hd__o2111ai_2 _15410_ (.A1(_13012_),
    .A2(_04839_),
    .B1(_13017_),
    .C1(_13021_),
    .D1(_13025_),
    .Y(_04878_));
 sky130_fd_sc_hd__a21boi_4 _15411_ (.A1(_04877_),
    .A2(_04878_),
    .B1_N(_13029_),
    .Y(_04879_));
 sky130_fd_sc_hd__nand2_1 _15412_ (.A(_04877_),
    .B(_04878_),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _15413_ (.A(_13029_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__o21ai_2 _15414_ (.A1(_04879_),
    .A2(_04881_),
    .B1(net348),
    .Y(_04882_));
 sky130_fd_sc_hd__o21ai_4 _15415_ (.A1(\w[62][11] ),
    .A2(net348),
    .B1(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1379 ();
 sky130_fd_sc_hd__nand2_1 _15417_ (.A(net123),
    .B(_04786_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21ai_0 _15418_ (.A1(_04786_),
    .A2(_04883_),
    .B1(_04885_),
    .Y(_00131_));
 sky130_fd_sc_hd__a2111oi_4 _15419_ (.A1(_04864_),
    .A2(_04865_),
    .B1(_13020_),
    .C1(_13024_),
    .D1(_13028_),
    .Y(_04886_));
 sky130_fd_sc_hd__or2_4 _15420_ (.A(_13025_),
    .B(_13024_),
    .X(_04887_));
 sky130_fd_sc_hd__a21oi_2 _15421_ (.A1(_13029_),
    .A2(_04887_),
    .B1(_13028_),
    .Y(_04888_));
 sky130_fd_sc_hd__nor2_2 _15422_ (.A(_04886_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__xnor2_1 _15423_ (.A(_13033_),
    .B(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand2_2 _15424_ (.A(net348),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_4 _15425_ (.A1(\w[62][12] ),
    .A2(net348),
    .B1(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1378 ();
 sky130_fd_sc_hd__nand2_1 _15427_ (.A(net111),
    .B(_04786_),
    .Y(_04894_));
 sky130_fd_sc_hd__o21ai_0 _15428_ (.A1(_04786_),
    .A2(_04892_),
    .B1(_04894_),
    .Y(_00132_));
 sky130_fd_sc_hd__or2_4 _15429_ (.A(_13028_),
    .B(_04879_),
    .X(_04895_));
 sky130_fd_sc_hd__a21o_1 _15430_ (.A1(_13033_),
    .A2(_04895_),
    .B1(_13032_),
    .X(_04896_));
 sky130_fd_sc_hd__xnor2_1 _15431_ (.A(_13037_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__nand2_4 _15432_ (.A(net348),
    .B(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__o21ai_4 _15433_ (.A1(\w[62][13] ),
    .A2(net348),
    .B1(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1377 ();
 sky130_fd_sc_hd__nand2_1 _15435_ (.A(net100),
    .B(_04786_),
    .Y(_04901_));
 sky130_fd_sc_hd__o21ai_0 _15436_ (.A1(_04786_),
    .A2(_04899_),
    .B1(_04901_),
    .Y(_00133_));
 sky130_fd_sc_hd__a21o_1 _15437_ (.A1(_13033_),
    .A2(_04889_),
    .B1(_13032_),
    .X(_04902_));
 sky130_fd_sc_hd__a21oi_1 _15438_ (.A1(_13037_),
    .A2(_04902_),
    .B1(_13036_),
    .Y(_04903_));
 sky130_fd_sc_hd__xor2_1 _15439_ (.A(_13041_),
    .B(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__nor2_2 _15440_ (.A(net363),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21oi_4 _15441_ (.A1(\w[62][14] ),
    .A2(net361),
    .B1(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1376 ();
 sky130_fd_sc_hd__nand2_1 _15443_ (.A(net89),
    .B(_04786_),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ai_0 _15444_ (.A1(_04786_),
    .A2(_04906_),
    .B1(_04908_),
    .Y(_00134_));
 sky130_fd_sc_hd__a21o_1 _15445_ (.A1(_13037_),
    .A2(_04896_),
    .B1(_13036_),
    .X(_04909_));
 sky130_fd_sc_hd__a21oi_2 _15446_ (.A1(_13041_),
    .A2(_04909_),
    .B1(_13040_),
    .Y(_04910_));
 sky130_fd_sc_hd__xnor2_4 _15447_ (.A(_13045_),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1375 ();
 sky130_fd_sc_hd__mux2i_4 _15449_ (.A0(\w[62][15] ),
    .A1(_04911_),
    .S(net348),
    .Y(_04913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1374 ();
 sky130_fd_sc_hd__nand2_1 _15451_ (.A(net78),
    .B(_04786_),
    .Y(_04915_));
 sky130_fd_sc_hd__o21ai_0 _15452_ (.A1(_04786_),
    .A2(_04913_),
    .B1(_04915_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand4_1 _15453_ (.A(_13033_),
    .B(_13037_),
    .C(_13041_),
    .D(_13045_),
    .Y(_04916_));
 sky130_fd_sc_hd__a21o_1 _15454_ (.A1(_13037_),
    .A2(_13032_),
    .B1(_13036_),
    .X(_04917_));
 sky130_fd_sc_hd__a21o_1 _15455_ (.A1(_13041_),
    .A2(_04917_),
    .B1(_13040_),
    .X(_04918_));
 sky130_fd_sc_hd__a21oi_2 _15456_ (.A1(_13045_),
    .A2(_04918_),
    .B1(_13044_),
    .Y(_04919_));
 sky130_fd_sc_hd__o31ai_2 _15457_ (.A1(_04886_),
    .A2(_04888_),
    .A3(_04916_),
    .B1(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__xnor2_1 _15458_ (.A(_13049_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_4 _15459_ (.A(net348),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21ai_4 _15460_ (.A1(\w[62][16] ),
    .A2(net348),
    .B1(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1373 ();
 sky130_fd_sc_hd__nand2_1 _15462_ (.A(net67),
    .B(_04786_),
    .Y(_04925_));
 sky130_fd_sc_hd__o21ai_0 _15463_ (.A1(_04786_),
    .A2(_04923_),
    .B1(_04925_),
    .Y(_00136_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1372 ();
 sky130_fd_sc_hd__nor2_1 _15465_ (.A(_13028_),
    .B(_04879_),
    .Y(_04927_));
 sky130_fd_sc_hd__o21ai_0 _15466_ (.A1(_04927_),
    .A2(_04916_),
    .B1(_04919_),
    .Y(_04928_));
 sky130_fd_sc_hd__a21oi_1 _15467_ (.A1(_13049_),
    .A2(_04928_),
    .B1(_13048_),
    .Y(_04929_));
 sky130_fd_sc_hd__xor2_2 _15468_ (.A(_13053_),
    .B(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__nor2_1 _15469_ (.A(net361),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__a21oi_4 _15470_ (.A1(\w[62][17] ),
    .A2(net361),
    .B1(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1371 ();
 sky130_fd_sc_hd__nand2_1 _15472_ (.A(net56),
    .B(_04786_),
    .Y(_04934_));
 sky130_fd_sc_hd__o21ai_0 _15473_ (.A1(_04786_),
    .A2(_04932_),
    .B1(_04934_),
    .Y(_00137_));
 sky130_fd_sc_hd__a21o_1 _15474_ (.A1(_13049_),
    .A2(_04920_),
    .B1(_13048_),
    .X(_04935_));
 sky130_fd_sc_hd__a21oi_1 _15475_ (.A1(_13053_),
    .A2(_04935_),
    .B1(_13052_),
    .Y(_04936_));
 sky130_fd_sc_hd__xor2_1 _15476_ (.A(_13057_),
    .B(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_1 _15477_ (.A(net363),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21oi_4 _15478_ (.A1(\w[62][18] ),
    .A2(net363),
    .B1(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1370 ();
 sky130_fd_sc_hd__nand2_1 _15480_ (.A(net45),
    .B(_04786_),
    .Y(_04941_));
 sky130_fd_sc_hd__o21ai_0 _15481_ (.A1(_04786_),
    .A2(_04939_),
    .B1(_04941_),
    .Y(_00138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1369 ();
 sky130_fd_sc_hd__nand3_1 _15483_ (.A(_13049_),
    .B(_13053_),
    .C(_13057_),
    .Y(_04943_));
 sky130_fd_sc_hd__nor2_2 _15484_ (.A(_04916_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__a21o_1 _15485_ (.A1(_13053_),
    .A2(_13048_),
    .B1(_13052_),
    .X(_04945_));
 sky130_fd_sc_hd__a21o_4 _15486_ (.A1(_13057_),
    .A2(_04945_),
    .B1(_13056_),
    .X(_04946_));
 sky130_fd_sc_hd__or2_4 _15487_ (.A(_04919_),
    .B(_04943_),
    .X(_04947_));
 sky130_fd_sc_hd__nand2b_2 _15488_ (.A_N(_04946_),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__a21oi_2 _15489_ (.A1(_04895_),
    .A2(_04944_),
    .B1(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__xnor2_4 _15490_ (.A(_13061_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__mux2i_4 _15491_ (.A0(\w[62][19] ),
    .A1(_04950_),
    .S(net348),
    .Y(_04951_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1368 ();
 sky130_fd_sc_hd__nand2_1 _15493_ (.A(net34),
    .B(_04786_),
    .Y(_04953_));
 sky130_fd_sc_hd__o21ai_0 _15494_ (.A1(_04786_),
    .A2(_04951_),
    .B1(_04953_),
    .Y(_00139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1367 ();
 sky130_fd_sc_hd__a21oi_1 _15496_ (.A1(_13061_),
    .A2(_04948_),
    .B1(_13060_),
    .Y(_04955_));
 sky130_fd_sc_hd__inv_1 _15497_ (.A(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__a31oi_1 _15498_ (.A1(_13061_),
    .A2(_04889_),
    .A3(_04944_),
    .B1(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__xor2_1 _15499_ (.A(_13065_),
    .B(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__nor2_1 _15500_ (.A(net363),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__a21oi_4 _15501_ (.A1(\w[62][20] ),
    .A2(net363),
    .B1(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1365 ();
 sky130_fd_sc_hd__nand2_1 _15504_ (.A(net23),
    .B(_04786_),
    .Y(_04963_));
 sky130_fd_sc_hd__o21ai_0 _15505_ (.A1(_04786_),
    .A2(_04960_),
    .B1(_04963_),
    .Y(_00141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1364 ();
 sky130_fd_sc_hd__nand4_1 _15507_ (.A(_13049_),
    .B(_13053_),
    .C(_13057_),
    .D(_13028_),
    .Y(_04965_));
 sky130_fd_sc_hd__o21ai_0 _15508_ (.A1(_04916_),
    .A2(_04965_),
    .B1(_04947_),
    .Y(_04966_));
 sky130_fd_sc_hd__a21oi_2 _15509_ (.A1(_04879_),
    .A2(_04944_),
    .B1(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nor3_2 _15510_ (.A(_13060_),
    .B(_13064_),
    .C(_04946_),
    .Y(_04968_));
 sky130_fd_sc_hd__or2_0 _15511_ (.A(_13061_),
    .B(_13060_),
    .X(_04969_));
 sky130_fd_sc_hd__a21oi_2 _15512_ (.A1(_13065_),
    .A2(_04969_),
    .B1(_13064_),
    .Y(_04970_));
 sky130_fd_sc_hd__a21oi_2 _15513_ (.A1(_04967_),
    .A2(_04968_),
    .B1(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__xnor2_2 _15514_ (.A(_13069_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_2 _15515_ (.A(net348),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__o21ai_4 _15516_ (.A1(\w[62][21] ),
    .A2(net348),
    .B1(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1363 ();
 sky130_fd_sc_hd__nand2_1 _15518_ (.A(net12),
    .B(_04786_),
    .Y(_04976_));
 sky130_fd_sc_hd__o21ai_0 _15519_ (.A1(_04786_),
    .A2(_04974_),
    .B1(_04976_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand3_1 _15520_ (.A(_13061_),
    .B(_13065_),
    .C(_04944_),
    .Y(_04977_));
 sky130_fd_sc_hd__nor3_2 _15521_ (.A(_04886_),
    .B(_04888_),
    .C(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__nor2b_2 _15522_ (.A(_04955_),
    .B_N(_13065_),
    .Y(_04979_));
 sky130_fd_sc_hd__o31ai_1 _15523_ (.A1(_13064_),
    .A2(_04978_),
    .A3(_04979_),
    .B1(_13069_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2b_1 _15524_ (.A_N(_13068_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__xnor2_1 _15525_ (.A(_13073_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_4 _15526_ (.A(net363),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__a21oi_4 _15527_ (.A1(\w[62][22] ),
    .A2(net362),
    .B1(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1362 ();
 sky130_fd_sc_hd__nand2_1 _15529_ (.A(net783),
    .B(_04786_),
    .Y(_04986_));
 sky130_fd_sc_hd__o21ai_0 _15530_ (.A1(_04786_),
    .A2(_04984_),
    .B1(_04986_),
    .Y(_00143_));
 sky130_fd_sc_hd__a21o_1 _15531_ (.A1(_13069_),
    .A2(_04971_),
    .B1(_13068_),
    .X(_04987_));
 sky130_fd_sc_hd__a21oi_2 _15532_ (.A1(_13073_),
    .A2(_04987_),
    .B1(_13072_),
    .Y(_04988_));
 sky130_fd_sc_hd__xnor2_2 _15533_ (.A(_13077_),
    .B(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__mux2i_4 _15534_ (.A0(\w[62][23] ),
    .A1(_04989_),
    .S(net348),
    .Y(_04990_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1361 ();
 sky130_fd_sc_hd__nand2_1 _15536_ (.A(net772),
    .B(_04786_),
    .Y(_04992_));
 sky130_fd_sc_hd__o21ai_0 _15537_ (.A1(_04786_),
    .A2(_04990_),
    .B1(_04992_),
    .Y(_00144_));
 sky130_fd_sc_hd__and3_1 _15538_ (.A(_13069_),
    .B(_13073_),
    .C(_13077_),
    .X(_04993_));
 sky130_fd_sc_hd__o31ai_2 _15539_ (.A1(_13064_),
    .A2(_04978_),
    .A3(_04979_),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__and2_4 _15540_ (.A(_13073_),
    .B(_13068_),
    .X(_04995_));
 sky130_fd_sc_hd__o21ai_2 _15541_ (.A1(_13072_),
    .A2(_04995_),
    .B1(_13077_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand3b_1 _15542_ (.A_N(_13076_),
    .B(_04994_),
    .C(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__xnor2_4 _15543_ (.A(_13081_),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__nor2_2 _15544_ (.A(net361),
    .B(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__a21oi_4 _15545_ (.A1(\w[62][24] ),
    .A2(net361),
    .B1(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1360 ();
 sky130_fd_sc_hd__nand2_1 _15547_ (.A(net761),
    .B(_04786_),
    .Y(_05002_));
 sky130_fd_sc_hd__o21ai_0 _15548_ (.A1(_04786_),
    .A2(_05000_),
    .B1(_05002_),
    .Y(_00145_));
 sky130_fd_sc_hd__nand4_1 _15549_ (.A(_13069_),
    .B(_13073_),
    .C(_13077_),
    .D(_13081_),
    .Y(_05003_));
 sky130_fd_sc_hd__a211oi_2 _15550_ (.A1(_04967_),
    .A2(_04968_),
    .B1(_04970_),
    .C1(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__o211a_4 _15551_ (.A1(_13072_),
    .A2(_04995_),
    .B1(_13077_),
    .C1(_13081_),
    .X(_05005_));
 sky130_fd_sc_hd__nor2_4 _15552_ (.A(_05004_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__a21oi_1 _15553_ (.A1(_13081_),
    .A2(_13076_),
    .B1(_13080_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_1 _15554_ (.A(_05006_),
    .B(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__xnor2_2 _15555_ (.A(_13085_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__nand2_1 _15556_ (.A(\w[62][25] ),
    .B(net361),
    .Y(_05010_));
 sky130_fd_sc_hd__o21a_4 _15557_ (.A1(net361),
    .A2(_05009_),
    .B1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1359 ();
 sky130_fd_sc_hd__nand2_1 _15559_ (.A(net750),
    .B(_04786_),
    .Y(_05013_));
 sky130_fd_sc_hd__o21ai_0 _15560_ (.A1(_04786_),
    .A2(_05011_),
    .B1(_05013_),
    .Y(_00146_));
 sky130_fd_sc_hd__nor3_2 _15561_ (.A(_13076_),
    .B(_13080_),
    .C(_13084_),
    .Y(_05014_));
 sky130_fd_sc_hd__or2_0 _15562_ (.A(_13081_),
    .B(_13080_),
    .X(_05015_));
 sky130_fd_sc_hd__a21oi_2 _15563_ (.A1(_13085_),
    .A2(_05015_),
    .B1(_13084_),
    .Y(_05016_));
 sky130_fd_sc_hd__a31oi_4 _15564_ (.A1(_04994_),
    .A2(_04996_),
    .A3(_05014_),
    .B1(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__xnor2_2 _15565_ (.A(_13089_),
    .B(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__nor2_4 _15566_ (.A(net361),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__a21oi_4 _15567_ (.A1(\w[62][26] ),
    .A2(net361),
    .B1(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1358 ();
 sky130_fd_sc_hd__nand2_1 _15569_ (.A(net739),
    .B(_04786_),
    .Y(_05022_));
 sky130_fd_sc_hd__o21ai_0 _15570_ (.A1(_04786_),
    .A2(_05020_),
    .B1(_05022_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand2_1 _15571_ (.A(_13085_),
    .B(_13089_),
    .Y(_05023_));
 sky130_fd_sc_hd__inv_1 _15572_ (.A(_13085_),
    .Y(_05024_));
 sky130_fd_sc_hd__o21bai_1 _15573_ (.A1(_05024_),
    .A2(_05007_),
    .B1_N(_13084_),
    .Y(_05025_));
 sky130_fd_sc_hd__a21oi_2 _15574_ (.A1(_13089_),
    .A2(_05025_),
    .B1(_13088_),
    .Y(_05026_));
 sky130_fd_sc_hd__o21ai_2 _15575_ (.A1(_05006_),
    .A2(_05023_),
    .B1(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__xor2_2 _15576_ (.A(_13093_),
    .B(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__mux2i_4 _15577_ (.A0(\w[62][27] ),
    .A1(_05028_),
    .S(net348),
    .Y(_05029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1357 ();
 sky130_fd_sc_hd__nand2_1 _15579_ (.A(net716),
    .B(_04786_),
    .Y(_05031_));
 sky130_fd_sc_hd__o21ai_0 _15580_ (.A1(_04786_),
    .A2(_05029_),
    .B1(_05031_),
    .Y(_00148_));
 sky130_fd_sc_hd__a21o_1 _15581_ (.A1(_13093_),
    .A2(_13088_),
    .B1(_13092_),
    .X(_05032_));
 sky130_fd_sc_hd__a31oi_1 _15582_ (.A1(_13089_),
    .A2(_13093_),
    .A3(_05017_),
    .B1(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__xnor2_2 _15583_ (.A(_13097_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__mux2i_4 _15584_ (.A0(\w[62][28] ),
    .A1(_05034_),
    .S(net348),
    .Y(_05035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1356 ();
 sky130_fd_sc_hd__nand2_1 _15586_ (.A(net605),
    .B(_04786_),
    .Y(_05037_));
 sky130_fd_sc_hd__o21ai_0 _15587_ (.A1(_04786_),
    .A2(_05035_),
    .B1(_05037_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand4_1 _15588_ (.A(_13085_),
    .B(_13089_),
    .C(_13093_),
    .D(_13097_),
    .Y(_05038_));
 sky130_fd_sc_hd__nor2b_1 _15589_ (.A(_05026_),
    .B_N(_13093_),
    .Y(_05039_));
 sky130_fd_sc_hd__o21a_1 _15590_ (.A1(_13092_),
    .A2(_05039_),
    .B1(_13097_),
    .X(_05040_));
 sky130_fd_sc_hd__nor2_1 _15591_ (.A(_13096_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__o21ai_2 _15592_ (.A1(_05006_),
    .A2(_05038_),
    .B1(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__xor2_4 _15593_ (.A(_13101_),
    .B(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__mux2i_4 _15594_ (.A0(\w[62][29] ),
    .A1(_05043_),
    .S(net348),
    .Y(_05044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1355 ();
 sky130_fd_sc_hd__nand2_1 _15596_ (.A(net223),
    .B(_04786_),
    .Y(_05046_));
 sky130_fd_sc_hd__o21ai_0 _15597_ (.A1(_04786_),
    .A2(_05044_),
    .B1(_05046_),
    .Y(_00150_));
 sky130_fd_sc_hd__a21oi_2 _15598_ (.A1(_13089_),
    .A2(_05017_),
    .B1(_13088_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_1 _15599_ (.A(_13097_),
    .B(_13101_),
    .Y(_05048_));
 sky130_fd_sc_hd__nor3_1 _15600_ (.A(_13105_),
    .B(net363),
    .C(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__nand2_1 _15601_ (.A(_13093_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__nand2b_1 _15602_ (.A_N(_13100_),
    .B(_13105_),
    .Y(_05051_));
 sky130_fd_sc_hd__nor3_1 _15603_ (.A(_13096_),
    .B(net363),
    .C(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__nand3b_1 _15604_ (.A_N(_13092_),
    .B(_05047_),
    .C(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__o21ai_0 _15605_ (.A1(_13093_),
    .A2(_13092_),
    .B1(_13097_),
    .Y(_05054_));
 sky130_fd_sc_hd__a21oi_1 _15606_ (.A1(_13101_),
    .A2(_13096_),
    .B1(_13100_),
    .Y(_05055_));
 sky130_fd_sc_hd__o22a_1 _15607_ (.A1(_13105_),
    .A2(_05055_),
    .B1(_05051_),
    .B2(_13101_),
    .X(_05056_));
 sky130_fd_sc_hd__nand2_2 _15608_ (.A(\w[62][30] ),
    .B(done),
    .Y(_05057_));
 sky130_fd_sc_hd__o21ai_0 _15609_ (.A1(net363),
    .A2(_05056_),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__a221oi_1 _15610_ (.A1(_05052_),
    .A2(_05054_),
    .B1(_05049_),
    .B2(_13092_),
    .C1(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__o211a_4 _15611_ (.A1(_05047_),
    .A2(_05050_),
    .B1(_05053_),
    .C1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1354 ();
 sky130_fd_sc_hd__nand2_1 _15613_ (.A(net112),
    .B(_04786_),
    .Y(_05062_));
 sky130_fd_sc_hd__o21ai_0 _15614_ (.A1(_04786_),
    .A2(_05060_),
    .B1(_05062_),
    .Y(_00152_));
 sky130_fd_sc_hd__xor2_1 _15615_ (.A(_11822_),
    .B(_11825_),
    .X(_05063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1350 ();
 sky130_fd_sc_hd__mux4_2 _15620_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net489),
    .S1(net494),
    .X(_05068_));
 sky130_fd_sc_hd__mux4_2 _15621_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net489),
    .S1(net494),
    .X(_05069_));
 sky130_fd_sc_hd__mux4_2 _15622_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net489),
    .S1(net494),
    .X(_05070_));
 sky130_fd_sc_hd__mux4_2 _15623_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net489),
    .S1(net494),
    .X(_05071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1349 ();
 sky130_fd_sc_hd__mux4_2 _15625_ (.A0(_05068_),
    .A1(_05069_),
    .A2(_05070_),
    .A3(_05071_),
    .S0(net482),
    .S1(net480),
    .X(_05073_));
 sky130_fd_sc_hd__mux4_2 _15626_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net488),
    .S1(net493),
    .X(_05074_));
 sky130_fd_sc_hd__mux4_2 _15627_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net488),
    .S1(net493),
    .X(_05075_));
 sky130_fd_sc_hd__mux4_2 _15628_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net488),
    .S1(net493),
    .X(_05076_));
 sky130_fd_sc_hd__mux4_2 _15629_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net488),
    .S1(net493),
    .X(_05077_));
 sky130_fd_sc_hd__mux4_2 _15630_ (.A0(_05074_),
    .A1(_05075_),
    .A2(_05076_),
    .A3(_05077_),
    .S0(net483),
    .S1(net481),
    .X(_05078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1348 ();
 sky130_fd_sc_hd__mux2i_4 _15632_ (.A0(_05073_),
    .A1(_05078_),
    .S(net479),
    .Y(_05080_));
 sky130_fd_sc_hd__xnor2_1 _15633_ (.A(_05063_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1344 ();
 sky130_fd_sc_hd__mux4_2 _15638_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05086_));
 sky130_fd_sc_hd__mux4_2 _15639_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05087_));
 sky130_fd_sc_hd__mux4_2 _15640_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05088_));
 sky130_fd_sc_hd__mux4_2 _15641_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1343 ();
 sky130_fd_sc_hd__mux4_2 _15643_ (.A0(_05086_),
    .A1(_05087_),
    .A2(_05088_),
    .A3(_05089_),
    .S0(net403),
    .S1(net402),
    .X(_05091_));
 sky130_fd_sc_hd__mux4_2 _15644_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05092_));
 sky130_fd_sc_hd__mux4_2 _15645_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05093_));
 sky130_fd_sc_hd__mux4_2 _15646_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05094_));
 sky130_fd_sc_hd__mux4_2 _15647_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net408),
    .S1(net414),
    .X(_05095_));
 sky130_fd_sc_hd__mux4_2 _15648_ (.A0(_05092_),
    .A1(_05093_),
    .A2(_05094_),
    .A3(_05095_),
    .S0(net403),
    .S1(net402),
    .X(_05096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1342 ();
 sky130_fd_sc_hd__mux2i_4 _15650_ (.A0(_05091_),
    .A1(_05096_),
    .S(net400),
    .Y(_05098_));
 sky130_fd_sc_hd__xnor2_4 _15651_ (.A(_11428_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_1 _15652_ (.A(_05081_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__xor2_1 _15653_ (.A(_11104_),
    .B(_11300_),
    .X(_05101_));
 sky130_fd_sc_hd__xnor2_1 _15654_ (.A(_11006_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__xnor2_2 _15655_ (.A(_05100_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__and2_4 _15656_ (.A(net348),
    .B(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__inv_1 _15657_ (.A(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__or3_4 _15658_ (.A(_13096_),
    .B(_13100_),
    .C(_05040_),
    .X(_05106_));
 sky130_fd_sc_hd__nor3_1 _15659_ (.A(_05004_),
    .B(_05005_),
    .C(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__clkinv_1 _15660_ (.A(_05038_),
    .Y(_05108_));
 sky130_fd_sc_hd__o221ai_2 _15661_ (.A1(_13101_),
    .A2(_13100_),
    .B1(_05108_),
    .B2(_05106_),
    .C1(_13105_),
    .Y(_05109_));
 sky130_fd_sc_hd__nor3_1 _15662_ (.A(_13104_),
    .B(net363),
    .C(_05103_),
    .Y(_05110_));
 sky130_fd_sc_hd__o21ai_0 _15663_ (.A1(_05107_),
    .A2(_05109_),
    .B1(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__o31a_1 _15664_ (.A1(_05105_),
    .A2(_05107_),
    .A3(_05109_),
    .B1(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__a22o_4 _15665_ (.A1(\w[62][31] ),
    .A2(net362),
    .B1(_05104_),
    .B2(_13104_),
    .X(_05113_));
 sky130_fd_sc_hd__mux2i_1 _15666_ (.A0(_05113_),
    .A1(net1),
    .S(_04786_),
    .Y(_05114_));
 sky130_fd_sc_hd__o21ai_0 _15667_ (.A1(_04786_),
    .A2(_05112_),
    .B1(_05114_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2b_4 _15668_ (.A(net1044),
    .B_N(_13536_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand2_8 _15669_ (.A(_09797_),
    .B(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1341 ();
 sky130_fd_sc_hd__mux2i_4 _15671_ (.A0(_13109_),
    .A1(\w[63][0] ),
    .S(net358),
    .Y(_05118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1339 ();
 sky130_fd_sc_hd__nand2_1 _15674_ (.A(net743),
    .B(_05116_),
    .Y(_05121_));
 sky130_fd_sc_hd__o21ai_0 _15675_ (.A1(_05116_),
    .A2(_05118_),
    .B1(_05121_),
    .Y(_00353_));
 sky130_fd_sc_hd__mux2i_4 _15676_ (.A0(_13112_),
    .A1(\w[63][1] ),
    .S(net358),
    .Y(_05122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1338 ();
 sky130_fd_sc_hd__nand2_1 _15678_ (.A(net742),
    .B(_05116_),
    .Y(_05124_));
 sky130_fd_sc_hd__o21ai_0 _15679_ (.A1(_05116_),
    .A2(_05122_),
    .B1(_05124_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand2_1 _15680_ (.A(_11850_),
    .B(_04797_),
    .Y(_05125_));
 sky130_fd_sc_hd__o21ai_4 _15681_ (.A1(\w[63][2] ),
    .A2(_04797_),
    .B1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1337 ();
 sky130_fd_sc_hd__nand2_1 _15683_ (.A(net741),
    .B(_05116_),
    .Y(_05128_));
 sky130_fd_sc_hd__o21ai_0 _15684_ (.A1(_05116_),
    .A2(_05126_),
    .B1(_05128_),
    .Y(_00375_));
 sky130_fd_sc_hd__nor2b_2 _15685_ (.A(_13120_),
    .B_N(_11849_),
    .Y(_05129_));
 sky130_fd_sc_hd__nor2b_4 _15686_ (.A(_11849_),
    .B_N(_13120_),
    .Y(_05130_));
 sky130_fd_sc_hd__o21ai_4 _15687_ (.A1(_05129_),
    .A2(_05130_),
    .B1(_04797_),
    .Y(_05131_));
 sky130_fd_sc_hd__o21ai_4 _15688_ (.A1(\w[63][3] ),
    .A2(_04797_),
    .B1(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1336 ();
 sky130_fd_sc_hd__nand2_1 _15690_ (.A(net740),
    .B(_05116_),
    .Y(_05134_));
 sky130_fd_sc_hd__o21ai_0 _15691_ (.A1(_05116_),
    .A2(_05132_),
    .B1(_05134_),
    .Y(_00378_));
 sky130_fd_sc_hd__clkinv_1 _15692_ (.A(_13124_),
    .Y(_05135_));
 sky130_fd_sc_hd__a21o_1 _15693_ (.A1(_13111_),
    .A2(_13116_),
    .B1(_13115_),
    .X(_05136_));
 sky130_fd_sc_hd__a21oi_2 _15694_ (.A1(_13120_),
    .A2(_05136_),
    .B1(_13119_),
    .Y(_05137_));
 sky130_fd_sc_hd__xnor2_1 _15695_ (.A(_05135_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_2 _15696_ (.A(_04797_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__o21ai_4 _15697_ (.A1(\w[63][4] ),
    .A2(_04797_),
    .B1(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1335 ();
 sky130_fd_sc_hd__nand2_1 _15699_ (.A(net738),
    .B(_05116_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21ai_0 _15700_ (.A1(_05116_),
    .A2(_05140_),
    .B1(_05142_),
    .Y(_00379_));
 sky130_fd_sc_hd__inv_2 _15701_ (.A(_13123_),
    .Y(_05143_));
 sky130_fd_sc_hd__o21ai_2 _15702_ (.A1(_13119_),
    .A2(_05130_),
    .B1(_13124_),
    .Y(_05144_));
 sky130_fd_sc_hd__a21boi_4 _15703_ (.A1(_05143_),
    .A2(_05144_),
    .B1_N(_13128_),
    .Y(_05145_));
 sky130_fd_sc_hd__nand2_1 _15704_ (.A(_05143_),
    .B(_05144_),
    .Y(_05146_));
 sky130_fd_sc_hd__nor2_1 _15705_ (.A(_13128_),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__o21ai_4 _15706_ (.A1(_05145_),
    .A2(_05147_),
    .B1(_04797_),
    .Y(_05148_));
 sky130_fd_sc_hd__o21ai_4 _15707_ (.A1(\w[63][5] ),
    .A2(_04797_),
    .B1(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1334 ();
 sky130_fd_sc_hd__nand2_1 _15709_ (.A(net737),
    .B(_05116_),
    .Y(_05151_));
 sky130_fd_sc_hd__o21ai_0 _15710_ (.A1(_05116_),
    .A2(_05149_),
    .B1(_05151_),
    .Y(_00380_));
 sky130_fd_sc_hd__clkinv_1 _15711_ (.A(_13132_),
    .Y(_05152_));
 sky130_fd_sc_hd__o21ai_2 _15712_ (.A1(_05135_),
    .A2(_05137_),
    .B1(_05143_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21oi_2 _15713_ (.A1(_13128_),
    .A2(_05153_),
    .B1(_13127_),
    .Y(_05154_));
 sky130_fd_sc_hd__xnor2_1 _15714_ (.A(_05152_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_2 _15715_ (.A(_04797_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__o21ai_4 _15716_ (.A1(\w[63][6] ),
    .A2(_04797_),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1333 ();
 sky130_fd_sc_hd__nand2_1 _15718_ (.A(net736),
    .B(_05116_),
    .Y(_05159_));
 sky130_fd_sc_hd__o21ai_0 _15719_ (.A1(_05116_),
    .A2(_05157_),
    .B1(_05159_),
    .Y(_00381_));
 sky130_fd_sc_hd__clkinvlp_2 _15720_ (.A(_13131_),
    .Y(_05160_));
 sky130_fd_sc_hd__o21ai_2 _15721_ (.A1(_13127_),
    .A2(_05145_),
    .B1(_13132_),
    .Y(_05161_));
 sky130_fd_sc_hd__a21boi_4 _15722_ (.A1(_05160_),
    .A2(_05161_),
    .B1_N(_13136_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_1 _15723_ (.A(_05160_),
    .B(_05161_),
    .Y(_05163_));
 sky130_fd_sc_hd__nor2_1 _15724_ (.A(_13136_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__o21ai_2 _15725_ (.A1(_05162_),
    .A2(_05164_),
    .B1(_04797_),
    .Y(_05165_));
 sky130_fd_sc_hd__o21ai_4 _15726_ (.A1(\w[63][7] ),
    .A2(_04797_),
    .B1(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1332 ();
 sky130_fd_sc_hd__nand2_1 _15728_ (.A(net735),
    .B(_05116_),
    .Y(_05168_));
 sky130_fd_sc_hd__o21ai_0 _15729_ (.A1(_05116_),
    .A2(_05166_),
    .B1(_05168_),
    .Y(_00382_));
 sky130_fd_sc_hd__o21ai_2 _15730_ (.A1(_05152_),
    .A2(_05154_),
    .B1(_05160_),
    .Y(_05169_));
 sky130_fd_sc_hd__a21oi_1 _15731_ (.A1(_13136_),
    .A2(_05169_),
    .B1(_13135_),
    .Y(_05170_));
 sky130_fd_sc_hd__xor2_1 _15732_ (.A(_13140_),
    .B(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nor2_1 _15733_ (.A(net359),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__a21oi_4 _15734_ (.A1(\w[63][8] ),
    .A2(net359),
    .B1(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1331 ();
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(net734),
    .B(_05116_),
    .Y(_05175_));
 sky130_fd_sc_hd__o21ai_0 _15737_ (.A1(_05116_),
    .A2(_05173_),
    .B1(_05175_),
    .Y(_00383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1330 ();
 sky130_fd_sc_hd__clkinv_1 _15739_ (.A(_13139_),
    .Y(_05177_));
 sky130_fd_sc_hd__o21ai_2 _15740_ (.A1(_13135_),
    .A2(_05162_),
    .B1(_13140_),
    .Y(_05178_));
 sky130_fd_sc_hd__nand2_1 _15741_ (.A(_05177_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__and2_4 _15742_ (.A(_13144_),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__nor2_1 _15743_ (.A(_13144_),
    .B(_05179_),
    .Y(_05181_));
 sky130_fd_sc_hd__o21ai_2 _15744_ (.A1(_05180_),
    .A2(_05181_),
    .B1(net348),
    .Y(_05182_));
 sky130_fd_sc_hd__o21ai_4 _15745_ (.A1(\w[63][9] ),
    .A2(net348),
    .B1(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1329 ();
 sky130_fd_sc_hd__nand2_1 _15747_ (.A(net733),
    .B(_05116_),
    .Y(_05185_));
 sky130_fd_sc_hd__o21ai_0 _15748_ (.A1(_05116_),
    .A2(_05183_),
    .B1(_05185_),
    .Y(_00384_));
 sky130_fd_sc_hd__a211o_4 _15749_ (.A1(_13136_),
    .A2(_05169_),
    .B1(_13139_),
    .C1(_13135_),
    .X(_05186_));
 sky130_fd_sc_hd__o21ai_0 _15750_ (.A1(_13140_),
    .A2(_13139_),
    .B1(_13144_),
    .Y(_05187_));
 sky130_fd_sc_hd__inv_2 _15751_ (.A(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__a21o_1 _15752_ (.A1(_05186_),
    .A2(_05188_),
    .B1(_13143_),
    .X(_05189_));
 sky130_fd_sc_hd__xnor2_1 _15753_ (.A(_13148_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nor2_2 _15754_ (.A(net364),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__a21oi_4 _15755_ (.A1(\w[63][10] ),
    .A2(net359),
    .B1(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1327 ();
 sky130_fd_sc_hd__nand2_1 _15758_ (.A(net732),
    .B(_05116_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21ai_0 _15759_ (.A1(_05116_),
    .A2(_05192_),
    .B1(_05195_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand3_2 _15760_ (.A(_13144_),
    .B(_13148_),
    .C(_13152_),
    .Y(_05196_));
 sky130_fd_sc_hd__a21oi_4 _15761_ (.A1(_05177_),
    .A2(_05178_),
    .B1(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__a21oi_2 _15762_ (.A1(_13148_),
    .A2(_13143_),
    .B1(_13147_),
    .Y(_05198_));
 sky130_fd_sc_hd__nor2b_4 _15763_ (.A(_05198_),
    .B_N(_13152_),
    .Y(_05199_));
 sky130_fd_sc_hd__nor2_2 _15764_ (.A(_05197_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__o21ai_0 _15765_ (.A1(_13143_),
    .A2(_05180_),
    .B1(_13148_),
    .Y(_05201_));
 sky130_fd_sc_hd__or3b_1 _15766_ (.A(_13152_),
    .B(_13147_),
    .C_N(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__and3_4 _15767_ (.A(net348),
    .B(_05200_),
    .C(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__a21oi_4 _15768_ (.A1(\w[63][11] ),
    .A2(net364),
    .B1(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1326 ();
 sky130_fd_sc_hd__nand2_1 _15770_ (.A(net731),
    .B(_05116_),
    .Y(_05206_));
 sky130_fd_sc_hd__o21ai_0 _15771_ (.A1(_05116_),
    .A2(_05204_),
    .B1(_05206_),
    .Y(_00355_));
 sky130_fd_sc_hd__inv_1 _15772_ (.A(_13156_),
    .Y(_05207_));
 sky130_fd_sc_hd__a2111oi_2 _15773_ (.A1(_05186_),
    .A2(_05188_),
    .B1(_13143_),
    .C1(_13147_),
    .D1(_13151_),
    .Y(_05208_));
 sky130_fd_sc_hd__or2_0 _15774_ (.A(_13148_),
    .B(_13147_),
    .X(_05209_));
 sky130_fd_sc_hd__a21oi_2 _15775_ (.A1(_13152_),
    .A2(_05209_),
    .B1(_13151_),
    .Y(_05210_));
 sky130_fd_sc_hd__or2_4 _15776_ (.A(_05208_),
    .B(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__xnor2_1 _15777_ (.A(_05207_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_1 _15778_ (.A(_04797_),
    .B(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__o21ai_4 _15779_ (.A1(\w[63][12] ),
    .A2(_04797_),
    .B1(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1325 ();
 sky130_fd_sc_hd__nand2_1 _15781_ (.A(net730),
    .B(_05116_),
    .Y(_05216_));
 sky130_fd_sc_hd__o21ai_0 _15782_ (.A1(_05116_),
    .A2(_05214_),
    .B1(_05216_),
    .Y(_00356_));
 sky130_fd_sc_hd__or3_1 _15783_ (.A(_13151_),
    .B(_05197_),
    .C(_05199_),
    .X(_05217_));
 sky130_fd_sc_hd__a21oi_1 _15784_ (.A1(_13156_),
    .A2(_05217_),
    .B1(_13155_),
    .Y(_05218_));
 sky130_fd_sc_hd__xor2_1 _15785_ (.A(_13160_),
    .B(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__nor2_4 _15786_ (.A(net364),
    .B(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__a21oi_4 _15787_ (.A1(\w[63][13] ),
    .A2(net364),
    .B1(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1324 ();
 sky130_fd_sc_hd__nand2_1 _15789_ (.A(net727),
    .B(_05116_),
    .Y(_05223_));
 sky130_fd_sc_hd__o21ai_0 _15790_ (.A1(_05116_),
    .A2(_05221_),
    .B1(_05223_),
    .Y(_00357_));
 sky130_fd_sc_hd__o21bai_1 _15791_ (.A1(_05207_),
    .A2(_05211_),
    .B1_N(_13155_),
    .Y(_05224_));
 sky130_fd_sc_hd__a21oi_1 _15792_ (.A1(_13160_),
    .A2(_05224_),
    .B1(_13159_),
    .Y(_05225_));
 sky130_fd_sc_hd__xor2_2 _15793_ (.A(_13164_),
    .B(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__nor2_2 _15794_ (.A(net358),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__a21oi_4 _15795_ (.A1(\w[63][14] ),
    .A2(net358),
    .B1(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1323 ();
 sky130_fd_sc_hd__nand2_1 _15797_ (.A(net715),
    .B(_05116_),
    .Y(_05230_));
 sky130_fd_sc_hd__o21ai_0 _15798_ (.A1(_05116_),
    .A2(_05228_),
    .B1(_05230_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand3_2 _15799_ (.A(_13156_),
    .B(_13160_),
    .C(_13164_),
    .Y(_05231_));
 sky130_fd_sc_hd__a21o_1 _15800_ (.A1(_13156_),
    .A2(_13151_),
    .B1(_13155_),
    .X(_05232_));
 sky130_fd_sc_hd__a21o_1 _15801_ (.A1(_13160_),
    .A2(_05232_),
    .B1(_13159_),
    .X(_05233_));
 sky130_fd_sc_hd__a21oi_2 _15802_ (.A1(_13164_),
    .A2(_05233_),
    .B1(_13163_),
    .Y(_05234_));
 sky130_fd_sc_hd__o21ai_2 _15803_ (.A1(_05200_),
    .A2(_05231_),
    .B1(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__xnor2_2 _15804_ (.A(_13168_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_2 _15805_ (.A(_04797_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__o21ai_4 _15806_ (.A1(\w[63][15] ),
    .A2(_04797_),
    .B1(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1322 ();
 sky130_fd_sc_hd__nand2_1 _15808_ (.A(net704),
    .B(_05116_),
    .Y(_05240_));
 sky130_fd_sc_hd__o21ai_0 _15809_ (.A1(_05116_),
    .A2(_05238_),
    .B1(_05240_),
    .Y(_00359_));
 sky130_fd_sc_hd__a21o_1 _15810_ (.A1(_13160_),
    .A2(_13155_),
    .B1(_13159_),
    .X(_05241_));
 sky130_fd_sc_hd__a21oi_1 _15811_ (.A1(_13164_),
    .A2(_05241_),
    .B1(_13163_),
    .Y(_05242_));
 sky130_fd_sc_hd__o21ai_0 _15812_ (.A1(_05211_),
    .A2(_05231_),
    .B1(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__a21oi_1 _15813_ (.A1(_13168_),
    .A2(_05243_),
    .B1(_13167_),
    .Y(_05244_));
 sky130_fd_sc_hd__xor2_1 _15814_ (.A(_13172_),
    .B(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__nor2_2 _15815_ (.A(net359),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21oi_4 _15816_ (.A1(\w[63][16] ),
    .A2(net359),
    .B1(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1321 ();
 sky130_fd_sc_hd__nand2_1 _15818_ (.A(net693),
    .B(_05116_),
    .Y(_05249_));
 sky130_fd_sc_hd__o21ai_0 _15819_ (.A1(_05116_),
    .A2(_05247_),
    .B1(_05249_),
    .Y(_00360_));
 sky130_fd_sc_hd__nand2_1 _15820_ (.A(_13168_),
    .B(_13172_),
    .Y(_05250_));
 sky130_fd_sc_hd__or2_4 _15821_ (.A(_05231_),
    .B(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__inv_1 _15822_ (.A(_13168_),
    .Y(_05252_));
 sky130_fd_sc_hd__o21bai_1 _15823_ (.A1(_05252_),
    .A2(_05234_),
    .B1_N(_13167_),
    .Y(_05253_));
 sky130_fd_sc_hd__a21oi_2 _15824_ (.A1(_13172_),
    .A2(_05253_),
    .B1(_13171_),
    .Y(_05254_));
 sky130_fd_sc_hd__o21ai_2 _15825_ (.A1(_05200_),
    .A2(_05251_),
    .B1(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__xnor2_4 _15826_ (.A(_13176_),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_2 _15827_ (.A(_04797_),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__o21ai_4 _15828_ (.A1(\w[63][17] ),
    .A2(_04797_),
    .B1(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1320 ();
 sky130_fd_sc_hd__nand2_1 _15830_ (.A(net682),
    .B(_05116_),
    .Y(_05260_));
 sky130_fd_sc_hd__o21ai_0 _15831_ (.A1(_05116_),
    .A2(_05258_),
    .B1(_05260_),
    .Y(_00361_));
 sky130_fd_sc_hd__o21bai_1 _15832_ (.A1(_05252_),
    .A2(_05242_),
    .B1_N(_13167_),
    .Y(_05261_));
 sky130_fd_sc_hd__a21oi_2 _15833_ (.A1(_13172_),
    .A2(_05261_),
    .B1(_13171_),
    .Y(_05262_));
 sky130_fd_sc_hd__o21ai_0 _15834_ (.A1(_05211_),
    .A2(_05251_),
    .B1(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__a21oi_1 _15835_ (.A1(_13176_),
    .A2(_05263_),
    .B1(_13175_),
    .Y(_05264_));
 sky130_fd_sc_hd__xor2_2 _15836_ (.A(_13180_),
    .B(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__nor2_1 _15837_ (.A(net358),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__a21oi_4 _15838_ (.A1(\w[63][18] ),
    .A2(net358),
    .B1(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1319 ();
 sky130_fd_sc_hd__nand2_1 _15840_ (.A(net671),
    .B(_05116_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_0 _15841_ (.A1(_05116_),
    .A2(_05267_),
    .B1(_05269_),
    .Y(_00362_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1318 ();
 sky130_fd_sc_hd__nand2_1 _15843_ (.A(_13176_),
    .B(_13180_),
    .Y(_05271_));
 sky130_fd_sc_hd__nor2_1 _15844_ (.A(_05251_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__o21ai_4 _15845_ (.A1(_05197_),
    .A2(_05199_),
    .B1(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__nor2_2 _15846_ (.A(_05254_),
    .B(_05271_),
    .Y(_05274_));
 sky130_fd_sc_hd__a21oi_4 _15847_ (.A1(_13180_),
    .A2(_13175_),
    .B1(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_1 _15848_ (.A(_05273_),
    .B(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__nor2_1 _15849_ (.A(_13179_),
    .B(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__xor2_1 _15850_ (.A(_13184_),
    .B(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__nor2_1 _15851_ (.A(net359),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__a21oi_4 _15852_ (.A1(\w[63][19] ),
    .A2(net359),
    .B1(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1317 ();
 sky130_fd_sc_hd__nand2_1 _15854_ (.A(net660),
    .B(_05116_),
    .Y(_05282_));
 sky130_fd_sc_hd__o21ai_0 _15855_ (.A1(_05116_),
    .A2(_05280_),
    .B1(_05282_),
    .Y(_00363_));
 sky130_fd_sc_hd__o21a_1 _15856_ (.A1(_13176_),
    .A2(_13175_),
    .B1(_13180_),
    .X(_05283_));
 sky130_fd_sc_hd__o21ai_2 _15857_ (.A1(_13179_),
    .A2(_05283_),
    .B1(_13184_),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2b_4 _15858_ (.A_N(_13183_),
    .B(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__nor3_2 _15859_ (.A(_13175_),
    .B(_13179_),
    .C(_13183_),
    .Y(_05286_));
 sky130_fd_sc_hd__o311ai_4 _15860_ (.A1(_05208_),
    .A2(_05210_),
    .A3(_05251_),
    .B1(_05262_),
    .C1(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__and3_4 _15861_ (.A(_13188_),
    .B(_05285_),
    .C(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__a21oi_2 _15862_ (.A1(_05285_),
    .A2(_05287_),
    .B1(_13188_),
    .Y(_05289_));
 sky130_fd_sc_hd__o21ai_4 _15863_ (.A1(_05288_),
    .A2(_05289_),
    .B1(net348),
    .Y(_05290_));
 sky130_fd_sc_hd__o21ai_4 _15864_ (.A1(\w[63][20] ),
    .A2(net348),
    .B1(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1315 ();
 sky130_fd_sc_hd__nand2_1 _15867_ (.A(net649),
    .B(_05116_),
    .Y(_05294_));
 sky130_fd_sc_hd__o21ai_0 _15868_ (.A1(_05116_),
    .A2(_05291_),
    .B1(_05294_),
    .Y(_00365_));
 sky130_fd_sc_hd__nor2_1 _15869_ (.A(_13179_),
    .B(_13183_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_0 _15870_ (.A1(_13184_),
    .A2(_13183_),
    .B1(_13188_),
    .Y(_05296_));
 sky130_fd_sc_hd__a31oi_1 _15871_ (.A1(_05273_),
    .A2(_05275_),
    .A3(_05295_),
    .B1(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__nor2_1 _15872_ (.A(_13187_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__xor2_1 _15873_ (.A(_13192_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__nor2_1 _15874_ (.A(net359),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__a21oi_4 _15875_ (.A1(\w[63][21] ),
    .A2(net359),
    .B1(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1314 ();
 sky130_fd_sc_hd__nand2_1 _15877_ (.A(net638),
    .B(_05116_),
    .Y(_05303_));
 sky130_fd_sc_hd__o21ai_0 _15878_ (.A1(_05116_),
    .A2(_05301_),
    .B1(_05303_),
    .Y(_00366_));
 sky130_fd_sc_hd__inv_2 _15879_ (.A(_13196_),
    .Y(_05304_));
 sky130_fd_sc_hd__a21o_4 _15880_ (.A1(_13192_),
    .A2(_13187_),
    .B1(_13191_),
    .X(_05305_));
 sky130_fd_sc_hd__a41oi_4 _15881_ (.A1(_13188_),
    .A2(_13192_),
    .A3(_05285_),
    .A4(_05287_),
    .B1(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__xnor2_2 _15882_ (.A(_05304_),
    .B(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__nand2_1 _15883_ (.A(_04797_),
    .B(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__o21ai_4 _15884_ (.A1(\w[63][22] ),
    .A2(_04797_),
    .B1(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1313 ();
 sky130_fd_sc_hd__nand2_1 _15886_ (.A(net627),
    .B(_05116_),
    .Y(_05311_));
 sky130_fd_sc_hd__o21ai_0 _15887_ (.A1(_05116_),
    .A2(_05309_),
    .B1(_05311_),
    .Y(_00367_));
 sky130_fd_sc_hd__nor3_2 _15888_ (.A(_13179_),
    .B(_13183_),
    .C(_05305_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2b_1 _15889_ (.A_N(_13187_),
    .B(_05296_),
    .Y(_05313_));
 sky130_fd_sc_hd__a21o_4 _15890_ (.A1(_13192_),
    .A2(_05313_),
    .B1(_13191_),
    .X(_05314_));
 sky130_fd_sc_hd__nand2_1 _15891_ (.A(_13196_),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__a31oi_2 _15892_ (.A1(_05273_),
    .A2(_05275_),
    .A3(_05312_),
    .B1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__o21a_4 _15893_ (.A1(_13195_),
    .A2(_05316_),
    .B1(_13200_),
    .X(_05317_));
 sky130_fd_sc_hd__nor3_1 _15894_ (.A(_13200_),
    .B(_13195_),
    .C(_05316_),
    .Y(_05318_));
 sky130_fd_sc_hd__o21ai_4 _15895_ (.A1(_05317_),
    .A2(_05318_),
    .B1(_04797_),
    .Y(_05319_));
 sky130_fd_sc_hd__o21ai_4 _15896_ (.A1(\w[63][23] ),
    .A2(_04797_),
    .B1(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1312 ();
 sky130_fd_sc_hd__nand2_1 _15898_ (.A(net616),
    .B(_05116_),
    .Y(_05322_));
 sky130_fd_sc_hd__o21ai_0 _15899_ (.A1(_05116_),
    .A2(_05320_),
    .B1(_05322_),
    .Y(_00368_));
 sky130_fd_sc_hd__o21bai_1 _15900_ (.A1(_05304_),
    .A2(_05306_),
    .B1_N(_13195_),
    .Y(_05323_));
 sky130_fd_sc_hd__a21oi_2 _15901_ (.A1(_13200_),
    .A2(_05323_),
    .B1(_13199_),
    .Y(_05324_));
 sky130_fd_sc_hd__xnor2_4 _15902_ (.A(_13204_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__mux2i_4 _15903_ (.A0(\w[63][24] ),
    .A1(_05325_),
    .S(_04797_),
    .Y(_05326_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1311 ();
 sky130_fd_sc_hd__nand2_1 _15905_ (.A(net604),
    .B(_05116_),
    .Y(_05328_));
 sky130_fd_sc_hd__o21ai_0 _15906_ (.A1(_05116_),
    .A2(_05326_),
    .B1(_05328_),
    .Y(_00369_));
 sky130_fd_sc_hd__o21ai_2 _15907_ (.A1(_13199_),
    .A2(_05317_),
    .B1(_13204_),
    .Y(_05329_));
 sky130_fd_sc_hd__nor2_2 _15908_ (.A(_13208_),
    .B(_13203_),
    .Y(_05330_));
 sky130_fd_sc_hd__a21o_1 _15909_ (.A1(_13200_),
    .A2(_13195_),
    .B1(_13199_),
    .X(_05331_));
 sky130_fd_sc_hd__a21o_4 _15910_ (.A1(_13204_),
    .A2(_05331_),
    .B1(_13203_),
    .X(_05332_));
 sky130_fd_sc_hd__and3_4 _15911_ (.A(_13196_),
    .B(_13200_),
    .C(_13204_),
    .X(_05333_));
 sky130_fd_sc_hd__nand2_1 _15912_ (.A(_05314_),
    .B(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__a31oi_1 _15913_ (.A1(_05273_),
    .A2(_05275_),
    .A3(_05312_),
    .B1(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__o21ai_0 _15914_ (.A1(_05332_),
    .A2(_05335_),
    .B1(_13208_),
    .Y(_05336_));
 sky130_fd_sc_hd__nand2_1 _15915_ (.A(_04797_),
    .B(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__a21oi_4 _15916_ (.A1(_05329_),
    .A2(_05330_),
    .B1(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__a21oi_4 _15917_ (.A1(\w[63][25] ),
    .A2(net358),
    .B1(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1310 ();
 sky130_fd_sc_hd__nand2_1 _15919_ (.A(net593),
    .B(_05116_),
    .Y(_05341_));
 sky130_fd_sc_hd__o21ai_0 _15920_ (.A1(_05116_),
    .A2(_05339_),
    .B1(_05341_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand2_2 _15921_ (.A(_13208_),
    .B(_05333_),
    .Y(_05342_));
 sky130_fd_sc_hd__a21oi_1 _15922_ (.A1(_13208_),
    .A2(_05332_),
    .B1(_13207_),
    .Y(_05343_));
 sky130_fd_sc_hd__o21ai_2 _15923_ (.A1(_05306_),
    .A2(_05342_),
    .B1(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__xnor2_1 _15924_ (.A(_13212_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_2 _15925_ (.A(_04797_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__o21ai_4 _15926_ (.A1(\w[63][26] ),
    .A2(_04797_),
    .B1(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1309 ();
 sky130_fd_sc_hd__nand2_1 _15928_ (.A(net582),
    .B(_05116_),
    .Y(_05349_));
 sky130_fd_sc_hd__o21ai_0 _15929_ (.A1(_05116_),
    .A2(_05347_),
    .B1(_05349_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_1 _15930_ (.A(_13212_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand3_1 _15931_ (.A(_05273_),
    .B(_05275_),
    .C(_05312_),
    .Y(_05351_));
 sky130_fd_sc_hd__nor2b_2 _15932_ (.A(_05342_),
    .B_N(_05314_),
    .Y(_05352_));
 sky130_fd_sc_hd__a21boi_4 _15933_ (.A1(_05351_),
    .A2(_05352_),
    .B1_N(_05343_),
    .Y(_05353_));
 sky130_fd_sc_hd__o21bai_2 _15934_ (.A1(_05350_),
    .A2(_05353_),
    .B1_N(_13211_),
    .Y(_05354_));
 sky130_fd_sc_hd__nor2_1 _15935_ (.A(_13216_),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__and2_0 _15936_ (.A(_13216_),
    .B(_05354_),
    .X(_05356_));
 sky130_fd_sc_hd__nand2_1 _15937_ (.A(\w[63][27] ),
    .B(net360),
    .Y(_05357_));
 sky130_fd_sc_hd__o31a_1 _15938_ (.A1(net360),
    .A2(_05355_),
    .A3(_05356_),
    .B1(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1308 ();
 sky130_fd_sc_hd__nand2_1 _15940_ (.A(net571),
    .B(_05116_),
    .Y(_05360_));
 sky130_fd_sc_hd__o21ai_0 _15941_ (.A1(_05116_),
    .A2(net538),
    .B1(_05360_),
    .Y(_00372_));
 sky130_fd_sc_hd__and4_4 _15942_ (.A(_13188_),
    .B(_13192_),
    .C(_13208_),
    .D(_05333_),
    .X(_05361_));
 sky130_fd_sc_hd__nand2_1 _15943_ (.A(_13208_),
    .B(_05332_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand3_1 _15944_ (.A(_13208_),
    .B(_05305_),
    .C(_05333_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_2 _15945_ (.A(_05362_),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__or3_4 _15946_ (.A(_13207_),
    .B(_13211_),
    .C(_13215_),
    .X(_05365_));
 sky130_fd_sc_hd__a311oi_4 _15947_ (.A1(_05285_),
    .A2(_05287_),
    .A3(_05361_),
    .B1(_05364_),
    .C1(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__or2_0 _15948_ (.A(_13212_),
    .B(_13211_),
    .X(_05367_));
 sky130_fd_sc_hd__a21oi_2 _15949_ (.A1(_13216_),
    .A2(_05367_),
    .B1(_13215_),
    .Y(_05368_));
 sky130_fd_sc_hd__nor2_1 _15950_ (.A(_05366_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__xnor2_1 _15951_ (.A(_13220_),
    .B(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__nor2_2 _15952_ (.A(net360),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__a21oi_4 _15953_ (.A1(\w[63][28] ),
    .A2(net360),
    .B1(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1307 ();
 sky130_fd_sc_hd__nand2_1 _15955_ (.A(net289),
    .B(_05116_),
    .Y(_05374_));
 sky130_fd_sc_hd__o21ai_0 _15956_ (.A1(_05116_),
    .A2(_05372_),
    .B1(_05374_),
    .Y(_00373_));
 sky130_fd_sc_hd__nand3_1 _15957_ (.A(_13212_),
    .B(_13216_),
    .C(_13220_),
    .Y(_05375_));
 sky130_fd_sc_hd__a21o_1 _15958_ (.A1(_13216_),
    .A2(_13211_),
    .B1(_13215_),
    .X(_05376_));
 sky130_fd_sc_hd__a21oi_1 _15959_ (.A1(_13220_),
    .A2(_05376_),
    .B1(_13219_),
    .Y(_05377_));
 sky130_fd_sc_hd__o21ai_2 _15960_ (.A1(_05353_),
    .A2(_05375_),
    .B1(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__xor2_2 _15961_ (.A(_13224_),
    .B(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2i_4 _15962_ (.A0(\w[63][29] ),
    .A1(_05379_),
    .S(_04797_),
    .Y(_05380_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1306 ();
 sky130_fd_sc_hd__nand2_1 _15964_ (.A(net278),
    .B(_05116_),
    .Y(_05382_));
 sky130_fd_sc_hd__o21ai_0 _15965_ (.A1(_05116_),
    .A2(_05380_),
    .B1(_05382_),
    .Y(_00374_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1305 ();
 sky130_fd_sc_hd__nand2_1 _15967_ (.A(_13220_),
    .B(_13224_),
    .Y(_05384_));
 sky130_fd_sc_hd__a21oi_1 _15968_ (.A1(_13224_),
    .A2(_13219_),
    .B1(_13223_),
    .Y(_05385_));
 sky130_fd_sc_hd__o31ai_1 _15969_ (.A1(_05366_),
    .A2(_05368_),
    .A3(_05384_),
    .B1(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__xnor2_1 _15970_ (.A(_13228_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__nor2_1 _15971_ (.A(net360),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__a21oi_4 _15972_ (.A1(\w[63][30] ),
    .A2(net360),
    .B1(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__a21oi_1 _15973_ (.A1(_09797_),
    .A2(_05115_),
    .B1(net267),
    .Y(_05390_));
 sky130_fd_sc_hd__a31oi_1 _15974_ (.A1(_09797_),
    .A2(_05115_),
    .A3(net1134),
    .B1(_05390_),
    .Y(_00376_));
 sky130_fd_sc_hd__nand2_1 _15975_ (.A(_13220_),
    .B(_05376_),
    .Y(_05391_));
 sky130_fd_sc_hd__nor3_1 _15976_ (.A(_13219_),
    .B(_13223_),
    .C(_13227_),
    .Y(_05392_));
 sky130_fd_sc_hd__o211ai_1 _15977_ (.A1(_05353_),
    .A2(_05375_),
    .B1(_05391_),
    .C1(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hd__nor3_1 _15978_ (.A(_13224_),
    .B(_13223_),
    .C(_13227_),
    .Y(_05394_));
 sky130_fd_sc_hd__nor2_1 _15979_ (.A(_13228_),
    .B(_13227_),
    .Y(_05395_));
 sky130_fd_sc_hd__nor2_1 _15980_ (.A(_05394_),
    .B(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__xor2_1 _15981_ (.A(_12070_),
    .B(_12073_),
    .X(_05397_));
 sky130_fd_sc_hd__mux4_2 _15982_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05398_));
 sky130_fd_sc_hd__mux4_2 _15983_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05399_));
 sky130_fd_sc_hd__mux4_2 _15984_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05400_));
 sky130_fd_sc_hd__mux4_2 _15985_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05401_));
 sky130_fd_sc_hd__mux4_2 _15986_ (.A0(_05398_),
    .A1(_05399_),
    .A2(_05400_),
    .A3(_05401_),
    .S0(net462),
    .S1(net460),
    .X(_05402_));
 sky130_fd_sc_hd__mux4_2 _15987_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05403_));
 sky130_fd_sc_hd__mux4_2 _15988_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05404_));
 sky130_fd_sc_hd__mux4_2 _15989_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05405_));
 sky130_fd_sc_hd__mux4_2 _15990_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net467),
    .S1(net475),
    .X(_05406_));
 sky130_fd_sc_hd__mux4_2 _15991_ (.A0(_05403_),
    .A1(_05404_),
    .A2(_05405_),
    .A3(_05406_),
    .S0(net462),
    .S1(net460),
    .X(_05407_));
 sky130_fd_sc_hd__mux2i_4 _15992_ (.A0(_05402_),
    .A1(_05407_),
    .S(\count16_2[5] ),
    .Y(_05408_));
 sky130_fd_sc_hd__xnor2_1 _15993_ (.A(_05397_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__mux4_2 _15994_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net387),
    .S1(net544),
    .X(_05410_));
 sky130_fd_sc_hd__mux4_2 _15995_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net387),
    .S1(net544),
    .X(_05411_));
 sky130_fd_sc_hd__mux4_2 _15996_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net387),
    .S1(net544),
    .X(_05412_));
 sky130_fd_sc_hd__mux4_2 _15997_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net387),
    .S1(net544),
    .X(_05413_));
 sky130_fd_sc_hd__mux4_2 _15998_ (.A0(_05410_),
    .A1(_05411_),
    .A2(_05412_),
    .A3(_05413_),
    .S0(net385),
    .S1(net382),
    .X(_05414_));
 sky130_fd_sc_hd__mux4_2 _15999_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net391),
    .S1(net397),
    .X(_05415_));
 sky130_fd_sc_hd__mux4_2 _16000_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net391),
    .S1(net397),
    .X(_05416_));
 sky130_fd_sc_hd__mux4_2 _16001_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net391),
    .S1(net397),
    .X(_05417_));
 sky130_fd_sc_hd__mux4_2 _16002_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net391),
    .S1(net397),
    .X(_05418_));
 sky130_fd_sc_hd__mux4_2 _16003_ (.A0(_05415_),
    .A1(_05416_),
    .A2(_05417_),
    .A3(_05418_),
    .S0(net384),
    .S1(net542),
    .X(_05419_));
 sky130_fd_sc_hd__mux2i_4 _16004_ (.A0(_05414_),
    .A1(_05419_),
    .S(net380),
    .Y(_05420_));
 sky130_fd_sc_hd__xnor2_4 _16005_ (.A(_03656_),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__xnor2_1 _16006_ (.A(_05409_),
    .B(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__xor2_1 _16007_ (.A(_03194_),
    .B(_03378_),
    .X(_05423_));
 sky130_fd_sc_hd__xnor2_1 _16008_ (.A(_02964_),
    .B(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__xnor2_1 _16009_ (.A(_05422_),
    .B(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__nor2_1 _16010_ (.A(net360),
    .B(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_1 _16011_ (.A(_04797_),
    .B(_05425_),
    .Y(_05427_));
 sky130_fd_sc_hd__a21oi_1 _16012_ (.A1(_05393_),
    .A2(_05396_),
    .B1(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__nor2_4 _16013_ (.A(\w[63][31] ),
    .B(_04797_),
    .Y(_05429_));
 sky130_fd_sc_hd__a311o_1 _16014_ (.A1(_05393_),
    .A2(_05396_),
    .A3(_05426_),
    .B1(_05428_),
    .C1(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1304 ();
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(net256),
    .B(_05116_),
    .Y(_05432_));
 sky130_fd_sc_hd__o21ai_0 _16017_ (.A1(_05116_),
    .A2(net1042),
    .B1(_05432_),
    .Y(_00377_));
 sky130_fd_sc_hd__nor2b_4 _16018_ (.A(net1044),
    .B_N(_13531_),
    .Y(_05433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1303 ();
 sky130_fd_sc_hd__nand2_8 _16020_ (.A(_09735_),
    .B(_05433_),
    .Y(_05435_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1301 ();
 sky130_fd_sc_hd__nand2_1 _16023_ (.A(net778),
    .B(_05435_),
    .Y(_05438_));
 sky130_fd_sc_hd__o21ai_0 _16024_ (.A1(_04790_),
    .A2(_05435_),
    .B1(_05438_),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _16025_ (.A(net777),
    .B(_05435_),
    .Y(_05439_));
 sky130_fd_sc_hd__o21ai_0 _16026_ (.A1(_04794_),
    .A2(_05435_),
    .B1(_05439_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _16027_ (.A(net776),
    .B(_05435_),
    .Y(_05440_));
 sky130_fd_sc_hd__o21ai_0 _16028_ (.A1(_04801_),
    .A2(_05435_),
    .B1(_05440_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand2_1 _16029_ (.A(net775),
    .B(_05435_),
    .Y(_05441_));
 sky130_fd_sc_hd__o21ai_0 _16030_ (.A1(_04808_),
    .A2(_05435_),
    .B1(_05441_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _16031_ (.A(net774),
    .B(_05435_),
    .Y(_05442_));
 sky130_fd_sc_hd__o21ai_0 _16032_ (.A1(_04817_),
    .A2(_05435_),
    .B1(_05442_),
    .Y(_00411_));
 sky130_fd_sc_hd__nand2_1 _16033_ (.A(net773),
    .B(_05435_),
    .Y(_05443_));
 sky130_fd_sc_hd__o21ai_0 _16034_ (.A1(_04826_),
    .A2(_05435_),
    .B1(_05443_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _16035_ (.A(net771),
    .B(_05435_),
    .Y(_05444_));
 sky130_fd_sc_hd__o21ai_0 _16036_ (.A1(_04834_),
    .A2(_05435_),
    .B1(_05444_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _16037_ (.A(net770),
    .B(_05435_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21ai_0 _16038_ (.A1(_04843_),
    .A2(_05435_),
    .B1(_05445_),
    .Y(_00414_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1300 ();
 sky130_fd_sc_hd__nand2_1 _16040_ (.A(net769),
    .B(_05435_),
    .Y(_05447_));
 sky130_fd_sc_hd__o21ai_0 _16041_ (.A1(_04852_),
    .A2(_05435_),
    .B1(_05447_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _16042_ (.A(net768),
    .B(_05435_),
    .Y(_05448_));
 sky130_fd_sc_hd__o21ai_0 _16043_ (.A1(_04860_),
    .A2(_05435_),
    .B1(_05448_),
    .Y(_00416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1299 ();
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(net767),
    .B(_05435_),
    .Y(_05450_));
 sky130_fd_sc_hd__o21ai_0 _16046_ (.A1(_04871_),
    .A2(_05435_),
    .B1(_05450_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _16047_ (.A(net766),
    .B(_05435_),
    .Y(_05451_));
 sky130_fd_sc_hd__o21ai_0 _16048_ (.A1(_04883_),
    .A2(_05435_),
    .B1(_05451_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _16049_ (.A(net765),
    .B(_05435_),
    .Y(_05452_));
 sky130_fd_sc_hd__o21ai_0 _16050_ (.A1(_04892_),
    .A2(_05435_),
    .B1(_05452_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _16051_ (.A(net764),
    .B(_05435_),
    .Y(_05453_));
 sky130_fd_sc_hd__o21ai_0 _16052_ (.A1(_04899_),
    .A2(_05435_),
    .B1(_05453_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _16053_ (.A(net763),
    .B(_05435_),
    .Y(_05454_));
 sky130_fd_sc_hd__o21ai_0 _16054_ (.A1(_04906_),
    .A2(_05435_),
    .B1(_05454_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _16055_ (.A(net762),
    .B(_05435_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21ai_0 _16056_ (.A1(_04913_),
    .A2(_05435_),
    .B1(_05455_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_1 _16057_ (.A(net760),
    .B(_05435_),
    .Y(_05456_));
 sky130_fd_sc_hd__o21ai_0 _16058_ (.A1(_04923_),
    .A2(_05435_),
    .B1(_05456_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand2_1 _16059_ (.A(net759),
    .B(_05435_),
    .Y(_05457_));
 sky130_fd_sc_hd__o21ai_0 _16060_ (.A1(_04932_),
    .A2(_05435_),
    .B1(_05457_),
    .Y(_00393_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1298 ();
 sky130_fd_sc_hd__nand2_1 _16062_ (.A(net758),
    .B(_05435_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21ai_0 _16063_ (.A1(_04939_),
    .A2(_05435_),
    .B1(_05459_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _16064_ (.A(net757),
    .B(_05435_),
    .Y(_05460_));
 sky130_fd_sc_hd__o21ai_0 _16065_ (.A1(_04951_),
    .A2(_05435_),
    .B1(_05460_),
    .Y(_00395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1297 ();
 sky130_fd_sc_hd__nand2_1 _16067_ (.A(net756),
    .B(_05435_),
    .Y(_05462_));
 sky130_fd_sc_hd__o21ai_0 _16068_ (.A1(_04960_),
    .A2(_05435_),
    .B1(_05462_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _16069_ (.A(net755),
    .B(_05435_),
    .Y(_05463_));
 sky130_fd_sc_hd__o21ai_0 _16070_ (.A1(_04974_),
    .A2(_05435_),
    .B1(_05463_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(net754),
    .B(_05435_),
    .Y(_05464_));
 sky130_fd_sc_hd__o21ai_0 _16072_ (.A1(_04984_),
    .A2(_05435_),
    .B1(_05464_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _16073_ (.A(net753),
    .B(_05435_),
    .Y(_05465_));
 sky130_fd_sc_hd__o21ai_0 _16074_ (.A1(_04990_),
    .A2(_05435_),
    .B1(_05465_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _16075_ (.A(net752),
    .B(_05435_),
    .Y(_05466_));
 sky130_fd_sc_hd__o21ai_0 _16076_ (.A1(_05000_),
    .A2(_05435_),
    .B1(_05466_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _16077_ (.A(net751),
    .B(_05435_),
    .Y(_05467_));
 sky130_fd_sc_hd__o21ai_0 _16078_ (.A1(_05011_),
    .A2(_05435_),
    .B1(_05467_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _16079_ (.A(net749),
    .B(_05435_),
    .Y(_05468_));
 sky130_fd_sc_hd__o21ai_0 _16080_ (.A1(_05020_),
    .A2(_05435_),
    .B1(_05468_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(net748),
    .B(_05435_),
    .Y(_05469_));
 sky130_fd_sc_hd__o21ai_0 _16082_ (.A1(_05029_),
    .A2(_05435_),
    .B1(_05469_),
    .Y(_00404_));
 sky130_fd_sc_hd__nand2_1 _16083_ (.A(net747),
    .B(_05435_),
    .Y(_05470_));
 sky130_fd_sc_hd__o21ai_0 _16084_ (.A1(_05035_),
    .A2(_05435_),
    .B1(_05470_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _16085_ (.A(net746),
    .B(_05435_),
    .Y(_05471_));
 sky130_fd_sc_hd__o21ai_0 _16086_ (.A1(_05044_),
    .A2(_05435_),
    .B1(_05471_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _16087_ (.A(net745),
    .B(_05435_),
    .Y(_05472_));
 sky130_fd_sc_hd__o21ai_0 _16088_ (.A1(_05060_),
    .A2(_05435_),
    .B1(_05472_),
    .Y(_00408_));
 sky130_fd_sc_hd__mux2i_1 _16089_ (.A0(_05113_),
    .A1(net744),
    .S(_05435_),
    .Y(_05473_));
 sky130_fd_sc_hd__o21ai_0 _16090_ (.A1(_05112_),
    .A2(_05435_),
    .B1(_05473_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2b_4 _16091_ (.A(net1044),
    .B_N(_13539_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand2_8 _16092_ (.A(_09797_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1295 ();
 sky130_fd_sc_hd__nand2_1 _16095_ (.A(net31),
    .B(_05475_),
    .Y(_05478_));
 sky130_fd_sc_hd__o21ai_0 _16096_ (.A1(_05118_),
    .A2(_05475_),
    .B1(_05478_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(net30),
    .B(_05475_),
    .Y(_05479_));
 sky130_fd_sc_hd__o21ai_0 _16098_ (.A1(_05122_),
    .A2(_05475_),
    .B1(_05479_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _16099_ (.A(net29),
    .B(_05475_),
    .Y(_05480_));
 sky130_fd_sc_hd__o21ai_0 _16100_ (.A1(_05126_),
    .A2(_05475_),
    .B1(_05480_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(net28),
    .B(_05475_),
    .Y(_05481_));
 sky130_fd_sc_hd__o21ai_0 _16102_ (.A1(_05132_),
    .A2(_05475_),
    .B1(_05481_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _16103_ (.A(net27),
    .B(_05475_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21ai_0 _16104_ (.A1(_05140_),
    .A2(_05475_),
    .B1(_05482_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _16105_ (.A(net26),
    .B(_05475_),
    .Y(_05483_));
 sky130_fd_sc_hd__o21ai_0 _16106_ (.A1(_05149_),
    .A2(_05475_),
    .B1(_05483_),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _16107_ (.A(net25),
    .B(_05475_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21ai_0 _16108_ (.A1(_05157_),
    .A2(_05475_),
    .B1(_05484_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(net24),
    .B(_05475_),
    .Y(_05485_));
 sky130_fd_sc_hd__o21ai_0 _16110_ (.A1(_05166_),
    .A2(_05475_),
    .B1(_05485_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _16111_ (.A(net22),
    .B(_05475_),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_0 _16112_ (.A1(_05173_),
    .A2(_05475_),
    .B1(_05486_),
    .Y(_00447_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1294 ();
 sky130_fd_sc_hd__nand2_1 _16114_ (.A(net21),
    .B(_05475_),
    .Y(_05488_));
 sky130_fd_sc_hd__o21ai_0 _16115_ (.A1(_05183_),
    .A2(_05475_),
    .B1(_05488_),
    .Y(_00448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1293 ();
 sky130_fd_sc_hd__nand2_1 _16117_ (.A(net20),
    .B(_05475_),
    .Y(_05490_));
 sky130_fd_sc_hd__o21ai_0 _16118_ (.A1(_05192_),
    .A2(_05475_),
    .B1(_05490_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _16119_ (.A(net19),
    .B(_05475_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_0 _16120_ (.A1(_05204_),
    .A2(_05475_),
    .B1(_05491_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _16121_ (.A(net18),
    .B(_05475_),
    .Y(_05492_));
 sky130_fd_sc_hd__o21ai_0 _16122_ (.A1(_05214_),
    .A2(_05475_),
    .B1(_05492_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _16123_ (.A(net17),
    .B(_05475_),
    .Y(_05493_));
 sky130_fd_sc_hd__o21ai_0 _16124_ (.A1(_05221_),
    .A2(_05475_),
    .B1(_05493_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _16125_ (.A(net16),
    .B(_05475_),
    .Y(_05494_));
 sky130_fd_sc_hd__o21ai_0 _16126_ (.A1(_05228_),
    .A2(_05475_),
    .B1(_05494_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _16127_ (.A(net15),
    .B(_05475_),
    .Y(_05495_));
 sky130_fd_sc_hd__o21ai_0 _16128_ (.A1(_05238_),
    .A2(_05475_),
    .B1(_05495_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _16129_ (.A(net14),
    .B(_05475_),
    .Y(_05496_));
 sky130_fd_sc_hd__o21ai_0 _16130_ (.A1(_05247_),
    .A2(_05475_),
    .B1(_05496_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _16131_ (.A(net13),
    .B(_05475_),
    .Y(_05497_));
 sky130_fd_sc_hd__o21ai_0 _16132_ (.A1(_05258_),
    .A2(_05475_),
    .B1(_05497_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _16133_ (.A(net11),
    .B(_05475_),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_0 _16134_ (.A1(_05267_),
    .A2(_05475_),
    .B1(_05498_),
    .Y(_00426_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1292 ();
 sky130_fd_sc_hd__nand2_1 _16136_ (.A(net10),
    .B(_05475_),
    .Y(_05500_));
 sky130_fd_sc_hd__o21ai_0 _16137_ (.A1(_05280_),
    .A2(_05475_),
    .B1(_05500_),
    .Y(_00427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1291 ();
 sky130_fd_sc_hd__nand2_1 _16139_ (.A(net9),
    .B(_05475_),
    .Y(_05502_));
 sky130_fd_sc_hd__o21ai_0 _16140_ (.A1(_05291_),
    .A2(_05475_),
    .B1(_05502_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(net8),
    .B(_05475_),
    .Y(_05503_));
 sky130_fd_sc_hd__o21ai_0 _16142_ (.A1(_05301_),
    .A2(_05475_),
    .B1(_05503_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _16143_ (.A(net7),
    .B(_05475_),
    .Y(_05504_));
 sky130_fd_sc_hd__o21ai_0 _16144_ (.A1(_05309_),
    .A2(_05475_),
    .B1(_05504_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _16145_ (.A(net6),
    .B(_05475_),
    .Y(_05505_));
 sky130_fd_sc_hd__o21ai_0 _16146_ (.A1(_05320_),
    .A2(_05475_),
    .B1(_05505_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _16147_ (.A(net5),
    .B(_05475_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21ai_0 _16148_ (.A1(_05326_),
    .A2(_05475_),
    .B1(_05506_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _16149_ (.A(net4),
    .B(_05475_),
    .Y(_05507_));
 sky130_fd_sc_hd__o21ai_0 _16150_ (.A1(_05339_),
    .A2(_05475_),
    .B1(_05507_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _16151_ (.A(net3),
    .B(_05475_),
    .Y(_05508_));
 sky130_fd_sc_hd__o21ai_0 _16152_ (.A1(_05347_),
    .A2(_05475_),
    .B1(_05508_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _16153_ (.A(net2),
    .B(_05475_),
    .Y(_05509_));
 sky130_fd_sc_hd__o21ai_0 _16154_ (.A1(net538),
    .A2(_05475_),
    .B1(_05509_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _16155_ (.A(net782),
    .B(_05475_),
    .Y(_05510_));
 sky130_fd_sc_hd__o21ai_0 _16156_ (.A1(_05372_),
    .A2(_05475_),
    .B1(_05510_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _16157_ (.A(net781),
    .B(_05475_),
    .Y(_05511_));
 sky130_fd_sc_hd__o21ai_0 _16158_ (.A1(_05380_),
    .A2(_05475_),
    .B1(_05511_),
    .Y(_00438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1289 ();
 sky130_fd_sc_hd__a21oi_1 _16161_ (.A1(_09797_),
    .A2(_05474_),
    .B1(net780),
    .Y(_05514_));
 sky130_fd_sc_hd__a31oi_1 _16162_ (.A1(_09797_),
    .A2(net1134),
    .A3(_05474_),
    .B1(_05514_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _16163_ (.A(net779),
    .B(_05475_),
    .Y(_05515_));
 sky130_fd_sc_hd__o21ai_0 _16164_ (.A1(net1042),
    .A2(_05475_),
    .B1(_05515_),
    .Y(_00441_));
 sky130_fd_sc_hd__nor2b_4 _16165_ (.A(net1044),
    .B_N(_13529_),
    .Y(_05516_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1288 ();
 sky130_fd_sc_hd__nand2_8 _16167_ (.A(_09735_),
    .B(_05516_),
    .Y(_05518_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1286 ();
 sky130_fd_sc_hd__nand2_1 _16170_ (.A(net66),
    .B(_05518_),
    .Y(_05521_));
 sky130_fd_sc_hd__o21ai_0 _16171_ (.A1(_04790_),
    .A2(_05518_),
    .B1(_05521_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _16172_ (.A(net65),
    .B(_05518_),
    .Y(_05522_));
 sky130_fd_sc_hd__o21ai_0 _16173_ (.A1(_04794_),
    .A2(_05518_),
    .B1(_05522_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _16174_ (.A(net64),
    .B(_05518_),
    .Y(_05523_));
 sky130_fd_sc_hd__o21ai_0 _16175_ (.A1(_04801_),
    .A2(_05518_),
    .B1(_05523_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _16176_ (.A(net63),
    .B(_05518_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_0 _16177_ (.A1(_04808_),
    .A2(_05518_),
    .B1(_05524_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _16178_ (.A(net62),
    .B(_05518_),
    .Y(_05525_));
 sky130_fd_sc_hd__o21ai_0 _16179_ (.A1(_04817_),
    .A2(_05518_),
    .B1(_05525_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _16180_ (.A(net61),
    .B(_05518_),
    .Y(_05526_));
 sky130_fd_sc_hd__o21ai_0 _16181_ (.A1(_04826_),
    .A2(_05518_),
    .B1(_05526_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _16182_ (.A(net60),
    .B(_05518_),
    .Y(_05527_));
 sky130_fd_sc_hd__o21ai_0 _16183_ (.A1(_04834_),
    .A2(_05518_),
    .B1(_05527_),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _16184_ (.A(net59),
    .B(_05518_),
    .Y(_05528_));
 sky130_fd_sc_hd__o21ai_0 _16185_ (.A1(_04843_),
    .A2(_05518_),
    .B1(_05528_),
    .Y(_00478_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1285 ();
 sky130_fd_sc_hd__nand2_1 _16187_ (.A(net58),
    .B(_05518_),
    .Y(_05530_));
 sky130_fd_sc_hd__o21ai_0 _16188_ (.A1(_04852_),
    .A2(_05518_),
    .B1(_05530_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _16189_ (.A(net57),
    .B(_05518_),
    .Y(_05531_));
 sky130_fd_sc_hd__o21ai_0 _16190_ (.A1(_04860_),
    .A2(_05518_),
    .B1(_05531_),
    .Y(_00480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1284 ();
 sky130_fd_sc_hd__nand2_1 _16192_ (.A(net55),
    .B(_05518_),
    .Y(_05533_));
 sky130_fd_sc_hd__o21ai_0 _16193_ (.A1(_04871_),
    .A2(_05518_),
    .B1(_05533_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _16194_ (.A(net54),
    .B(_05518_),
    .Y(_05534_));
 sky130_fd_sc_hd__o21ai_0 _16195_ (.A1(_04883_),
    .A2(_05518_),
    .B1(_05534_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _16196_ (.A(net53),
    .B(_05518_),
    .Y(_05535_));
 sky130_fd_sc_hd__o21ai_0 _16197_ (.A1(_04892_),
    .A2(_05518_),
    .B1(_05535_),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _16198_ (.A(net52),
    .B(_05518_),
    .Y(_05536_));
 sky130_fd_sc_hd__o21ai_0 _16199_ (.A1(_04899_),
    .A2(_05518_),
    .B1(_05536_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _16200_ (.A(net51),
    .B(_05518_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_0 _16201_ (.A1(_04906_),
    .A2(_05518_),
    .B1(_05537_),
    .Y(_00454_));
 sky130_fd_sc_hd__nand2_1 _16202_ (.A(net50),
    .B(_05518_),
    .Y(_05538_));
 sky130_fd_sc_hd__o21ai_0 _16203_ (.A1(_04913_),
    .A2(_05518_),
    .B1(_05538_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _16204_ (.A(net49),
    .B(_05518_),
    .Y(_05539_));
 sky130_fd_sc_hd__o21ai_0 _16205_ (.A1(_04923_),
    .A2(_05518_),
    .B1(_05539_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _16206_ (.A(net48),
    .B(_05518_),
    .Y(_05540_));
 sky130_fd_sc_hd__o21ai_0 _16207_ (.A1(_04932_),
    .A2(_05518_),
    .B1(_05540_),
    .Y(_00457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1283 ();
 sky130_fd_sc_hd__nand2_1 _16209_ (.A(net47),
    .B(_05518_),
    .Y(_05542_));
 sky130_fd_sc_hd__o21ai_0 _16210_ (.A1(_04939_),
    .A2(_05518_),
    .B1(_05542_),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _16211_ (.A(net46),
    .B(_05518_),
    .Y(_05543_));
 sky130_fd_sc_hd__o21ai_0 _16212_ (.A1(_04951_),
    .A2(_05518_),
    .B1(_05543_),
    .Y(_00459_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1282 ();
 sky130_fd_sc_hd__nand2_1 _16214_ (.A(net44),
    .B(_05518_),
    .Y(_05545_));
 sky130_fd_sc_hd__o21ai_0 _16215_ (.A1(_04960_),
    .A2(_05518_),
    .B1(_05545_),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _16216_ (.A(net43),
    .B(_05518_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21ai_0 _16217_ (.A1(_04974_),
    .A2(_05518_),
    .B1(_05546_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _16218_ (.A(net42),
    .B(_05518_),
    .Y(_05547_));
 sky130_fd_sc_hd__o21ai_0 _16219_ (.A1(_04984_),
    .A2(_05518_),
    .B1(_05547_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _16220_ (.A(net41),
    .B(_05518_),
    .Y(_05548_));
 sky130_fd_sc_hd__o21ai_0 _16221_ (.A1(_04990_),
    .A2(_05518_),
    .B1(_05548_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _16222_ (.A(net40),
    .B(_05518_),
    .Y(_05549_));
 sky130_fd_sc_hd__o21ai_0 _16223_ (.A1(_05000_),
    .A2(_05518_),
    .B1(_05549_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _16224_ (.A(net39),
    .B(_05518_),
    .Y(_05550_));
 sky130_fd_sc_hd__o21ai_0 _16225_ (.A1(_05011_),
    .A2(_05518_),
    .B1(_05550_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _16226_ (.A(net38),
    .B(_05518_),
    .Y(_05551_));
 sky130_fd_sc_hd__o21ai_0 _16227_ (.A1(_05020_),
    .A2(_05518_),
    .B1(_05551_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _16228_ (.A(net37),
    .B(_05518_),
    .Y(_05552_));
 sky130_fd_sc_hd__o21ai_0 _16229_ (.A1(_05029_),
    .A2(_05518_),
    .B1(_05552_),
    .Y(_00468_));
 sky130_fd_sc_hd__nand2_1 _16230_ (.A(net36),
    .B(_05518_),
    .Y(_05553_));
 sky130_fd_sc_hd__o21ai_0 _16231_ (.A1(_05035_),
    .A2(_05518_),
    .B1(_05553_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _16232_ (.A(net35),
    .B(_05518_),
    .Y(_05554_));
 sky130_fd_sc_hd__o21ai_0 _16233_ (.A1(_05044_),
    .A2(_05518_),
    .B1(_05554_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _16234_ (.A(net33),
    .B(_05518_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21ai_0 _16235_ (.A1(_05060_),
    .A2(_05518_),
    .B1(_05555_),
    .Y(_00472_));
 sky130_fd_sc_hd__mux2i_1 _16236_ (.A0(_05113_),
    .A1(net32),
    .S(_05518_),
    .Y(_05556_));
 sky130_fd_sc_hd__o21ai_0 _16237_ (.A1(_05112_),
    .A2(_05518_),
    .B1(_05556_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2b_4 _16238_ (.A(net1044),
    .B_N(_13537_),
    .Y(_05557_));
 sky130_fd_sc_hd__nand2_8 _16239_ (.A(_09797_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1280 ();
 sky130_fd_sc_hd__nand2_1 _16242_ (.A(net102),
    .B(_05558_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21ai_0 _16243_ (.A1(_05118_),
    .A2(_05558_),
    .B1(_05561_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _16244_ (.A(net101),
    .B(_05558_),
    .Y(_05562_));
 sky130_fd_sc_hd__o21ai_0 _16245_ (.A1(_05122_),
    .A2(_05558_),
    .B1(_05562_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _16246_ (.A(net99),
    .B(_05558_),
    .Y(_05563_));
 sky130_fd_sc_hd__o21ai_0 _16247_ (.A1(_05126_),
    .A2(_05558_),
    .B1(_05563_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _16248_ (.A(net98),
    .B(_05558_),
    .Y(_05564_));
 sky130_fd_sc_hd__o21ai_0 _16249_ (.A1(_05132_),
    .A2(_05558_),
    .B1(_05564_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _16250_ (.A(net97),
    .B(_05558_),
    .Y(_05565_));
 sky130_fd_sc_hd__o21ai_0 _16251_ (.A1(_05140_),
    .A2(_05558_),
    .B1(_05565_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _16252_ (.A(net96),
    .B(_05558_),
    .Y(_05566_));
 sky130_fd_sc_hd__o21ai_0 _16253_ (.A1(_05149_),
    .A2(_05558_),
    .B1(_05566_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _16254_ (.A(net95),
    .B(_05558_),
    .Y(_05567_));
 sky130_fd_sc_hd__o21ai_0 _16255_ (.A1(_05157_),
    .A2(_05558_),
    .B1(_05567_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _16256_ (.A(net94),
    .B(_05558_),
    .Y(_05568_));
 sky130_fd_sc_hd__o21ai_0 _16257_ (.A1(_05166_),
    .A2(_05558_),
    .B1(_05568_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _16258_ (.A(net93),
    .B(_05558_),
    .Y(_05569_));
 sky130_fd_sc_hd__o21ai_0 _16259_ (.A1(_05173_),
    .A2(_05558_),
    .B1(_05569_),
    .Y(_00511_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1279 ();
 sky130_fd_sc_hd__nand2_1 _16261_ (.A(net92),
    .B(_05558_),
    .Y(_05571_));
 sky130_fd_sc_hd__o21ai_0 _16262_ (.A1(_05183_),
    .A2(_05558_),
    .B1(_05571_),
    .Y(_00512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1278 ();
 sky130_fd_sc_hd__nand2_1 _16264_ (.A(net91),
    .B(_05558_),
    .Y(_05573_));
 sky130_fd_sc_hd__o21ai_0 _16265_ (.A1(_05192_),
    .A2(_05558_),
    .B1(_05573_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _16266_ (.A(net90),
    .B(_05558_),
    .Y(_05574_));
 sky130_fd_sc_hd__o21ai_0 _16267_ (.A1(_05204_),
    .A2(_05558_),
    .B1(_05574_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _16268_ (.A(net88),
    .B(_05558_),
    .Y(_05575_));
 sky130_fd_sc_hd__o21ai_0 _16269_ (.A1(_05214_),
    .A2(_05558_),
    .B1(_05575_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _16270_ (.A(net87),
    .B(_05558_),
    .Y(_05576_));
 sky130_fd_sc_hd__o21ai_0 _16271_ (.A1(_05221_),
    .A2(_05558_),
    .B1(_05576_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _16272_ (.A(net86),
    .B(_05558_),
    .Y(_05577_));
 sky130_fd_sc_hd__o21ai_0 _16273_ (.A1(_05228_),
    .A2(_05558_),
    .B1(_05577_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _16274_ (.A(net85),
    .B(_05558_),
    .Y(_05578_));
 sky130_fd_sc_hd__o21ai_0 _16275_ (.A1(_05238_),
    .A2(_05558_),
    .B1(_05578_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _16276_ (.A(net84),
    .B(_05558_),
    .Y(_05579_));
 sky130_fd_sc_hd__o21ai_0 _16277_ (.A1(_05247_),
    .A2(_05558_),
    .B1(_05579_),
    .Y(_00488_));
 sky130_fd_sc_hd__nand2_1 _16278_ (.A(net83),
    .B(_05558_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ai_0 _16279_ (.A1(_05258_),
    .A2(_05558_),
    .B1(_05580_),
    .Y(_00489_));
 sky130_fd_sc_hd__nand2_1 _16280_ (.A(net82),
    .B(_05558_),
    .Y(_05581_));
 sky130_fd_sc_hd__o21ai_0 _16281_ (.A1(_05267_),
    .A2(_05558_),
    .B1(_05581_),
    .Y(_00490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1277 ();
 sky130_fd_sc_hd__nand2_1 _16283_ (.A(net81),
    .B(_05558_),
    .Y(_05583_));
 sky130_fd_sc_hd__o21ai_0 _16284_ (.A1(_05280_),
    .A2(_05558_),
    .B1(_05583_),
    .Y(_00491_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1276 ();
 sky130_fd_sc_hd__nand2_2 _16286_ (.A(net80),
    .B(_05558_),
    .Y(_05585_));
 sky130_fd_sc_hd__o21ai_0 _16287_ (.A1(_05291_),
    .A2(_05558_),
    .B1(_05585_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _16288_ (.A(net79),
    .B(_05558_),
    .Y(_05586_));
 sky130_fd_sc_hd__o21ai_0 _16289_ (.A1(_05301_),
    .A2(_05558_),
    .B1(_05586_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _16290_ (.A(net77),
    .B(_05558_),
    .Y(_05587_));
 sky130_fd_sc_hd__o21ai_0 _16291_ (.A1(_05309_),
    .A2(_05558_),
    .B1(_05587_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand2_1 _16292_ (.A(net76),
    .B(_05558_),
    .Y(_05588_));
 sky130_fd_sc_hd__o21ai_0 _16293_ (.A1(_05320_),
    .A2(_05558_),
    .B1(_05588_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _16294_ (.A(net75),
    .B(_05558_),
    .Y(_05589_));
 sky130_fd_sc_hd__o21ai_0 _16295_ (.A1(_05326_),
    .A2(_05558_),
    .B1(_05589_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _16296_ (.A(net74),
    .B(_05558_),
    .Y(_05590_));
 sky130_fd_sc_hd__o21ai_0 _16297_ (.A1(_05339_),
    .A2(_05558_),
    .B1(_05590_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _16298_ (.A(net73),
    .B(_05558_),
    .Y(_05591_));
 sky130_fd_sc_hd__o21ai_0 _16299_ (.A1(_05347_),
    .A2(_05558_),
    .B1(_05591_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _16300_ (.A(net72),
    .B(_05558_),
    .Y(_05592_));
 sky130_fd_sc_hd__o21ai_0 _16301_ (.A1(net538),
    .A2(_05558_),
    .B1(_05592_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _16302_ (.A(net71),
    .B(_05558_),
    .Y(_05593_));
 sky130_fd_sc_hd__o21ai_0 _16303_ (.A1(_05372_),
    .A2(_05558_),
    .B1(_05593_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _16304_ (.A(net70),
    .B(_05558_),
    .Y(_05594_));
 sky130_fd_sc_hd__o21ai_0 _16305_ (.A1(_05380_),
    .A2(_05558_),
    .B1(_05594_),
    .Y(_00502_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1275 ();
 sky130_fd_sc_hd__a21oi_1 _16307_ (.A1(_09797_),
    .A2(_05557_),
    .B1(net69),
    .Y(_05596_));
 sky130_fd_sc_hd__a31oi_1 _16308_ (.A1(_09797_),
    .A2(net1134),
    .A3(_05557_),
    .B1(_05596_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _16309_ (.A(net68),
    .B(_05558_),
    .Y(_05597_));
 sky130_fd_sc_hd__o21ai_0 _16310_ (.A1(net1042),
    .A2(_05558_),
    .B1(_05597_),
    .Y(_00505_));
 sky130_fd_sc_hd__nor2b_4 _16311_ (.A(net1044),
    .B_N(_13533_),
    .Y(_05598_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1274 ();
 sky130_fd_sc_hd__nand2_8 _16313_ (.A(_09735_),
    .B(_05598_),
    .Y(_05600_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1272 ();
 sky130_fd_sc_hd__nand2_1 _16316_ (.A(net138),
    .B(_05600_),
    .Y(_05603_));
 sky130_fd_sc_hd__o21ai_0 _16317_ (.A1(_04790_),
    .A2(_05600_),
    .B1(_05603_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _16318_ (.A(net137),
    .B(_05600_),
    .Y(_05604_));
 sky130_fd_sc_hd__o21ai_0 _16319_ (.A1(_04794_),
    .A2(_05600_),
    .B1(_05604_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _16320_ (.A(net136),
    .B(_05600_),
    .Y(_05605_));
 sky130_fd_sc_hd__o21ai_0 _16321_ (.A1(_04801_),
    .A2(_05600_),
    .B1(_05605_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _16322_ (.A(net135),
    .B(_05600_),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_0 _16323_ (.A1(_04808_),
    .A2(_05600_),
    .B1(_05606_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _16324_ (.A(net133),
    .B(_05600_),
    .Y(_05607_));
 sky130_fd_sc_hd__o21ai_0 _16325_ (.A1(_04817_),
    .A2(_05600_),
    .B1(_05607_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand2_1 _16326_ (.A(net132),
    .B(_05600_),
    .Y(_05608_));
 sky130_fd_sc_hd__o21ai_0 _16327_ (.A1(_04826_),
    .A2(_05600_),
    .B1(_05608_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(net131),
    .B(_05600_),
    .Y(_05609_));
 sky130_fd_sc_hd__o21ai_0 _16329_ (.A1(_04834_),
    .A2(_05600_),
    .B1(_05609_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _16330_ (.A(net130),
    .B(_05600_),
    .Y(_05610_));
 sky130_fd_sc_hd__o21ai_0 _16331_ (.A1(_04843_),
    .A2(_05600_),
    .B1(_05610_),
    .Y(_00542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1271 ();
 sky130_fd_sc_hd__nand2_1 _16333_ (.A(net129),
    .B(_05600_),
    .Y(_05612_));
 sky130_fd_sc_hd__o21ai_0 _16334_ (.A1(_04852_),
    .A2(_05600_),
    .B1(_05612_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _16335_ (.A(net128),
    .B(_05600_),
    .Y(_05613_));
 sky130_fd_sc_hd__o21ai_0 _16336_ (.A1(_04860_),
    .A2(_05600_),
    .B1(_05613_),
    .Y(_00544_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1270 ();
 sky130_fd_sc_hd__nand2_1 _16338_ (.A(net127),
    .B(_05600_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_0 _16339_ (.A1(_04871_),
    .A2(_05600_),
    .B1(_05615_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _16340_ (.A(net126),
    .B(_05600_),
    .Y(_05616_));
 sky130_fd_sc_hd__o21ai_0 _16341_ (.A1(_04883_),
    .A2(_05600_),
    .B1(_05616_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _16342_ (.A(net125),
    .B(_05600_),
    .Y(_05617_));
 sky130_fd_sc_hd__o21ai_0 _16343_ (.A1(_04892_),
    .A2(_05600_),
    .B1(_05617_),
    .Y(_00516_));
 sky130_fd_sc_hd__nand2_1 _16344_ (.A(net124),
    .B(_05600_),
    .Y(_05618_));
 sky130_fd_sc_hd__o21ai_0 _16345_ (.A1(_04899_),
    .A2(_05600_),
    .B1(_05618_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _16346_ (.A(net122),
    .B(_05600_),
    .Y(_05619_));
 sky130_fd_sc_hd__o21ai_0 _16347_ (.A1(_04906_),
    .A2(_05600_),
    .B1(_05619_),
    .Y(_00518_));
 sky130_fd_sc_hd__nand2_1 _16348_ (.A(net121),
    .B(_05600_),
    .Y(_05620_));
 sky130_fd_sc_hd__o21ai_0 _16349_ (.A1(_04913_),
    .A2(_05600_),
    .B1(_05620_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _16350_ (.A(net120),
    .B(_05600_),
    .Y(_05621_));
 sky130_fd_sc_hd__o21ai_0 _16351_ (.A1(_04923_),
    .A2(_05600_),
    .B1(_05621_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _16352_ (.A(net119),
    .B(_05600_),
    .Y(_05622_));
 sky130_fd_sc_hd__o21ai_0 _16353_ (.A1(_04932_),
    .A2(_05600_),
    .B1(_05622_),
    .Y(_00521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1269 ();
 sky130_fd_sc_hd__nand2_1 _16355_ (.A(net118),
    .B(_05600_),
    .Y(_05624_));
 sky130_fd_sc_hd__o21ai_0 _16356_ (.A1(_04939_),
    .A2(_05600_),
    .B1(_05624_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_1 _16357_ (.A(net117),
    .B(_05600_),
    .Y(_05625_));
 sky130_fd_sc_hd__o21ai_0 _16358_ (.A1(_04951_),
    .A2(_05600_),
    .B1(_05625_),
    .Y(_00523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1268 ();
 sky130_fd_sc_hd__nand2_1 _16360_ (.A(net116),
    .B(_05600_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21ai_0 _16361_ (.A1(_04960_),
    .A2(_05600_),
    .B1(_05627_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _16362_ (.A(net115),
    .B(_05600_),
    .Y(_05628_));
 sky130_fd_sc_hd__o21ai_0 _16363_ (.A1(_04974_),
    .A2(_05600_),
    .B1(_05628_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _16364_ (.A(net114),
    .B(_05600_),
    .Y(_05629_));
 sky130_fd_sc_hd__o21ai_0 _16365_ (.A1(_04984_),
    .A2(_05600_),
    .B1(_05629_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _16366_ (.A(net113),
    .B(_05600_),
    .Y(_05630_));
 sky130_fd_sc_hd__o21ai_0 _16367_ (.A1(_04990_),
    .A2(_05600_),
    .B1(_05630_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _16368_ (.A(net110),
    .B(_05600_),
    .Y(_05631_));
 sky130_fd_sc_hd__o21ai_0 _16369_ (.A1(_05000_),
    .A2(_05600_),
    .B1(_05631_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _16370_ (.A(net109),
    .B(_05600_),
    .Y(_05632_));
 sky130_fd_sc_hd__o21ai_0 _16371_ (.A1(_05011_),
    .A2(_05600_),
    .B1(_05632_),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _16372_ (.A(net108),
    .B(_05600_),
    .Y(_05633_));
 sky130_fd_sc_hd__o21ai_0 _16373_ (.A1(_05020_),
    .A2(_05600_),
    .B1(_05633_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _16374_ (.A(net107),
    .B(_05600_),
    .Y(_05634_));
 sky130_fd_sc_hd__o21ai_0 _16375_ (.A1(_05029_),
    .A2(_05600_),
    .B1(_05634_),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _16376_ (.A(net106),
    .B(_05600_),
    .Y(_05635_));
 sky130_fd_sc_hd__o21ai_0 _16377_ (.A1(_05035_),
    .A2(_05600_),
    .B1(_05635_),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2_1 _16378_ (.A(net105),
    .B(_05600_),
    .Y(_05636_));
 sky130_fd_sc_hd__o21ai_0 _16379_ (.A1(_05044_),
    .A2(_05600_),
    .B1(_05636_),
    .Y(_00534_));
 sky130_fd_sc_hd__nand2_1 _16380_ (.A(net104),
    .B(_05600_),
    .Y(_05637_));
 sky130_fd_sc_hd__o21ai_0 _16381_ (.A1(_05060_),
    .A2(_05600_),
    .B1(_05637_),
    .Y(_00536_));
 sky130_fd_sc_hd__mux2i_1 _16382_ (.A0(_05113_),
    .A1(net103),
    .S(_05600_),
    .Y(_05638_));
 sky130_fd_sc_hd__o21ai_0 _16383_ (.A1(_05112_),
    .A2(_05600_),
    .B1(_05638_),
    .Y(_00537_));
 sky130_fd_sc_hd__nor4_4 _16384_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(net1043),
    .D(_09803_),
    .Y(_05639_));
 sky130_fd_sc_hd__nor2_1 _16385_ (.A(net173),
    .B(net1073),
    .Y(_05640_));
 sky130_fd_sc_hd__a21oi_1 _16386_ (.A1(_05118_),
    .A2(net1073),
    .B1(_05640_),
    .Y(_00545_));
 sky130_fd_sc_hd__nor2_1 _16387_ (.A(net172),
    .B(net1073),
    .Y(_05641_));
 sky130_fd_sc_hd__a21oi_1 _16388_ (.A1(_05122_),
    .A2(net1073),
    .B1(_05641_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand2_8 _16389_ (.A(_09731_),
    .B(_09836_),
    .Y(_05642_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1266 ();
 sky130_fd_sc_hd__nand2_1 _16392_ (.A(net171),
    .B(_05642_),
    .Y(_05645_));
 sky130_fd_sc_hd__o21ai_0 _16393_ (.A1(_05126_),
    .A2(_05642_),
    .B1(_05645_),
    .Y(_00567_));
 sky130_fd_sc_hd__nor2_1 _16394_ (.A(net170),
    .B(net1073),
    .Y(_05646_));
 sky130_fd_sc_hd__a21oi_1 _16395_ (.A1(_05132_),
    .A2(net1073),
    .B1(_05646_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _16396_ (.A(net169),
    .B(_05642_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_0 _16397_ (.A1(_05140_),
    .A2(_05642_),
    .B1(_05647_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _16398_ (.A(net168),
    .B(_05642_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_0 _16399_ (.A1(_05149_),
    .A2(_05642_),
    .B1(_05648_),
    .Y(_00572_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1265 ();
 sky130_fd_sc_hd__nand2_1 _16401_ (.A(net166),
    .B(_05642_),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_0 _16402_ (.A1(_05157_),
    .A2(_05642_),
    .B1(_05650_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _16403_ (.A(net165),
    .B(_05642_),
    .Y(_05651_));
 sky130_fd_sc_hd__o21ai_0 _16404_ (.A1(_05166_),
    .A2(_05642_),
    .B1(_05651_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _16405_ (.A(net164),
    .B(_05642_),
    .Y(_05652_));
 sky130_fd_sc_hd__o21ai_0 _16406_ (.A1(_05173_),
    .A2(_05642_),
    .B1(_05652_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _16407_ (.A(net163),
    .B(_05642_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21ai_0 _16408_ (.A1(_05183_),
    .A2(_05642_),
    .B1(_05653_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _16409_ (.A(net162),
    .B(_05642_),
    .Y(_05654_));
 sky130_fd_sc_hd__o21ai_0 _16410_ (.A1(_05192_),
    .A2(_05642_),
    .B1(_05654_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _16411_ (.A(net161),
    .B(_05642_),
    .Y(_05655_));
 sky130_fd_sc_hd__o21ai_0 _16412_ (.A1(_05204_),
    .A2(_05642_),
    .B1(_05655_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _16413_ (.A(net160),
    .B(_05642_),
    .Y(_05656_));
 sky130_fd_sc_hd__o21ai_0 _16414_ (.A1(_05214_),
    .A2(_05642_),
    .B1(_05656_),
    .Y(_00548_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1264 ();
 sky130_fd_sc_hd__nand2_1 _16416_ (.A(net159),
    .B(_05642_),
    .Y(_05658_));
 sky130_fd_sc_hd__o21ai_0 _16417_ (.A1(_05221_),
    .A2(_05642_),
    .B1(_05658_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _16418_ (.A(net158),
    .B(_05642_),
    .Y(_05659_));
 sky130_fd_sc_hd__o21ai_0 _16419_ (.A1(_05228_),
    .A2(_05642_),
    .B1(_05659_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _16420_ (.A(net157),
    .B(_05642_),
    .Y(_05660_));
 sky130_fd_sc_hd__o21ai_0 _16421_ (.A1(_05238_),
    .A2(_05642_),
    .B1(_05660_),
    .Y(_00551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1263 ();
 sky130_fd_sc_hd__nand2_1 _16423_ (.A(net155),
    .B(_05642_),
    .Y(_05662_));
 sky130_fd_sc_hd__o21ai_0 _16424_ (.A1(_05247_),
    .A2(_05642_),
    .B1(_05662_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _16425_ (.A(net154),
    .B(_05642_),
    .Y(_05663_));
 sky130_fd_sc_hd__o21ai_0 _16426_ (.A1(_05258_),
    .A2(_05642_),
    .B1(_05663_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_1 _16427_ (.A(net153),
    .B(_05642_),
    .Y(_05664_));
 sky130_fd_sc_hd__o21ai_0 _16428_ (.A1(_05267_),
    .A2(_05642_),
    .B1(_05664_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _16429_ (.A(net152),
    .B(_05642_),
    .Y(_05665_));
 sky130_fd_sc_hd__o21ai_0 _16430_ (.A1(_05280_),
    .A2(_05642_),
    .B1(_05665_),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _16431_ (.A(net151),
    .B(_05642_),
    .Y(_05666_));
 sky130_fd_sc_hd__o21ai_0 _16432_ (.A1(_05291_),
    .A2(_05642_),
    .B1(_05666_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(net150),
    .B(_05642_),
    .Y(_05667_));
 sky130_fd_sc_hd__o21ai_0 _16434_ (.A1(_05301_),
    .A2(_05642_),
    .B1(_05667_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_1 _16435_ (.A(net149),
    .B(_05642_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21ai_0 _16436_ (.A1(_05309_),
    .A2(_05642_),
    .B1(_05668_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _16437_ (.A(net148),
    .B(_05642_),
    .Y(_05669_));
 sky130_fd_sc_hd__o21ai_0 _16438_ (.A1(_05320_),
    .A2(_05642_),
    .B1(_05669_),
    .Y(_00560_));
 sky130_fd_sc_hd__nand2_1 _16439_ (.A(net147),
    .B(_05642_),
    .Y(_05670_));
 sky130_fd_sc_hd__o21ai_0 _16440_ (.A1(_05326_),
    .A2(_05642_),
    .B1(_05670_),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_1 _16441_ (.A(net146),
    .B(_05642_),
    .Y(_05671_));
 sky130_fd_sc_hd__o21ai_0 _16442_ (.A1(_05339_),
    .A2(_05642_),
    .B1(_05671_),
    .Y(_00562_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(net144),
    .B(_05642_),
    .Y(_05672_));
 sky130_fd_sc_hd__o21ai_0 _16444_ (.A1(_05347_),
    .A2(_05642_),
    .B1(_05672_),
    .Y(_00563_));
 sky130_fd_sc_hd__nor2_1 _16445_ (.A(net143),
    .B(net1073),
    .Y(_05673_));
 sky130_fd_sc_hd__a21oi_1 _16446_ (.A1(net538),
    .A2(net1073),
    .B1(_05673_),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_1 _16447_ (.A(net142),
    .B(_05642_),
    .Y(_05674_));
 sky130_fd_sc_hd__o21ai_0 _16448_ (.A1(_05372_),
    .A2(_05642_),
    .B1(_05674_),
    .Y(_00565_));
 sky130_fd_sc_hd__nand2_1 _16449_ (.A(net141),
    .B(_05642_),
    .Y(_05675_));
 sky130_fd_sc_hd__o21ai_0 _16450_ (.A1(_05380_),
    .A2(_05642_),
    .B1(_05675_),
    .Y(_00566_));
 sky130_fd_sc_hd__nor2_1 _16451_ (.A(net140),
    .B(_05639_),
    .Y(_05676_));
 sky130_fd_sc_hd__a21oi_1 _16452_ (.A1(net1134),
    .A2(_05639_),
    .B1(_05676_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _16453_ (.A(net139),
    .B(_05642_),
    .Y(_05677_));
 sky130_fd_sc_hd__o21ai_0 _16454_ (.A1(net1042),
    .A2(_05642_),
    .B1(_05677_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_8 _16455_ (.A(_09739_),
    .B(_04784_),
    .Y(_05678_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1261 ();
 sky130_fd_sc_hd__nand2_1 _16458_ (.A(net208),
    .B(_05678_),
    .Y(_05681_));
 sky130_fd_sc_hd__o21ai_0 _16459_ (.A1(_04790_),
    .A2(_05678_),
    .B1(_05681_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _16460_ (.A(net207),
    .B(_05678_),
    .Y(_05682_));
 sky130_fd_sc_hd__o21ai_0 _16461_ (.A1(_04794_),
    .A2(_05678_),
    .B1(_05682_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _16462_ (.A(net206),
    .B(_05678_),
    .Y(_05683_));
 sky130_fd_sc_hd__o21ai_0 _16463_ (.A1(_04801_),
    .A2(_05678_),
    .B1(_05683_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _16464_ (.A(net205),
    .B(_05678_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21ai_0 _16465_ (.A1(_04808_),
    .A2(_05678_),
    .B1(_05684_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _16466_ (.A(net204),
    .B(_05678_),
    .Y(_05685_));
 sky130_fd_sc_hd__o21ai_0 _16467_ (.A1(_04817_),
    .A2(_05678_),
    .B1(_05685_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _16468_ (.A(net203),
    .B(_05678_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21ai_0 _16469_ (.A1(_04826_),
    .A2(_05678_),
    .B1(_05686_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _16470_ (.A(net202),
    .B(_05678_),
    .Y(_05687_));
 sky130_fd_sc_hd__o21ai_0 _16471_ (.A1(_04834_),
    .A2(_05678_),
    .B1(_05687_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _16472_ (.A(net201),
    .B(_05678_),
    .Y(_05688_));
 sky130_fd_sc_hd__o21ai_0 _16473_ (.A1(_04843_),
    .A2(_05678_),
    .B1(_05688_),
    .Y(_00606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1260 ();
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(net199),
    .B(_05678_),
    .Y(_05690_));
 sky130_fd_sc_hd__o21ai_0 _16476_ (.A1(_04852_),
    .A2(_05678_),
    .B1(_05690_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _16477_ (.A(net198),
    .B(_05678_),
    .Y(_05691_));
 sky130_fd_sc_hd__o21ai_0 _16478_ (.A1(_04860_),
    .A2(_05678_),
    .B1(_05691_),
    .Y(_00608_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1259 ();
 sky130_fd_sc_hd__nand2_1 _16480_ (.A(net197),
    .B(_05678_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_0 _16481_ (.A1(_04871_),
    .A2(_05678_),
    .B1(_05693_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _16482_ (.A(net196),
    .B(_05678_),
    .Y(_05694_));
 sky130_fd_sc_hd__o21ai_0 _16483_ (.A1(_04883_),
    .A2(_05678_),
    .B1(_05694_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _16484_ (.A(net195),
    .B(_05678_),
    .Y(_05695_));
 sky130_fd_sc_hd__o21ai_0 _16485_ (.A1(_04892_),
    .A2(_05678_),
    .B1(_05695_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_1 _16486_ (.A(net194),
    .B(_05678_),
    .Y(_05696_));
 sky130_fd_sc_hd__o21ai_0 _16487_ (.A1(_04899_),
    .A2(_05678_),
    .B1(_05696_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_1 _16488_ (.A(net193),
    .B(_05678_),
    .Y(_05697_));
 sky130_fd_sc_hd__o21ai_0 _16489_ (.A1(_04906_),
    .A2(_05678_),
    .B1(_05697_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _16490_ (.A(net192),
    .B(_05678_),
    .Y(_05698_));
 sky130_fd_sc_hd__o21ai_0 _16491_ (.A1(_04913_),
    .A2(_05678_),
    .B1(_05698_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _16492_ (.A(net191),
    .B(_05678_),
    .Y(_05699_));
 sky130_fd_sc_hd__o21ai_0 _16493_ (.A1(_04923_),
    .A2(_05678_),
    .B1(_05699_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _16494_ (.A(net190),
    .B(_05678_),
    .Y(_05700_));
 sky130_fd_sc_hd__o21ai_0 _16495_ (.A1(_04932_),
    .A2(_05678_),
    .B1(_05700_),
    .Y(_00585_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1258 ();
 sky130_fd_sc_hd__nand2_1 _16497_ (.A(net188),
    .B(_05678_),
    .Y(_05702_));
 sky130_fd_sc_hd__o21ai_0 _16498_ (.A1(_04939_),
    .A2(_05678_),
    .B1(_05702_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _16499_ (.A(net187),
    .B(_05678_),
    .Y(_05703_));
 sky130_fd_sc_hd__o21ai_0 _16500_ (.A1(_04951_),
    .A2(_05678_),
    .B1(_05703_),
    .Y(_00587_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1257 ();
 sky130_fd_sc_hd__nand2_1 _16502_ (.A(net186),
    .B(_05678_),
    .Y(_05705_));
 sky130_fd_sc_hd__o21ai_0 _16503_ (.A1(_04960_),
    .A2(_05678_),
    .B1(_05705_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _16504_ (.A(net185),
    .B(_05678_),
    .Y(_05706_));
 sky130_fd_sc_hd__o21ai_0 _16505_ (.A1(_04974_),
    .A2(_05678_),
    .B1(_05706_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _16506_ (.A(net184),
    .B(_05678_),
    .Y(_05707_));
 sky130_fd_sc_hd__o21ai_0 _16507_ (.A1(_04984_),
    .A2(_05678_),
    .B1(_05707_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand2_1 _16508_ (.A(net183),
    .B(_05678_),
    .Y(_05708_));
 sky130_fd_sc_hd__o21ai_0 _16509_ (.A1(_04990_),
    .A2(_05678_),
    .B1(_05708_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _16510_ (.A(net182),
    .B(_05678_),
    .Y(_05709_));
 sky130_fd_sc_hd__o21ai_0 _16511_ (.A1(_05000_),
    .A2(_05678_),
    .B1(_05709_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _16512_ (.A(net181),
    .B(_05678_),
    .Y(_05710_));
 sky130_fd_sc_hd__o21ai_0 _16513_ (.A1(_05011_),
    .A2(_05678_),
    .B1(_05710_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _16514_ (.A(net180),
    .B(_05678_),
    .Y(_05711_));
 sky130_fd_sc_hd__o21ai_0 _16515_ (.A1(_05020_),
    .A2(_05678_),
    .B1(_05711_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _16516_ (.A(net179),
    .B(_05678_),
    .Y(_05712_));
 sky130_fd_sc_hd__o21ai_0 _16517_ (.A1(_05029_),
    .A2(_05678_),
    .B1(_05712_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _16518_ (.A(net177),
    .B(_05678_),
    .Y(_05713_));
 sky130_fd_sc_hd__o21ai_0 _16519_ (.A1(_05035_),
    .A2(_05678_),
    .B1(_05713_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _16520_ (.A(net176),
    .B(_05678_),
    .Y(_05714_));
 sky130_fd_sc_hd__o21ai_0 _16521_ (.A1(_05044_),
    .A2(_05678_),
    .B1(_05714_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _16522_ (.A(net175),
    .B(_05678_),
    .Y(_05715_));
 sky130_fd_sc_hd__o21ai_0 _16523_ (.A1(_05060_),
    .A2(_05678_),
    .B1(_05715_),
    .Y(_00600_));
 sky130_fd_sc_hd__mux2i_1 _16524_ (.A0(_05113_),
    .A1(net174),
    .S(_05678_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_0 _16525_ (.A1(_05112_),
    .A2(_05678_),
    .B1(_05716_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_8 _16526_ (.A(_09784_),
    .B(_05115_),
    .Y(_05717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1255 ();
 sky130_fd_sc_hd__nand2_1 _16529_ (.A(net244),
    .B(_05717_),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ai_0 _16530_ (.A1(_05118_),
    .A2(_05717_),
    .B1(_05720_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _16531_ (.A(net243),
    .B(_05717_),
    .Y(_05721_));
 sky130_fd_sc_hd__o21ai_0 _16532_ (.A1(_05122_),
    .A2(_05717_),
    .B1(_05721_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _16533_ (.A(net242),
    .B(_05717_),
    .Y(_05722_));
 sky130_fd_sc_hd__o21ai_0 _16534_ (.A1(_05126_),
    .A2(_05717_),
    .B1(_05722_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _16535_ (.A(net241),
    .B(_05717_),
    .Y(_05723_));
 sky130_fd_sc_hd__o21ai_0 _16536_ (.A1(_05132_),
    .A2(_05717_),
    .B1(_05723_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _16537_ (.A(net240),
    .B(_05717_),
    .Y(_05724_));
 sky130_fd_sc_hd__o21ai_0 _16538_ (.A1(_05140_),
    .A2(_05717_),
    .B1(_05724_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _16539_ (.A(net239),
    .B(_05717_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_0 _16540_ (.A1(_05149_),
    .A2(_05717_),
    .B1(_05725_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _16541_ (.A(net238),
    .B(_05717_),
    .Y(_05726_));
 sky130_fd_sc_hd__o21ai_0 _16542_ (.A1(_05157_),
    .A2(_05717_),
    .B1(_05726_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _16543_ (.A(net237),
    .B(_05717_),
    .Y(_05727_));
 sky130_fd_sc_hd__o21ai_0 _16544_ (.A1(_05166_),
    .A2(_05717_),
    .B1(_05727_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _16545_ (.A(net236),
    .B(_05717_),
    .Y(_05728_));
 sky130_fd_sc_hd__o21ai_0 _16546_ (.A1(_05173_),
    .A2(_05717_),
    .B1(_05728_),
    .Y(_00639_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1254 ();
 sky130_fd_sc_hd__nand2_1 _16548_ (.A(net235),
    .B(_05717_),
    .Y(_05730_));
 sky130_fd_sc_hd__o21ai_0 _16549_ (.A1(_05183_),
    .A2(_05717_),
    .B1(_05730_),
    .Y(_00640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1253 ();
 sky130_fd_sc_hd__nand2_1 _16551_ (.A(net233),
    .B(_05717_),
    .Y(_05732_));
 sky130_fd_sc_hd__o21ai_0 _16552_ (.A1(_05192_),
    .A2(_05717_),
    .B1(_05732_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _16553_ (.A(net232),
    .B(_05717_),
    .Y(_05733_));
 sky130_fd_sc_hd__o21ai_0 _16554_ (.A1(_05204_),
    .A2(_05717_),
    .B1(_05733_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _16555_ (.A(net231),
    .B(_05717_),
    .Y(_05734_));
 sky130_fd_sc_hd__o21ai_0 _16556_ (.A1(_05214_),
    .A2(_05717_),
    .B1(_05734_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _16557_ (.A(net230),
    .B(_05717_),
    .Y(_05735_));
 sky130_fd_sc_hd__o21ai_0 _16558_ (.A1(_05221_),
    .A2(_05717_),
    .B1(_05735_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _16559_ (.A(net229),
    .B(_05717_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21ai_0 _16560_ (.A1(_05228_),
    .A2(_05717_),
    .B1(_05736_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _16561_ (.A(net228),
    .B(_05717_),
    .Y(_05737_));
 sky130_fd_sc_hd__o21ai_0 _16562_ (.A1(_05238_),
    .A2(_05717_),
    .B1(_05737_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _16563_ (.A(net227),
    .B(_05717_),
    .Y(_05738_));
 sky130_fd_sc_hd__o21ai_0 _16564_ (.A1(_05247_),
    .A2(_05717_),
    .B1(_05738_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _16565_ (.A(net226),
    .B(_05717_),
    .Y(_05739_));
 sky130_fd_sc_hd__o21ai_0 _16566_ (.A1(_05258_),
    .A2(_05717_),
    .B1(_05739_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _16567_ (.A(net225),
    .B(_05717_),
    .Y(_05740_));
 sky130_fd_sc_hd__o21ai_0 _16568_ (.A1(_05267_),
    .A2(_05717_),
    .B1(_05740_),
    .Y(_00618_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1252 ();
 sky130_fd_sc_hd__nand2_1 _16570_ (.A(net224),
    .B(_05717_),
    .Y(_05742_));
 sky130_fd_sc_hd__o21ai_0 _16571_ (.A1(_05280_),
    .A2(_05717_),
    .B1(_05742_),
    .Y(_00619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1251 ();
 sky130_fd_sc_hd__nand2_1 _16573_ (.A(net221),
    .B(_05717_),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ai_0 _16574_ (.A1(_05291_),
    .A2(_05717_),
    .B1(_05744_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _16575_ (.A(net220),
    .B(_05717_),
    .Y(_05745_));
 sky130_fd_sc_hd__o21ai_0 _16576_ (.A1(_05301_),
    .A2(_05717_),
    .B1(_05745_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _16577_ (.A(net219),
    .B(_05717_),
    .Y(_05746_));
 sky130_fd_sc_hd__o21ai_0 _16578_ (.A1(_05309_),
    .A2(_05717_),
    .B1(_05746_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _16579_ (.A(net218),
    .B(_05717_),
    .Y(_05747_));
 sky130_fd_sc_hd__o21ai_0 _16580_ (.A1(_05320_),
    .A2(_05717_),
    .B1(_05747_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _16581_ (.A(net217),
    .B(_05717_),
    .Y(_05748_));
 sky130_fd_sc_hd__o21ai_0 _16582_ (.A1(_05326_),
    .A2(_05717_),
    .B1(_05748_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _16583_ (.A(net216),
    .B(_05717_),
    .Y(_05749_));
 sky130_fd_sc_hd__o21ai_0 _16584_ (.A1(_05339_),
    .A2(_05717_),
    .B1(_05749_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _16585_ (.A(net215),
    .B(_05717_),
    .Y(_05750_));
 sky130_fd_sc_hd__o21ai_0 _16586_ (.A1(_05347_),
    .A2(_05717_),
    .B1(_05750_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _16587_ (.A(net214),
    .B(_05717_),
    .Y(_05751_));
 sky130_fd_sc_hd__o21ai_0 _16588_ (.A1(net538),
    .A2(_05717_),
    .B1(_05751_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _16589_ (.A(net213),
    .B(_05717_),
    .Y(_05752_));
 sky130_fd_sc_hd__o21ai_0 _16590_ (.A1(_05372_),
    .A2(_05717_),
    .B1(_05752_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _16591_ (.A(net212),
    .B(_05717_),
    .Y(_05753_));
 sky130_fd_sc_hd__o21ai_0 _16592_ (.A1(_05380_),
    .A2(_05717_),
    .B1(_05753_),
    .Y(_00630_));
 sky130_fd_sc_hd__a21oi_1 _16593_ (.A1(_09784_),
    .A2(_05115_),
    .B1(net210),
    .Y(_05754_));
 sky130_fd_sc_hd__a31oi_1 _16594_ (.A1(_09784_),
    .A2(_05115_),
    .A3(net1134),
    .B1(_05754_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _16595_ (.A(net209),
    .B(_05717_),
    .Y(_05755_));
 sky130_fd_sc_hd__o21ai_0 _16596_ (.A1(net1042),
    .A2(_05717_),
    .B1(_05755_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_8 _16597_ (.A(_09739_),
    .B(_05433_),
    .Y(_05756_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1249 ();
 sky130_fd_sc_hd__nand2_1 _16600_ (.A(net280),
    .B(_05756_),
    .Y(_05759_));
 sky130_fd_sc_hd__o21ai_0 _16601_ (.A1(_04790_),
    .A2(_05756_),
    .B1(_05759_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _16602_ (.A(net279),
    .B(_05756_),
    .Y(_05760_));
 sky130_fd_sc_hd__o21ai_0 _16603_ (.A1(_04794_),
    .A2(_05756_),
    .B1(_05760_),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _16604_ (.A(net277),
    .B(_05756_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_0 _16605_ (.A1(_04801_),
    .A2(_05756_),
    .B1(_05761_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2_1 _16606_ (.A(net276),
    .B(_05756_),
    .Y(_05762_));
 sky130_fd_sc_hd__o21ai_0 _16607_ (.A1(_04808_),
    .A2(_05756_),
    .B1(_05762_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _16608_ (.A(net275),
    .B(_05756_),
    .Y(_05763_));
 sky130_fd_sc_hd__o21ai_0 _16609_ (.A1(_04817_),
    .A2(_05756_),
    .B1(_05763_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _16610_ (.A(net274),
    .B(_05756_),
    .Y(_05764_));
 sky130_fd_sc_hd__o21ai_0 _16611_ (.A1(_04826_),
    .A2(_05756_),
    .B1(_05764_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _16612_ (.A(net273),
    .B(_05756_),
    .Y(_05765_));
 sky130_fd_sc_hd__o21ai_0 _16613_ (.A1(_04834_),
    .A2(_05756_),
    .B1(_05765_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _16614_ (.A(net272),
    .B(_05756_),
    .Y(_05766_));
 sky130_fd_sc_hd__o21ai_0 _16615_ (.A1(_04843_),
    .A2(_05756_),
    .B1(_05766_),
    .Y(_00190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1248 ();
 sky130_fd_sc_hd__nand2_1 _16617_ (.A(net271),
    .B(_05756_),
    .Y(_05768_));
 sky130_fd_sc_hd__o21ai_0 _16618_ (.A1(_04852_),
    .A2(_05756_),
    .B1(_05768_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _16619_ (.A(net270),
    .B(_05756_),
    .Y(_05769_));
 sky130_fd_sc_hd__o21ai_0 _16620_ (.A1(_04860_),
    .A2(_05756_),
    .B1(_05769_),
    .Y(_00192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1247 ();
 sky130_fd_sc_hd__nand2_1 _16622_ (.A(net269),
    .B(_05756_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_0 _16623_ (.A1(_04871_),
    .A2(_05756_),
    .B1(_05771_),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _16624_ (.A(net268),
    .B(_05756_),
    .Y(_05772_));
 sky130_fd_sc_hd__o21ai_0 _16625_ (.A1(_04883_),
    .A2(_05756_),
    .B1(_05772_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _16626_ (.A(net266),
    .B(_05756_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21ai_0 _16627_ (.A1(_04892_),
    .A2(_05756_),
    .B1(_05773_),
    .Y(_00164_));
 sky130_fd_sc_hd__nand2_1 _16628_ (.A(net265),
    .B(_05756_),
    .Y(_05774_));
 sky130_fd_sc_hd__o21ai_0 _16629_ (.A1(_04899_),
    .A2(_05756_),
    .B1(_05774_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _16630_ (.A(net264),
    .B(_05756_),
    .Y(_05775_));
 sky130_fd_sc_hd__o21ai_0 _16631_ (.A1(_04906_),
    .A2(_05756_),
    .B1(_05775_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand2_1 _16632_ (.A(net263),
    .B(_05756_),
    .Y(_05776_));
 sky130_fd_sc_hd__o21ai_0 _16633_ (.A1(_04913_),
    .A2(_05756_),
    .B1(_05776_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _16634_ (.A(net262),
    .B(_05756_),
    .Y(_05777_));
 sky130_fd_sc_hd__o21ai_0 _16635_ (.A1(_04923_),
    .A2(_05756_),
    .B1(_05777_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _16636_ (.A(net261),
    .B(_05756_),
    .Y(_05778_));
 sky130_fd_sc_hd__o21ai_0 _16637_ (.A1(_04932_),
    .A2(_05756_),
    .B1(_05778_),
    .Y(_00169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1246 ();
 sky130_fd_sc_hd__nand2_1 _16639_ (.A(net260),
    .B(_05756_),
    .Y(_05780_));
 sky130_fd_sc_hd__o21ai_0 _16640_ (.A1(_04939_),
    .A2(_05756_),
    .B1(_05780_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_1 _16641_ (.A(net259),
    .B(_05756_),
    .Y(_05781_));
 sky130_fd_sc_hd__o21ai_0 _16642_ (.A1(_04951_),
    .A2(_05756_),
    .B1(_05781_),
    .Y(_00171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1245 ();
 sky130_fd_sc_hd__nand2_1 _16644_ (.A(net258),
    .B(_05756_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21ai_0 _16645_ (.A1(_04960_),
    .A2(_05756_),
    .B1(_05783_),
    .Y(_00173_));
 sky130_fd_sc_hd__nand2_1 _16646_ (.A(net257),
    .B(_05756_),
    .Y(_05784_));
 sky130_fd_sc_hd__o21ai_0 _16647_ (.A1(_04974_),
    .A2(_05756_),
    .B1(_05784_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _16648_ (.A(net255),
    .B(_05756_),
    .Y(_05785_));
 sky130_fd_sc_hd__o21ai_0 _16649_ (.A1(_04984_),
    .A2(_05756_),
    .B1(_05785_),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _16650_ (.A(net254),
    .B(_05756_),
    .Y(_05786_));
 sky130_fd_sc_hd__o21ai_0 _16651_ (.A1(_04990_),
    .A2(_05756_),
    .B1(_05786_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand2_1 _16652_ (.A(net253),
    .B(_05756_),
    .Y(_05787_));
 sky130_fd_sc_hd__o21ai_0 _16653_ (.A1(_05000_),
    .A2(_05756_),
    .B1(_05787_),
    .Y(_00177_));
 sky130_fd_sc_hd__nand2_1 _16654_ (.A(net252),
    .B(_05756_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21ai_0 _16655_ (.A1(_05011_),
    .A2(_05756_),
    .B1(_05788_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _16656_ (.A(net251),
    .B(_05756_),
    .Y(_05789_));
 sky130_fd_sc_hd__o21ai_0 _16657_ (.A1(_05020_),
    .A2(_05756_),
    .B1(_05789_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _16658_ (.A(net250),
    .B(_05756_),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ai_0 _16659_ (.A1(_05029_),
    .A2(_05756_),
    .B1(_05790_),
    .Y(_00180_));
 sky130_fd_sc_hd__nand2_1 _16660_ (.A(net249),
    .B(_05756_),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_0 _16661_ (.A1(_05035_),
    .A2(_05756_),
    .B1(_05791_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _16662_ (.A(net248),
    .B(_05756_),
    .Y(_05792_));
 sky130_fd_sc_hd__o21ai_0 _16663_ (.A1(_05044_),
    .A2(_05756_),
    .B1(_05792_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _16664_ (.A(net247),
    .B(_05756_),
    .Y(_05793_));
 sky130_fd_sc_hd__o21ai_0 _16665_ (.A1(_05060_),
    .A2(_05756_),
    .B1(_05793_),
    .Y(_00184_));
 sky130_fd_sc_hd__mux2i_1 _16666_ (.A0(_05113_),
    .A1(net246),
    .S(_05756_),
    .Y(_05794_));
 sky130_fd_sc_hd__o21ai_0 _16667_ (.A1(_05112_),
    .A2(_05756_),
    .B1(_05794_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_8 _16668_ (.A(_09784_),
    .B(_05474_),
    .Y(_05795_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1243 ();
 sky130_fd_sc_hd__nand2_1 _16671_ (.A(net586),
    .B(_05795_),
    .Y(_05798_));
 sky130_fd_sc_hd__o21ai_0 _16672_ (.A1(_05118_),
    .A2(_05795_),
    .B1(_05798_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _16673_ (.A(net585),
    .B(_05795_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ai_0 _16674_ (.A1(_05122_),
    .A2(_05795_),
    .B1(_05799_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _16675_ (.A(net584),
    .B(_05795_),
    .Y(_05800_));
 sky130_fd_sc_hd__o21ai_0 _16676_ (.A1(_05126_),
    .A2(_05795_),
    .B1(_05800_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _16677_ (.A(net583),
    .B(_05795_),
    .Y(_05801_));
 sky130_fd_sc_hd__o21ai_0 _16678_ (.A1(_05132_),
    .A2(_05795_),
    .B1(_05801_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _16679_ (.A(net581),
    .B(_05795_),
    .Y(_05802_));
 sky130_fd_sc_hd__o21ai_0 _16680_ (.A1(_05140_),
    .A2(_05795_),
    .B1(_05802_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _16681_ (.A(net580),
    .B(_05795_),
    .Y(_05803_));
 sky130_fd_sc_hd__o21ai_0 _16682_ (.A1(_05149_),
    .A2(_05795_),
    .B1(_05803_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _16683_ (.A(net579),
    .B(_05795_),
    .Y(_05804_));
 sky130_fd_sc_hd__o21ai_0 _16684_ (.A1(_05157_),
    .A2(_05795_),
    .B1(_05804_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _16685_ (.A(net578),
    .B(_05795_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_0 _16686_ (.A1(_05166_),
    .A2(_05795_),
    .B1(_05805_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _16687_ (.A(net577),
    .B(_05795_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21ai_0 _16688_ (.A1(_05173_),
    .A2(_05795_),
    .B1(_05806_),
    .Y(_00223_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1242 ();
 sky130_fd_sc_hd__nand2_2 _16690_ (.A(net576),
    .B(_05795_),
    .Y(_05808_));
 sky130_fd_sc_hd__o21ai_0 _16691_ (.A1(_05183_),
    .A2(_05795_),
    .B1(_05808_),
    .Y(_00224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1241 ();
 sky130_fd_sc_hd__nand2_1 _16693_ (.A(net575),
    .B(_05795_),
    .Y(_05810_));
 sky130_fd_sc_hd__o21ai_0 _16694_ (.A1(_05192_),
    .A2(_05795_),
    .B1(_05810_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _16695_ (.A(net574),
    .B(_05795_),
    .Y(_05811_));
 sky130_fd_sc_hd__o21ai_0 _16696_ (.A1(_05204_),
    .A2(_05795_),
    .B1(_05811_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _16697_ (.A(net573),
    .B(_05795_),
    .Y(_05812_));
 sky130_fd_sc_hd__o21ai_0 _16698_ (.A1(_05214_),
    .A2(_05795_),
    .B1(_05812_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _16699_ (.A(net572),
    .B(_05795_),
    .Y(_05813_));
 sky130_fd_sc_hd__o21ai_0 _16700_ (.A1(_05221_),
    .A2(_05795_),
    .B1(_05813_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand2_1 _16701_ (.A(net570),
    .B(_05795_),
    .Y(_05814_));
 sky130_fd_sc_hd__o21ai_0 _16702_ (.A1(_05228_),
    .A2(_05795_),
    .B1(_05814_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _16703_ (.A(net569),
    .B(_05795_),
    .Y(_05815_));
 sky130_fd_sc_hd__o21ai_0 _16704_ (.A1(_05238_),
    .A2(_05795_),
    .B1(_05815_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _16705_ (.A(net568),
    .B(_05795_),
    .Y(_05816_));
 sky130_fd_sc_hd__o21ai_0 _16706_ (.A1(_05247_),
    .A2(_05795_),
    .B1(_05816_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _16707_ (.A(net567),
    .B(_05795_),
    .Y(_05817_));
 sky130_fd_sc_hd__o21ai_0 _16708_ (.A1(_05258_),
    .A2(_05795_),
    .B1(_05817_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _16709_ (.A(net566),
    .B(_05795_),
    .Y(_05818_));
 sky130_fd_sc_hd__o21ai_0 _16710_ (.A1(_05267_),
    .A2(_05795_),
    .B1(_05818_),
    .Y(_00202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1240 ();
 sky130_fd_sc_hd__nand2_1 _16712_ (.A(net565),
    .B(_05795_),
    .Y(_05820_));
 sky130_fd_sc_hd__o21ai_0 _16713_ (.A1(_05280_),
    .A2(_05795_),
    .B1(_05820_),
    .Y(_00203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1239 ();
 sky130_fd_sc_hd__nand2_1 _16715_ (.A(net564),
    .B(_05795_),
    .Y(_05822_));
 sky130_fd_sc_hd__o21ai_0 _16716_ (.A1(_05291_),
    .A2(_05795_),
    .B1(_05822_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _16717_ (.A(net563),
    .B(_05795_),
    .Y(_05823_));
 sky130_fd_sc_hd__o21ai_0 _16718_ (.A1(_05301_),
    .A2(_05795_),
    .B1(_05823_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _16719_ (.A(net562),
    .B(_05795_),
    .Y(_05824_));
 sky130_fd_sc_hd__o21ai_0 _16720_ (.A1(_05309_),
    .A2(_05795_),
    .B1(_05824_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_1 _16721_ (.A(net561),
    .B(_05795_),
    .Y(_05825_));
 sky130_fd_sc_hd__o21ai_0 _16722_ (.A1(_05320_),
    .A2(_05795_),
    .B1(_05825_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _16723_ (.A(net288),
    .B(_05795_),
    .Y(_05826_));
 sky130_fd_sc_hd__o21ai_0 _16724_ (.A1(_05326_),
    .A2(_05795_),
    .B1(_05826_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _16725_ (.A(net287),
    .B(_05795_),
    .Y(_05827_));
 sky130_fd_sc_hd__o21ai_0 _16726_ (.A1(_05339_),
    .A2(_05795_),
    .B1(_05827_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _16727_ (.A(net286),
    .B(_05795_),
    .Y(_05828_));
 sky130_fd_sc_hd__o21ai_0 _16728_ (.A1(_05347_),
    .A2(_05795_),
    .B1(_05828_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _16729_ (.A(net285),
    .B(_05795_),
    .Y(_05829_));
 sky130_fd_sc_hd__o21ai_0 _16730_ (.A1(net538),
    .A2(_05795_),
    .B1(_05829_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _16731_ (.A(net284),
    .B(_05795_),
    .Y(_05830_));
 sky130_fd_sc_hd__o21ai_0 _16732_ (.A1(_05372_),
    .A2(_05795_),
    .B1(_05830_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _16733_ (.A(net283),
    .B(_05795_),
    .Y(_05831_));
 sky130_fd_sc_hd__o21ai_0 _16734_ (.A1(_05380_),
    .A2(_05795_),
    .B1(_05831_),
    .Y(_00214_));
 sky130_fd_sc_hd__a21oi_1 _16735_ (.A1(_09784_),
    .A2(_05474_),
    .B1(net282),
    .Y(_05832_));
 sky130_fd_sc_hd__a31oi_1 _16736_ (.A1(_09784_),
    .A2(net1134),
    .A3(_05474_),
    .B1(_05832_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _16737_ (.A(net281),
    .B(_05795_),
    .Y(_05833_));
 sky130_fd_sc_hd__o21ai_0 _16738_ (.A1(net1042),
    .A2(_05795_),
    .B1(_05833_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_8 _16739_ (.A(_09739_),
    .B(_05516_),
    .Y(_05834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1237 ();
 sky130_fd_sc_hd__nand2_1 _16742_ (.A(net622),
    .B(_05834_),
    .Y(_05837_));
 sky130_fd_sc_hd__o21ai_0 _16743_ (.A1(_04790_),
    .A2(_05834_),
    .B1(_05837_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _16744_ (.A(net621),
    .B(_05834_),
    .Y(_05838_));
 sky130_fd_sc_hd__o21ai_0 _16745_ (.A1(_04794_),
    .A2(_05834_),
    .B1(_05838_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _16746_ (.A(net620),
    .B(_05834_),
    .Y(_05839_));
 sky130_fd_sc_hd__o21ai_0 _16747_ (.A1(_04801_),
    .A2(_05834_),
    .B1(_05839_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _16748_ (.A(net619),
    .B(_05834_),
    .Y(_05840_));
 sky130_fd_sc_hd__o21ai_0 _16749_ (.A1(_04808_),
    .A2(_05834_),
    .B1(_05840_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _16750_ (.A(net618),
    .B(_05834_),
    .Y(_05841_));
 sky130_fd_sc_hd__o21ai_0 _16751_ (.A1(_04817_),
    .A2(_05834_),
    .B1(_05841_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(net617),
    .B(_05834_),
    .Y(_05842_));
 sky130_fd_sc_hd__o21ai_0 _16753_ (.A1(_04826_),
    .A2(_05834_),
    .B1(_05842_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _16754_ (.A(net615),
    .B(_05834_),
    .Y(_05843_));
 sky130_fd_sc_hd__o21ai_0 _16755_ (.A1(_04834_),
    .A2(_05834_),
    .B1(_05843_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _16756_ (.A(net614),
    .B(_05834_),
    .Y(_05844_));
 sky130_fd_sc_hd__o21ai_0 _16757_ (.A1(_04843_),
    .A2(_05834_),
    .B1(_05844_),
    .Y(_00254_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1236 ();
 sky130_fd_sc_hd__nand2_1 _16759_ (.A(net613),
    .B(_05834_),
    .Y(_05846_));
 sky130_fd_sc_hd__o21ai_0 _16760_ (.A1(_04852_),
    .A2(_05834_),
    .B1(_05846_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _16761_ (.A(net612),
    .B(_05834_),
    .Y(_05847_));
 sky130_fd_sc_hd__o21ai_0 _16762_ (.A1(_04860_),
    .A2(_05834_),
    .B1(_05847_),
    .Y(_00256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1235 ();
 sky130_fd_sc_hd__nand2_1 _16764_ (.A(net611),
    .B(_05834_),
    .Y(_05849_));
 sky130_fd_sc_hd__o21ai_0 _16765_ (.A1(_04871_),
    .A2(_05834_),
    .B1(_05849_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _16766_ (.A(net610),
    .B(_05834_),
    .Y(_05850_));
 sky130_fd_sc_hd__o21ai_0 _16767_ (.A1(_04883_),
    .A2(_05834_),
    .B1(_05850_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _16768_ (.A(net609),
    .B(_05834_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_0 _16769_ (.A1(_04892_),
    .A2(_05834_),
    .B1(_05851_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _16770_ (.A(net608),
    .B(_05834_),
    .Y(_05852_));
 sky130_fd_sc_hd__o21ai_0 _16771_ (.A1(_04899_),
    .A2(_05834_),
    .B1(_05852_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _16772_ (.A(net607),
    .B(_05834_),
    .Y(_05853_));
 sky130_fd_sc_hd__o21ai_0 _16773_ (.A1(_04906_),
    .A2(_05834_),
    .B1(_05853_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _16774_ (.A(net606),
    .B(_05834_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_0 _16775_ (.A1(_04913_),
    .A2(_05834_),
    .B1(_05854_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _16776_ (.A(net603),
    .B(_05834_),
    .Y(_05855_));
 sky130_fd_sc_hd__o21ai_0 _16777_ (.A1(_04923_),
    .A2(_05834_),
    .B1(_05855_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _16778_ (.A(net602),
    .B(_05834_),
    .Y(_05856_));
 sky130_fd_sc_hd__o21ai_0 _16779_ (.A1(_04932_),
    .A2(_05834_),
    .B1(_05856_),
    .Y(_00233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1234 ();
 sky130_fd_sc_hd__nand2_1 _16781_ (.A(net601),
    .B(_05834_),
    .Y(_05858_));
 sky130_fd_sc_hd__o21ai_0 _16782_ (.A1(_04939_),
    .A2(_05834_),
    .B1(_05858_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _16783_ (.A(net600),
    .B(_05834_),
    .Y(_05859_));
 sky130_fd_sc_hd__o21ai_0 _16784_ (.A1(_04951_),
    .A2(_05834_),
    .B1(_05859_),
    .Y(_00235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1233 ();
 sky130_fd_sc_hd__nand2_1 _16786_ (.A(net599),
    .B(_05834_),
    .Y(_05861_));
 sky130_fd_sc_hd__o21ai_0 _16787_ (.A1(_04960_),
    .A2(_05834_),
    .B1(_05861_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _16788_ (.A(net598),
    .B(_05834_),
    .Y(_05862_));
 sky130_fd_sc_hd__o21ai_0 _16789_ (.A1(_04974_),
    .A2(_05834_),
    .B1(_05862_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _16790_ (.A(net597),
    .B(_05834_),
    .Y(_05863_));
 sky130_fd_sc_hd__o21ai_0 _16791_ (.A1(_04984_),
    .A2(_05834_),
    .B1(_05863_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _16792_ (.A(net596),
    .B(_05834_),
    .Y(_05864_));
 sky130_fd_sc_hd__o21ai_0 _16793_ (.A1(_04990_),
    .A2(_05834_),
    .B1(_05864_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _16794_ (.A(net595),
    .B(_05834_),
    .Y(_05865_));
 sky130_fd_sc_hd__o21ai_0 _16795_ (.A1(_05000_),
    .A2(_05834_),
    .B1(_05865_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _16796_ (.A(net594),
    .B(_05834_),
    .Y(_05866_));
 sky130_fd_sc_hd__o21ai_0 _16797_ (.A1(_05011_),
    .A2(_05834_),
    .B1(_05866_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _16798_ (.A(net592),
    .B(_05834_),
    .Y(_05867_));
 sky130_fd_sc_hd__o21ai_0 _16799_ (.A1(_05020_),
    .A2(_05834_),
    .B1(_05867_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _16800_ (.A(net591),
    .B(_05834_),
    .Y(_05868_));
 sky130_fd_sc_hd__o21ai_0 _16801_ (.A1(_05029_),
    .A2(_05834_),
    .B1(_05868_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _16802_ (.A(net590),
    .B(_05834_),
    .Y(_05869_));
 sky130_fd_sc_hd__o21ai_0 _16803_ (.A1(_05035_),
    .A2(_05834_),
    .B1(_05869_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _16804_ (.A(net589),
    .B(_05834_),
    .Y(_05870_));
 sky130_fd_sc_hd__o21ai_0 _16805_ (.A1(_05044_),
    .A2(_05834_),
    .B1(_05870_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(net588),
    .B(_05834_),
    .Y(_05871_));
 sky130_fd_sc_hd__o21ai_0 _16807_ (.A1(_05060_),
    .A2(_05834_),
    .B1(_05871_),
    .Y(_00248_));
 sky130_fd_sc_hd__mux2i_1 _16808_ (.A0(_05113_),
    .A1(net587),
    .S(_05834_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21ai_0 _16809_ (.A1(_05112_),
    .A2(_05834_),
    .B1(_05872_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_8 _16810_ (.A(_09784_),
    .B(_05557_),
    .Y(_05873_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1231 ();
 sky130_fd_sc_hd__nand2_1 _16813_ (.A(net657),
    .B(_05873_),
    .Y(_05876_));
 sky130_fd_sc_hd__o21ai_0 _16814_ (.A1(_05118_),
    .A2(_05873_),
    .B1(_05876_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _16815_ (.A(net656),
    .B(_05873_),
    .Y(_05877_));
 sky130_fd_sc_hd__o21ai_0 _16816_ (.A1(_05122_),
    .A2(_05873_),
    .B1(_05877_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _16817_ (.A(net655),
    .B(_05873_),
    .Y(_05878_));
 sky130_fd_sc_hd__o21ai_0 _16818_ (.A1(_05126_),
    .A2(_05873_),
    .B1(_05878_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _16819_ (.A(net654),
    .B(_05873_),
    .Y(_05879_));
 sky130_fd_sc_hd__o21ai_0 _16820_ (.A1(_05132_),
    .A2(_05873_),
    .B1(_05879_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(net653),
    .B(_05873_),
    .Y(_05880_));
 sky130_fd_sc_hd__o21ai_0 _16822_ (.A1(_05140_),
    .A2(_05873_),
    .B1(_05880_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _16823_ (.A(net652),
    .B(_05873_),
    .Y(_05881_));
 sky130_fd_sc_hd__o21ai_0 _16824_ (.A1(_05149_),
    .A2(_05873_),
    .B1(_05881_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _16825_ (.A(net651),
    .B(_05873_),
    .Y(_05882_));
 sky130_fd_sc_hd__o21ai_0 _16826_ (.A1(_05157_),
    .A2(_05873_),
    .B1(_05882_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _16827_ (.A(net650),
    .B(_05873_),
    .Y(_05883_));
 sky130_fd_sc_hd__o21ai_0 _16828_ (.A1(_05166_),
    .A2(_05873_),
    .B1(_05883_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _16829_ (.A(net648),
    .B(_05873_),
    .Y(_05884_));
 sky130_fd_sc_hd__o21ai_0 _16830_ (.A1(_05173_),
    .A2(_05873_),
    .B1(_05884_),
    .Y(_00287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1230 ();
 sky130_fd_sc_hd__nand2_1 _16832_ (.A(net647),
    .B(_05873_),
    .Y(_05886_));
 sky130_fd_sc_hd__o21ai_0 _16833_ (.A1(_05183_),
    .A2(_05873_),
    .B1(_05886_),
    .Y(_00288_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1229 ();
 sky130_fd_sc_hd__nand2_1 _16835_ (.A(net646),
    .B(_05873_),
    .Y(_05888_));
 sky130_fd_sc_hd__o21ai_0 _16836_ (.A1(_05192_),
    .A2(_05873_),
    .B1(_05888_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _16837_ (.A(net645),
    .B(_05873_),
    .Y(_05889_));
 sky130_fd_sc_hd__o21ai_0 _16838_ (.A1(_05204_),
    .A2(_05873_),
    .B1(_05889_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _16839_ (.A(net644),
    .B(_05873_),
    .Y(_05890_));
 sky130_fd_sc_hd__o21ai_0 _16840_ (.A1(_05214_),
    .A2(_05873_),
    .B1(_05890_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _16841_ (.A(net643),
    .B(_05873_),
    .Y(_05891_));
 sky130_fd_sc_hd__o21ai_0 _16842_ (.A1(_05221_),
    .A2(_05873_),
    .B1(_05891_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _16843_ (.A(net642),
    .B(_05873_),
    .Y(_05892_));
 sky130_fd_sc_hd__o21ai_0 _16844_ (.A1(_05228_),
    .A2(_05873_),
    .B1(_05892_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _16845_ (.A(net641),
    .B(_05873_),
    .Y(_05893_));
 sky130_fd_sc_hd__o21ai_0 _16846_ (.A1(_05238_),
    .A2(_05873_),
    .B1(_05893_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _16847_ (.A(net640),
    .B(_05873_),
    .Y(_05894_));
 sky130_fd_sc_hd__o21ai_0 _16848_ (.A1(_05247_),
    .A2(_05873_),
    .B1(_05894_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _16849_ (.A(net639),
    .B(_05873_),
    .Y(_05895_));
 sky130_fd_sc_hd__o21ai_0 _16850_ (.A1(_05258_),
    .A2(_05873_),
    .B1(_05895_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _16851_ (.A(net637),
    .B(_05873_),
    .Y(_05896_));
 sky130_fd_sc_hd__o21ai_0 _16852_ (.A1(_05267_),
    .A2(_05873_),
    .B1(_05896_),
    .Y(_00266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1228 ();
 sky130_fd_sc_hd__nand2_1 _16854_ (.A(net636),
    .B(_05873_),
    .Y(_05898_));
 sky130_fd_sc_hd__o21ai_0 _16855_ (.A1(_05280_),
    .A2(_05873_),
    .B1(_05898_),
    .Y(_00267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1227 ();
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(net635),
    .B(_05873_),
    .Y(_05900_));
 sky130_fd_sc_hd__o21ai_0 _16858_ (.A1(_05291_),
    .A2(_05873_),
    .B1(_05900_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _16859_ (.A(net634),
    .B(_05873_),
    .Y(_05901_));
 sky130_fd_sc_hd__o21ai_0 _16860_ (.A1(_05301_),
    .A2(_05873_),
    .B1(_05901_),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _16861_ (.A(net633),
    .B(_05873_),
    .Y(_05902_));
 sky130_fd_sc_hd__o21ai_0 _16862_ (.A1(_05309_),
    .A2(_05873_),
    .B1(_05902_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _16863_ (.A(net632),
    .B(_05873_),
    .Y(_05903_));
 sky130_fd_sc_hd__o21ai_0 _16864_ (.A1(_05320_),
    .A2(_05873_),
    .B1(_05903_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _16865_ (.A(net631),
    .B(_05873_),
    .Y(_05904_));
 sky130_fd_sc_hd__o21ai_0 _16866_ (.A1(_05326_),
    .A2(_05873_),
    .B1(_05904_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(net630),
    .B(_05873_),
    .Y(_05905_));
 sky130_fd_sc_hd__o21ai_0 _16868_ (.A1(_05339_),
    .A2(_05873_),
    .B1(_05905_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _16869_ (.A(net629),
    .B(_05873_),
    .Y(_05906_));
 sky130_fd_sc_hd__o21ai_0 _16870_ (.A1(_05347_),
    .A2(_05873_),
    .B1(_05906_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _16871_ (.A(net628),
    .B(_05873_),
    .Y(_05907_));
 sky130_fd_sc_hd__o21ai_0 _16872_ (.A1(net538),
    .A2(_05873_),
    .B1(_05907_),
    .Y(_00276_));
 sky130_fd_sc_hd__nand2_1 _16873_ (.A(net626),
    .B(_05873_),
    .Y(_05908_));
 sky130_fd_sc_hd__o21ai_0 _16874_ (.A1(_05372_),
    .A2(_05873_),
    .B1(_05908_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _16875_ (.A(net625),
    .B(_05873_),
    .Y(_05909_));
 sky130_fd_sc_hd__o21ai_0 _16876_ (.A1(_05380_),
    .A2(_05873_),
    .B1(_05909_),
    .Y(_00278_));
 sky130_fd_sc_hd__a21oi_1 _16877_ (.A1(_09784_),
    .A2(_05557_),
    .B1(net624),
    .Y(_05910_));
 sky130_fd_sc_hd__a31oi_1 _16878_ (.A1(_09784_),
    .A2(net1134),
    .A3(_05557_),
    .B1(_05910_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _16879_ (.A(net623),
    .B(_05873_),
    .Y(_05911_));
 sky130_fd_sc_hd__o21ai_0 _16880_ (.A1(net1042),
    .A2(_05873_),
    .B1(_05911_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_8 _16881_ (.A(_09739_),
    .B(_05598_),
    .Y(_05912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1225 ();
 sky130_fd_sc_hd__nand2_1 _16884_ (.A(net692),
    .B(_05912_),
    .Y(_05915_));
 sky130_fd_sc_hd__o21ai_0 _16885_ (.A1(_04790_),
    .A2(_05912_),
    .B1(_05915_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _16886_ (.A(net691),
    .B(_05912_),
    .Y(_05916_));
 sky130_fd_sc_hd__o21ai_0 _16887_ (.A1(_04794_),
    .A2(_05912_),
    .B1(_05916_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _16888_ (.A(net690),
    .B(_05912_),
    .Y(_05917_));
 sky130_fd_sc_hd__o21ai_0 _16889_ (.A1(_04801_),
    .A2(_05912_),
    .B1(_05917_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _16890_ (.A(net689),
    .B(_05912_),
    .Y(_05918_));
 sky130_fd_sc_hd__o21ai_0 _16891_ (.A1(_04808_),
    .A2(_05912_),
    .B1(_05918_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(net688),
    .B(_05912_),
    .Y(_05919_));
 sky130_fd_sc_hd__o21ai_0 _16893_ (.A1(_04817_),
    .A2(_05912_),
    .B1(_05919_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _16894_ (.A(net687),
    .B(_05912_),
    .Y(_05920_));
 sky130_fd_sc_hd__o21ai_0 _16895_ (.A1(_04826_),
    .A2(_05912_),
    .B1(_05920_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _16896_ (.A(net686),
    .B(_05912_),
    .Y(_05921_));
 sky130_fd_sc_hd__o21ai_0 _16897_ (.A1(_04834_),
    .A2(_05912_),
    .B1(_05921_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _16898_ (.A(net685),
    .B(_05912_),
    .Y(_05922_));
 sky130_fd_sc_hd__o21ai_0 _16899_ (.A1(_04843_),
    .A2(_05912_),
    .B1(_05922_),
    .Y(_00318_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1224 ();
 sky130_fd_sc_hd__nand2_1 _16901_ (.A(net684),
    .B(_05912_),
    .Y(_05924_));
 sky130_fd_sc_hd__o21ai_0 _16902_ (.A1(_04852_),
    .A2(_05912_),
    .B1(_05924_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _16903_ (.A(net683),
    .B(_05912_),
    .Y(_05925_));
 sky130_fd_sc_hd__o21ai_0 _16904_ (.A1(_04860_),
    .A2(_05912_),
    .B1(_05925_),
    .Y(_00320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1223 ();
 sky130_fd_sc_hd__nand2_1 _16906_ (.A(net681),
    .B(_05912_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21ai_0 _16907_ (.A1(_04871_),
    .A2(_05912_),
    .B1(_05927_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _16908_ (.A(net680),
    .B(_05912_),
    .Y(_05928_));
 sky130_fd_sc_hd__o21ai_0 _16909_ (.A1(_04883_),
    .A2(_05912_),
    .B1(_05928_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _16910_ (.A(net679),
    .B(_05912_),
    .Y(_05929_));
 sky130_fd_sc_hd__o21ai_0 _16911_ (.A1(_04892_),
    .A2(_05912_),
    .B1(_05929_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _16912_ (.A(net678),
    .B(_05912_),
    .Y(_05930_));
 sky130_fd_sc_hd__o21ai_0 _16913_ (.A1(_04899_),
    .A2(_05912_),
    .B1(_05930_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _16914_ (.A(net677),
    .B(_05912_),
    .Y(_05931_));
 sky130_fd_sc_hd__o21ai_0 _16915_ (.A1(_04906_),
    .A2(_05912_),
    .B1(_05931_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _16916_ (.A(net676),
    .B(_05912_),
    .Y(_05932_));
 sky130_fd_sc_hd__o21ai_0 _16917_ (.A1(_04913_),
    .A2(_05912_),
    .B1(_05932_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _16918_ (.A(net675),
    .B(_05912_),
    .Y(_05933_));
 sky130_fd_sc_hd__o21ai_0 _16919_ (.A1(_04923_),
    .A2(_05912_),
    .B1(_05933_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _16920_ (.A(net674),
    .B(_05912_),
    .Y(_05934_));
 sky130_fd_sc_hd__o21ai_0 _16921_ (.A1(_04932_),
    .A2(_05912_),
    .B1(_05934_),
    .Y(_00297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1222 ();
 sky130_fd_sc_hd__nand2_1 _16923_ (.A(net673),
    .B(_05912_),
    .Y(_05936_));
 sky130_fd_sc_hd__o21ai_0 _16924_ (.A1(_04939_),
    .A2(_05912_),
    .B1(_05936_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _16925_ (.A(net672),
    .B(_05912_),
    .Y(_05937_));
 sky130_fd_sc_hd__o21ai_0 _16926_ (.A1(_04951_),
    .A2(_05912_),
    .B1(_05937_),
    .Y(_00299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1221 ();
 sky130_fd_sc_hd__nand2_1 _16928_ (.A(net670),
    .B(_05912_),
    .Y(_05939_));
 sky130_fd_sc_hd__o21ai_0 _16929_ (.A1(_04960_),
    .A2(_05912_),
    .B1(_05939_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _16930_ (.A(net669),
    .B(_05912_),
    .Y(_05940_));
 sky130_fd_sc_hd__o21ai_0 _16931_ (.A1(_04974_),
    .A2(_05912_),
    .B1(_05940_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _16932_ (.A(net668),
    .B(_05912_),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_0 _16933_ (.A1(_04984_),
    .A2(_05912_),
    .B1(_05941_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _16934_ (.A(net667),
    .B(_05912_),
    .Y(_05942_));
 sky130_fd_sc_hd__o21ai_0 _16935_ (.A1(_04990_),
    .A2(_05912_),
    .B1(_05942_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _16936_ (.A(net666),
    .B(_05912_),
    .Y(_05943_));
 sky130_fd_sc_hd__o21ai_0 _16937_ (.A1(_05000_),
    .A2(_05912_),
    .B1(_05943_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _16938_ (.A(net665),
    .B(_05912_),
    .Y(_05944_));
 sky130_fd_sc_hd__o21ai_0 _16939_ (.A1(_05011_),
    .A2(_05912_),
    .B1(_05944_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _16940_ (.A(net664),
    .B(_05912_),
    .Y(_05945_));
 sky130_fd_sc_hd__o21ai_0 _16941_ (.A1(_05020_),
    .A2(_05912_),
    .B1(_05945_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _16942_ (.A(net663),
    .B(_05912_),
    .Y(_05946_));
 sky130_fd_sc_hd__o21ai_0 _16943_ (.A1(_05029_),
    .A2(_05912_),
    .B1(_05946_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _16944_ (.A(net662),
    .B(_05912_),
    .Y(_05947_));
 sky130_fd_sc_hd__o21ai_0 _16945_ (.A1(_05035_),
    .A2(_05912_),
    .B1(_05947_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand2_1 _16946_ (.A(net661),
    .B(_05912_),
    .Y(_05948_));
 sky130_fd_sc_hd__o21ai_0 _16947_ (.A1(_05044_),
    .A2(_05912_),
    .B1(_05948_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _16948_ (.A(net659),
    .B(_05912_),
    .Y(_05949_));
 sky130_fd_sc_hd__o21ai_0 _16949_ (.A1(_05060_),
    .A2(_05912_),
    .B1(_05949_),
    .Y(_00312_));
 sky130_fd_sc_hd__mux2i_1 _16950_ (.A0(_05113_),
    .A1(net658),
    .S(_05912_),
    .Y(_05950_));
 sky130_fd_sc_hd__o21ai_0 _16951_ (.A1(_05112_),
    .A2(_05912_),
    .B1(_05950_),
    .Y(_00313_));
 sky130_fd_sc_hd__nor2b_4 _16952_ (.A(net1044),
    .B_N(_13541_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand2_8 _16953_ (.A(_09784_),
    .B(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1219 ();
 sky130_fd_sc_hd__nand2_1 _16956_ (.A(net729),
    .B(_05952_),
    .Y(_05955_));
 sky130_fd_sc_hd__o21ai_0 _16957_ (.A1(_05118_),
    .A2(_05952_),
    .B1(_05955_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _16958_ (.A(net728),
    .B(_05952_),
    .Y(_05956_));
 sky130_fd_sc_hd__o21ai_0 _16959_ (.A1(_05122_),
    .A2(_05952_),
    .B1(_05956_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _16960_ (.A(net726),
    .B(_05952_),
    .Y(_05957_));
 sky130_fd_sc_hd__o21ai_0 _16961_ (.A1(_05126_),
    .A2(_05952_),
    .B1(_05957_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _16962_ (.A(net725),
    .B(_05952_),
    .Y(_05958_));
 sky130_fd_sc_hd__o21ai_0 _16963_ (.A1(_05132_),
    .A2(_05952_),
    .B1(_05958_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _16964_ (.A(net724),
    .B(_05952_),
    .Y(_05959_));
 sky130_fd_sc_hd__o21ai_0 _16965_ (.A1(_05140_),
    .A2(_05952_),
    .B1(_05959_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _16966_ (.A(net723),
    .B(_05952_),
    .Y(_05960_));
 sky130_fd_sc_hd__o21ai_0 _16967_ (.A1(_05149_),
    .A2(_05952_),
    .B1(_05960_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(net722),
    .B(_05952_),
    .Y(_05961_));
 sky130_fd_sc_hd__o21ai_0 _16969_ (.A1(_05157_),
    .A2(_05952_),
    .B1(_05961_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(net721),
    .B(_05952_),
    .Y(_05962_));
 sky130_fd_sc_hd__o21ai_0 _16971_ (.A1(_05166_),
    .A2(_05952_),
    .B1(_05962_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _16972_ (.A(net720),
    .B(_05952_),
    .Y(_05963_));
 sky130_fd_sc_hd__o21ai_0 _16973_ (.A1(_05173_),
    .A2(_05952_),
    .B1(_05963_),
    .Y(_00351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1218 ();
 sky130_fd_sc_hd__nand2_1 _16975_ (.A(net719),
    .B(_05952_),
    .Y(_05965_));
 sky130_fd_sc_hd__o21ai_0 _16976_ (.A1(_05183_),
    .A2(_05952_),
    .B1(_05965_),
    .Y(_00352_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1217 ();
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(net718),
    .B(_05952_),
    .Y(_05967_));
 sky130_fd_sc_hd__o21ai_0 _16979_ (.A1(_05192_),
    .A2(_05952_),
    .B1(_05967_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _16980_ (.A(net717),
    .B(_05952_),
    .Y(_05968_));
 sky130_fd_sc_hd__o21ai_0 _16981_ (.A1(_05204_),
    .A2(_05952_),
    .B1(_05968_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _16982_ (.A(net714),
    .B(_05952_),
    .Y(_05969_));
 sky130_fd_sc_hd__o21ai_0 _16983_ (.A1(_05214_),
    .A2(_05952_),
    .B1(_05969_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(net713),
    .B(_05952_),
    .Y(_05970_));
 sky130_fd_sc_hd__o21ai_0 _16985_ (.A1(_05221_),
    .A2(_05952_),
    .B1(_05970_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _16986_ (.A(net712),
    .B(_05952_),
    .Y(_05971_));
 sky130_fd_sc_hd__o21ai_0 _16987_ (.A1(_05228_),
    .A2(_05952_),
    .B1(_05971_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _16988_ (.A(net711),
    .B(_05952_),
    .Y(_05972_));
 sky130_fd_sc_hd__o21ai_0 _16989_ (.A1(_05238_),
    .A2(_05952_),
    .B1(_05972_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _16990_ (.A(net710),
    .B(_05952_),
    .Y(_05973_));
 sky130_fd_sc_hd__o21ai_0 _16991_ (.A1(_05247_),
    .A2(_05952_),
    .B1(_05973_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _16992_ (.A(net709),
    .B(_05952_),
    .Y(_05974_));
 sky130_fd_sc_hd__o21ai_0 _16993_ (.A1(_05258_),
    .A2(_05952_),
    .B1(_05974_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _16994_ (.A(net708),
    .B(_05952_),
    .Y(_05975_));
 sky130_fd_sc_hd__o21ai_0 _16995_ (.A1(_05267_),
    .A2(_05952_),
    .B1(_05975_),
    .Y(_00330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1216 ();
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(net707),
    .B(_05952_),
    .Y(_05977_));
 sky130_fd_sc_hd__o21ai_0 _16998_ (.A1(_05280_),
    .A2(_05952_),
    .B1(_05977_),
    .Y(_00331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1215 ();
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(net706),
    .B(_05952_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21ai_0 _17001_ (.A1(_05291_),
    .A2(_05952_),
    .B1(_05979_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _17002_ (.A(net705),
    .B(_05952_),
    .Y(_05980_));
 sky130_fd_sc_hd__o21ai_0 _17003_ (.A1(_05301_),
    .A2(_05952_),
    .B1(_05980_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _17004_ (.A(net703),
    .B(_05952_),
    .Y(_05981_));
 sky130_fd_sc_hd__o21ai_0 _17005_ (.A1(_05309_),
    .A2(_05952_),
    .B1(_05981_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _17006_ (.A(net702),
    .B(_05952_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21ai_0 _17007_ (.A1(_05320_),
    .A2(_05952_),
    .B1(_05982_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _17008_ (.A(net701),
    .B(_05952_),
    .Y(_05983_));
 sky130_fd_sc_hd__o21ai_0 _17009_ (.A1(_05326_),
    .A2(_05952_),
    .B1(_05983_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _17010_ (.A(net700),
    .B(_05952_),
    .Y(_05984_));
 sky130_fd_sc_hd__o21ai_0 _17011_ (.A1(_05339_),
    .A2(_05952_),
    .B1(_05984_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(net699),
    .B(_05952_),
    .Y(_05985_));
 sky130_fd_sc_hd__o21ai_0 _17013_ (.A1(_05347_),
    .A2(_05952_),
    .B1(_05985_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _17014_ (.A(net698),
    .B(_05952_),
    .Y(_05986_));
 sky130_fd_sc_hd__o21ai_0 _17015_ (.A1(net538),
    .A2(_05952_),
    .B1(_05986_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_1 _17016_ (.A(net697),
    .B(_05952_),
    .Y(_05987_));
 sky130_fd_sc_hd__o21ai_0 _17017_ (.A1(_05372_),
    .A2(_05952_),
    .B1(_05987_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(net696),
    .B(_05952_),
    .Y(_05988_));
 sky130_fd_sc_hd__o21ai_0 _17019_ (.A1(_05380_),
    .A2(_05952_),
    .B1(_05988_),
    .Y(_00342_));
 sky130_fd_sc_hd__a21oi_1 _17020_ (.A1(_09784_),
    .A2(_05951_),
    .B1(net695),
    .Y(_05989_));
 sky130_fd_sc_hd__a31oi_1 _17021_ (.A1(_09784_),
    .A2(net1134),
    .A3(_05951_),
    .B1(_05989_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _17022_ (.A(net694),
    .B(_05952_),
    .Y(_05990_));
 sky130_fd_sc_hd__o21ai_0 _17023_ (.A1(net1042),
    .A2(_05952_),
    .B1(_05990_),
    .Y(_00345_));
 sky130_fd_sc_hd__or2_0 _17024_ (.A(\hash.reset ),
    .B(\hash.CA2.f_dash[0] ),
    .X(_12653_));
 sky130_fd_sc_hd__inv_1 _17025_ (.A(_12653_),
    .Y(_00875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1214 ();
 sky130_fd_sc_hd__nor2_1 _17027_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[0] ),
    .Y(_00843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1208 ();
 sky130_fd_sc_hd__clkinvlp_4 _17034_ (.A(_12109_),
    .Y(_05998_));
 sky130_fd_sc_hd__nor2_2 _17035_ (.A(net349),
    .B(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__inv_1 _17036_ (.A(_05999_),
    .Y(\hash.CA1.S0.X[2] ));
 sky130_fd_sc_hd__xnor2_1 _17037_ (.A(_13544_),
    .B(_05999_),
    .Y(_00680_));
 sky130_fd_sc_hd__xor2_2 _17038_ (.A(_12108_),
    .B(_13255_),
    .X(_06000_));
 sky130_fd_sc_hd__nor2_4 _17039_ (.A(net349),
    .B(_06000_),
    .Y(\hash.CA1.S0.X[3] ));
 sky130_fd_sc_hd__inv_1 _17040_ (.A(_00658_),
    .Y(\hash.CA1.S0.X[0] ));
 sky130_fd_sc_hd__or3_4 _17041_ (.A(_13241_),
    .B(_05998_),
    .C(\hash.CA1.S0.X[0] ),
    .X(_06001_));
 sky130_fd_sc_hd__xor2_1 _17042_ (.A(\hash.CA1.S0.X[3] ),
    .B(_06001_),
    .X(_00683_));
 sky130_fd_sc_hd__clkinv_16 _17043_ (.A(net349),
    .Y(_06002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1204 ();
 sky130_fd_sc_hd__a21o_4 _17048_ (.A1(_13240_),
    .A2(_13248_),
    .B1(_13247_),
    .X(_06007_));
 sky130_fd_sc_hd__a21oi_1 _17049_ (.A1(_13255_),
    .A2(_06007_),
    .B1(_13254_),
    .Y(_06008_));
 sky130_fd_sc_hd__xnor2_2 _17050_ (.A(_13262_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__and2_4 _17051_ (.A(_06002_),
    .B(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1203 ();
 sky130_fd_sc_hd__a211oi_1 _17053_ (.A1(_13544_),
    .A2(_12109_),
    .B1(_06000_),
    .C1(net349),
    .Y(_06011_));
 sky130_fd_sc_hd__xor2_1 _17054_ (.A(_06010_),
    .B(_06011_),
    .X(_00684_));
 sky130_fd_sc_hd__nor2b_2 _17055_ (.A(_12108_),
    .B_N(_13255_),
    .Y(_06012_));
 sky130_fd_sc_hd__o21a_1 _17056_ (.A1(_13254_),
    .A2(_06012_),
    .B1(_13262_),
    .X(_06013_));
 sky130_fd_sc_hd__o21ai_2 _17057_ (.A1(_13261_),
    .A2(_06013_),
    .B1(_13269_),
    .Y(_06014_));
 sky130_fd_sc_hd__or3_4 _17058_ (.A(_13269_),
    .B(_13261_),
    .C(_06013_),
    .X(_06015_));
 sky130_fd_sc_hd__a21oi_4 _17059_ (.A1(_06014_),
    .A2(_06015_),
    .B1(net349),
    .Y(_06016_));
 sky130_fd_sc_hd__clkinvlp_2 _17060_ (.A(_06016_),
    .Y(\hash.CA1.S0.X[5] ));
 sky130_fd_sc_hd__nand4_1 _17061_ (.A(_06002_),
    .B(\hash.CA1.S0.X[3] ),
    .C(_06001_),
    .D(_06009_),
    .Y(_06017_));
 sky130_fd_sc_hd__xnor2_1 _17062_ (.A(_06016_),
    .B(_06017_),
    .Y(_00685_));
 sky130_fd_sc_hd__nor2_1 _17063_ (.A(net349),
    .B(_13276_),
    .Y(_06018_));
 sky130_fd_sc_hd__nor2b_1 _17064_ (.A(net349),
    .B_N(_13276_),
    .Y(_06019_));
 sky130_fd_sc_hd__or2_4 _17065_ (.A(_13254_),
    .B(_13261_),
    .X(_06020_));
 sky130_fd_sc_hd__a21oi_2 _17066_ (.A1(_13255_),
    .A2(_06007_),
    .B1(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__o21ai_2 _17067_ (.A1(_13262_),
    .A2(_13261_),
    .B1(_13269_),
    .Y(_06022_));
 sky130_fd_sc_hd__o21bai_2 _17068_ (.A1(_06021_),
    .A2(_06022_),
    .B1_N(_13268_),
    .Y(_06023_));
 sky130_fd_sc_hd__mux2_8 _17069_ (.A0(_06018_),
    .A1(_06019_),
    .S(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__inv_4 _17070_ (.A(_06024_),
    .Y(\hash.CA1.S0.X[6] ));
 sky130_fd_sc_hd__nand3_1 _17071_ (.A(_06002_),
    .B(_06009_),
    .C(_06011_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2_1 _17072_ (.A(_06016_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__xnor2_1 _17073_ (.A(\hash.CA1.S0.X[6] ),
    .B(_06026_),
    .Y(_00686_));
 sky130_fd_sc_hd__o21a_1 _17074_ (.A1(_13262_),
    .A2(_13261_),
    .B1(_13269_),
    .X(_06027_));
 sky130_fd_sc_hd__o211a_2 _17075_ (.A1(_06012_),
    .A2(_06020_),
    .B1(_06027_),
    .C1(_13276_),
    .X(_06028_));
 sky130_fd_sc_hd__a21o_4 _17076_ (.A1(_13276_),
    .A2(_13268_),
    .B1(_13275_),
    .X(_06029_));
 sky130_fd_sc_hd__or3_4 _17077_ (.A(_13283_),
    .B(_06028_),
    .C(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__o21ai_2 _17078_ (.A1(_06028_),
    .A2(_06029_),
    .B1(_13283_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand3_4 _17079_ (.A(_06002_),
    .B(_06030_),
    .C(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__inv_4 _17080_ (.A(_06032_),
    .Y(\hash.CA1.S0.X[7] ));
 sky130_fd_sc_hd__a31oi_2 _17081_ (.A1(_06016_),
    .A2(_06017_),
    .A3(_06024_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__nand3_1 _17082_ (.A(_06016_),
    .B(_06017_),
    .C(_06024_),
    .Y(_06034_));
 sky130_fd_sc_hd__nor2_1 _17083_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__nor2_1 _17084_ (.A(_06033_),
    .B(_06035_),
    .Y(_00687_));
 sky130_fd_sc_hd__nor2_1 _17085_ (.A(net350),
    .B(_13290_),
    .Y(_06036_));
 sky130_fd_sc_hd__nor2b_1 _17086_ (.A(net349),
    .B_N(_13290_),
    .Y(_06037_));
 sky130_fd_sc_hd__nor2_1 _17087_ (.A(_13268_),
    .B(_13275_),
    .Y(_06038_));
 sky130_fd_sc_hd__o21ai_0 _17088_ (.A1(_06021_),
    .A2(_06022_),
    .B1(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__nor2_1 _17089_ (.A(_13276_),
    .B(_13275_),
    .Y(_06040_));
 sky130_fd_sc_hd__inv_1 _17090_ (.A(_06040_),
    .Y(_06041_));
 sky130_fd_sc_hd__a31oi_2 _17091_ (.A1(_13283_),
    .A2(_06039_),
    .A3(_06041_),
    .B1(_13282_),
    .Y(_06042_));
 sky130_fd_sc_hd__mux2_8 _17092_ (.A0(_06036_),
    .A1(_06037_),
    .S(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1202 ();
 sky130_fd_sc_hd__a31oi_2 _17094_ (.A1(_06016_),
    .A2(_06024_),
    .A3(_06025_),
    .B1(_06032_),
    .Y(_06044_));
 sky130_fd_sc_hd__xor2_1 _17095_ (.A(_06043_),
    .B(_06044_),
    .X(_00688_));
 sky130_fd_sc_hd__o211ai_1 _17096_ (.A1(_06012_),
    .A2(_06020_),
    .B1(_06027_),
    .C1(_13276_),
    .Y(_06045_));
 sky130_fd_sc_hd__nor3_2 _17097_ (.A(_13282_),
    .B(_13289_),
    .C(_06029_),
    .Y(_06046_));
 sky130_fd_sc_hd__o21a_1 _17098_ (.A1(_13283_),
    .A2(_13282_),
    .B1(_13290_),
    .X(_06047_));
 sky130_fd_sc_hd__nor2_1 _17099_ (.A(_13289_),
    .B(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__a21oi_1 _17100_ (.A1(_06045_),
    .A2(_06046_),
    .B1(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__xnor2_2 _17101_ (.A(_13297_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_8 _17102_ (.A(_06002_),
    .B(_06050_),
    .Y(\hash.CA1.S0.X[9] ));
 sky130_fd_sc_hd__nand2_1 _17103_ (.A(_06033_),
    .B(_06043_),
    .Y(_06051_));
 sky130_fd_sc_hd__xor2_1 _17104_ (.A(\hash.CA1.S0.X[9] ),
    .B(_06051_),
    .X(_00689_));
 sky130_fd_sc_hd__a21oi_2 _17105_ (.A1(_13297_),
    .A2(_13289_),
    .B1(_13282_),
    .Y(_06052_));
 sky130_fd_sc_hd__and2_0 _17106_ (.A(_06038_),
    .B(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__o21ai_1 _17107_ (.A1(_06021_),
    .A2(_06022_),
    .B1(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__o21ai_2 _17108_ (.A1(_13289_),
    .A2(_06047_),
    .B1(_13297_),
    .Y(_06055_));
 sky130_fd_sc_hd__a21oi_2 _17109_ (.A1(_06040_),
    .A2(_06052_),
    .B1(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__a21oi_1 _17110_ (.A1(_06054_),
    .A2(_06056_),
    .B1(_13296_),
    .Y(_06057_));
 sky130_fd_sc_hd__xnor2_2 _17111_ (.A(_13304_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__nor2_4 _17112_ (.A(net349),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__inv_6 _17113_ (.A(_06059_),
    .Y(\hash.CA1.S0.X[10] ));
 sky130_fd_sc_hd__a21oi_1 _17114_ (.A1(_06043_),
    .A2(_06044_),
    .B1(\hash.CA1.S0.X[9] ),
    .Y(_06060_));
 sky130_fd_sc_hd__xnor2_1 _17115_ (.A(_06059_),
    .B(_06060_),
    .Y(_00659_));
 sky130_fd_sc_hd__inv_1 _17116_ (.A(_13304_),
    .Y(_06061_));
 sky130_fd_sc_hd__a211oi_4 _17117_ (.A1(_06045_),
    .A2(_06046_),
    .B1(_06061_),
    .C1(net1098),
    .Y(_06062_));
 sky130_fd_sc_hd__a21o_1 _17118_ (.A1(_13304_),
    .A2(_13296_),
    .B1(_13303_),
    .X(_06063_));
 sky130_fd_sc_hd__nor2_2 _17119_ (.A(_06062_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__xnor2_2 _17120_ (.A(_13311_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_8 _17121_ (.A(_06002_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__inv_1 _17122_ (.A(_06066_),
    .Y(\hash.CA1.S0.X[11] ));
 sky130_fd_sc_hd__a2111oi_2 _17123_ (.A1(_06033_),
    .A2(_06043_),
    .B1(\hash.CA1.S0.X[9] ),
    .C1(_06058_),
    .D1(net349),
    .Y(_06067_));
 sky130_fd_sc_hd__xor2_1 _17124_ (.A(_06066_),
    .B(_06067_),
    .X(_00660_));
 sky130_fd_sc_hd__or2_0 _17125_ (.A(_13311_),
    .B(_13310_),
    .X(_06068_));
 sky130_fd_sc_hd__o31ai_1 _17126_ (.A1(_13304_),
    .A2(_13303_),
    .A3(_13310_),
    .B1(_06068_),
    .Y(_06069_));
 sky130_fd_sc_hd__or3_1 _17127_ (.A(_13296_),
    .B(_13303_),
    .C(_13310_),
    .X(_06070_));
 sky130_fd_sc_hd__a21oi_2 _17128_ (.A1(_06054_),
    .A2(_06056_),
    .B1(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__or2_4 _17129_ (.A(_06069_),
    .B(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__xor2_4 _17130_ (.A(_13318_),
    .B(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__nor2_4 _17131_ (.A(net349),
    .B(_06073_),
    .Y(\hash.CA1.S0.X[12] ));
 sky130_fd_sc_hd__a2111oi_0 _17132_ (.A1(_06043_),
    .A2(_06044_),
    .B1(\hash.CA1.S0.X[9] ),
    .C1(_06058_),
    .D1(net349),
    .Y(_06074_));
 sky130_fd_sc_hd__nor2_2 _17133_ (.A(_06066_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__xor2_1 _17134_ (.A(\hash.CA1.S0.X[12] ),
    .B(_06075_),
    .X(_00661_));
 sky130_fd_sc_hd__or3_4 _17135_ (.A(_13310_),
    .B(_13317_),
    .C(_06063_),
    .X(_06076_));
 sky130_fd_sc_hd__a21o_1 _17136_ (.A1(_13318_),
    .A2(_06068_),
    .B1(_13317_),
    .X(_06077_));
 sky130_fd_sc_hd__o21ai_4 _17137_ (.A1(_06076_),
    .A2(_06062_),
    .B1(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__xnor2_2 _17138_ (.A(_13325_),
    .B(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__nor2_2 _17139_ (.A(net349),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__inv_1 _17140_ (.A(_06080_),
    .Y(\hash.CA1.S0.X[13] ));
 sky130_fd_sc_hd__nor4_2 _17141_ (.A(net349),
    .B(_06066_),
    .C(_06067_),
    .D(_06073_),
    .Y(_06081_));
 sky130_fd_sc_hd__xnor2_1 _17142_ (.A(\hash.CA1.S0.X[13] ),
    .B(_06081_),
    .Y(_00662_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1201 ();
 sky130_fd_sc_hd__clkinv_1 _17144_ (.A(_13332_),
    .Y(_06083_));
 sky130_fd_sc_hd__nor3_1 _17145_ (.A(_06083_),
    .B(_13317_),
    .C(_13324_),
    .Y(_06084_));
 sky130_fd_sc_hd__o21ai_0 _17146_ (.A1(_13318_),
    .A2(_13317_),
    .B1(_13325_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand2b_1 _17147_ (.A_N(_13324_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__nand2_1 _17148_ (.A(_13332_),
    .B(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__nand2_1 _17149_ (.A(_13318_),
    .B(_13325_),
    .Y(_06088_));
 sky130_fd_sc_hd__a21oi_1 _17150_ (.A1(_13325_),
    .A2(_13317_),
    .B1(_13324_),
    .Y(_06089_));
 sky130_fd_sc_hd__o311ai_0 _17151_ (.A1(_06069_),
    .A2(_06071_),
    .A3(_06088_),
    .B1(_06089_),
    .C1(_06083_),
    .Y(_06090_));
 sky130_fd_sc_hd__a22oi_2 _17152_ (.A1(_06072_),
    .A2(_06084_),
    .B1(_06087_),
    .B2(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__nand2_8 _17153_ (.A(_06002_),
    .B(_06091_),
    .Y(\hash.CA1.S0.X[14] ));
 sky130_fd_sc_hd__nand2_1 _17154_ (.A(\hash.CA1.S0.X[12] ),
    .B(_06075_),
    .Y(_06092_));
 sky130_fd_sc_hd__nand2_1 _17155_ (.A(_06080_),
    .B(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__xnor2_1 _17156_ (.A(\hash.CA1.S0.X[14] ),
    .B(_06093_),
    .Y(_00663_));
 sky130_fd_sc_hd__a21oi_2 _17157_ (.A1(_13332_),
    .A2(_13324_),
    .B1(_13331_),
    .Y(_06094_));
 sky130_fd_sc_hd__nor2_1 _17158_ (.A(_13325_),
    .B(_13324_),
    .Y(_06095_));
 sky130_fd_sc_hd__nor2_1 _17159_ (.A(_06083_),
    .B(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__nor2_1 _17160_ (.A(_13331_),
    .B(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__a21oi_1 _17161_ (.A1(_06078_),
    .A2(_06094_),
    .B1(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__xnor2_2 _17162_ (.A(_13339_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__nand2_4 _17163_ (.A(_06002_),
    .B(_06099_),
    .Y(\hash.CA1.S0.X[15] ));
 sky130_fd_sc_hd__or3_1 _17164_ (.A(\hash.CA1.S0.X[13] ),
    .B(_06081_),
    .C(\hash.CA1.S0.X[14] ),
    .X(_06100_));
 sky130_fd_sc_hd__xnor2_1 _17165_ (.A(\hash.CA1.S0.X[15] ),
    .B(_06100_),
    .Y(_00664_));
 sky130_fd_sc_hd__or4_4 _17166_ (.A(_06083_),
    .B(_06069_),
    .C(_06071_),
    .D(_06088_),
    .X(_06101_));
 sky130_fd_sc_hd__a21o_4 _17167_ (.A1(_13325_),
    .A2(_13317_),
    .B1(_13324_),
    .X(_06102_));
 sky130_fd_sc_hd__nand2_1 _17168_ (.A(_13332_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__nor2_1 _17169_ (.A(_13331_),
    .B(_13338_),
    .Y(_06104_));
 sky130_fd_sc_hd__nor2_1 _17170_ (.A(_13339_),
    .B(_13338_),
    .Y(_06105_));
 sky130_fd_sc_hd__a31oi_2 _17171_ (.A1(_06101_),
    .A2(_06103_),
    .A3(_06104_),
    .B1(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__xor2_2 _17172_ (.A(_13346_),
    .B(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__nor2_4 _17173_ (.A(net349),
    .B(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__clkinv_1 _17174_ (.A(_06108_),
    .Y(\hash.CA1.S0.X[16] ));
 sky130_fd_sc_hd__nand4_1 _17175_ (.A(_06002_),
    .B(_06080_),
    .C(_06091_),
    .D(_06099_),
    .Y(_06109_));
 sky130_fd_sc_hd__a21oi_2 _17176_ (.A1(\hash.CA1.S0.X[12] ),
    .A2(_06075_),
    .B1(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__xnor2_1 _17177_ (.A(_06108_),
    .B(_06110_),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_1 _17178_ (.A(_13345_),
    .Y(_06111_));
 sky130_fd_sc_hd__o21ai_2 _17179_ (.A1(_13331_),
    .A2(_06096_),
    .B1(_13339_),
    .Y(_06112_));
 sky130_fd_sc_hd__a21oi_1 _17180_ (.A1(_06078_),
    .A2(_06094_),
    .B1(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__o21ai_2 _17181_ (.A1(_13338_),
    .A2(_06113_),
    .B1(_13346_),
    .Y(_06114_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1200 ();
 sky130_fd_sc_hd__a21boi_2 _17183_ (.A1(_06111_),
    .A2(_06114_),
    .B1_N(_13353_),
    .Y(_06116_));
 sky130_fd_sc_hd__nor3b_2 _17184_ (.A(_13353_),
    .B(_13345_),
    .C_N(_06114_),
    .Y(_06117_));
 sky130_fd_sc_hd__nor3_4 _17185_ (.A(net350),
    .B(_06116_),
    .C(_06117_),
    .Y(\hash.CA1.S0.X[17] ));
 sky130_fd_sc_hd__or3_4 _17186_ (.A(_06081_),
    .B(_06107_),
    .C(_06109_),
    .X(_06118_));
 sky130_fd_sc_hd__xor2_1 _17187_ (.A(\hash.CA1.S0.X[17] ),
    .B(_06118_),
    .X(_00666_));
 sky130_fd_sc_hd__a21o_1 _17188_ (.A1(_13345_),
    .A2(_13353_),
    .B1(_13352_),
    .X(_06119_));
 sky130_fd_sc_hd__a31oi_1 _17189_ (.A1(_13346_),
    .A2(_13353_),
    .A3(_06106_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__xnor2_2 _17190_ (.A(_13360_),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__nand2_4 _17191_ (.A(_06002_),
    .B(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__inv_4 _17192_ (.A(_06122_),
    .Y(\hash.CA1.S0.X[18] ));
 sky130_fd_sc_hd__nand2_2 _17193_ (.A(_06108_),
    .B(_06110_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _17194_ (.A(\hash.CA1.S0.X[17] ),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__xnor2_1 _17195_ (.A(\hash.CA1.S0.X[18] ),
    .B(_06124_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_2 _17196_ (.A(_13346_),
    .B(_13353_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand3_1 _17197_ (.A(_13339_),
    .B(_13346_),
    .C(_13353_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand3_1 _17198_ (.A(_13346_),
    .B(_13353_),
    .C(_13338_),
    .Y(_06127_));
 sky130_fd_sc_hd__o21ai_1 _17199_ (.A1(_06094_),
    .A2(_06126_),
    .B1(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__nor2_1 _17200_ (.A(_06119_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__o31ai_1 _17201_ (.A1(_06078_),
    .A2(_06112_),
    .A3(_06125_),
    .B1(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__a21oi_1 _17202_ (.A1(_13360_),
    .A2(_06130_),
    .B1(_13359_),
    .Y(_06131_));
 sky130_fd_sc_hd__xnor2_2 _17203_ (.A(_13367_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__nor2_4 _17204_ (.A(net349),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__clkinvlp_2 _17205_ (.A(_06133_),
    .Y(\hash.CA1.S0.X[19] ));
 sky130_fd_sc_hd__nand2_2 _17206_ (.A(\hash.CA1.S0.X[17] ),
    .B(_06118_),
    .Y(_06134_));
 sky130_fd_sc_hd__o21ai_4 _17207_ (.A1(_06134_),
    .A2(_06122_),
    .B1(_06133_),
    .Y(_06135_));
 sky130_fd_sc_hd__or3_4 _17208_ (.A(_06134_),
    .B(_06122_),
    .C(_06133_),
    .X(_06136_));
 sky130_fd_sc_hd__nand2_1 _17209_ (.A(_06135_),
    .B(_06136_),
    .Y(_00668_));
 sky130_fd_sc_hd__a21oi_2 _17210_ (.A1(_13332_),
    .A2(_06102_),
    .B1(_13331_),
    .Y(_06137_));
 sky130_fd_sc_hd__nand2_1 _17211_ (.A(_13360_),
    .B(_13367_),
    .Y(_06138_));
 sky130_fd_sc_hd__nor2_1 _17212_ (.A(_06125_),
    .B(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__nand2_2 _17213_ (.A(_13339_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__a21oi_4 _17214_ (.A1(_06101_),
    .A2(_06137_),
    .B1(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__a21oi_1 _17215_ (.A1(_13353_),
    .A2(_13345_),
    .B1(_13352_),
    .Y(_06142_));
 sky130_fd_sc_hd__a21boi_0 _17216_ (.A1(_06142_),
    .A2(_06127_),
    .B1_N(_13360_),
    .Y(_06143_));
 sky130_fd_sc_hd__o21ai_2 _17217_ (.A1(_13359_),
    .A2(_06143_),
    .B1(_13367_),
    .Y(_06144_));
 sky130_fd_sc_hd__nand2b_4 _17218_ (.A_N(_13366_),
    .B(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__or3_4 _17219_ (.A(_13374_),
    .B(_06141_),
    .C(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__o21ai_2 _17220_ (.A1(_06141_),
    .A2(_06145_),
    .B1(_13374_),
    .Y(_06147_));
 sky130_fd_sc_hd__and3_4 _17221_ (.A(_06002_),
    .B(_06146_),
    .C(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1199 ();
 sky130_fd_sc_hd__a31oi_2 _17223_ (.A1(\hash.CA1.S0.X[17] ),
    .A2(\hash.CA1.S0.X[18] ),
    .A3(_06123_),
    .B1(\hash.CA1.S0.X[19] ),
    .Y(_06149_));
 sky130_fd_sc_hd__xnor2_1 _17224_ (.A(_06148_),
    .B(_06149_),
    .Y(_00670_));
 sky130_fd_sc_hd__nor4_4 _17225_ (.A(_06119_),
    .B(_13366_),
    .C(_13359_),
    .D(_06128_),
    .Y(_06150_));
 sky130_fd_sc_hd__o31ai_4 _17226_ (.A1(_06125_),
    .A2(_06112_),
    .A3(_06078_),
    .B1(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__o21ai_0 _17227_ (.A1(_13360_),
    .A2(_13359_),
    .B1(_13367_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2b_2 _17228_ (.A_N(_13366_),
    .B(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__a31o_4 _17229_ (.A1(_06151_),
    .A2(_13374_),
    .A3(_06153_),
    .B1(_13373_),
    .X(_06154_));
 sky130_fd_sc_hd__xor2_2 _17230_ (.A(_13381_),
    .B(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__and2_4 _17231_ (.A(_06002_),
    .B(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1198 ();
 sky130_fd_sc_hd__nand2_1 _17233_ (.A(_06135_),
    .B(_06148_),
    .Y(_06157_));
 sky130_fd_sc_hd__xnor2_1 _17234_ (.A(_06156_),
    .B(_06157_),
    .Y(_00671_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1197 ();
 sky130_fd_sc_hd__or3_4 _17236_ (.A(_13373_),
    .B(_13380_),
    .C(_06145_),
    .X(_06159_));
 sky130_fd_sc_hd__nor3_1 _17237_ (.A(_13374_),
    .B(_13373_),
    .C(_13380_),
    .Y(_06160_));
 sky130_fd_sc_hd__nor2_1 _17238_ (.A(_13381_),
    .B(_13380_),
    .Y(_06161_));
 sky130_fd_sc_hd__nor2_1 _17239_ (.A(_06160_),
    .B(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__o21ai_4 _17240_ (.A1(_06159_),
    .A2(_06141_),
    .B1(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__xor2_4 _17241_ (.A(_06163_),
    .B(_13388_),
    .X(_06164_));
 sky130_fd_sc_hd__nor2_4 _17242_ (.A(net350),
    .B(_06164_),
    .Y(\hash.CA1.S0.X[22] ));
 sky130_fd_sc_hd__nand4_1 _17243_ (.A(_06002_),
    .B(_06146_),
    .C(_06147_),
    .D(_06155_),
    .Y(_06165_));
 sky130_fd_sc_hd__nor2_1 _17244_ (.A(_06149_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__xor2_1 _17245_ (.A(\hash.CA1.S0.X[22] ),
    .B(_06166_),
    .X(_00672_));
 sky130_fd_sc_hd__a21o_1 _17246_ (.A1(_13381_),
    .A2(_06154_),
    .B1(_13380_),
    .X(_06167_));
 sky130_fd_sc_hd__a211o_4 _17247_ (.A1(_13388_),
    .A2(_06167_),
    .B1(_13387_),
    .C1(_13395_),
    .X(_06168_));
 sky130_fd_sc_hd__a211o_4 _17248_ (.A1(_06154_),
    .A2(_13381_),
    .B1(_13387_),
    .C1(_13380_),
    .X(_06169_));
 sky130_fd_sc_hd__o21a_4 _17249_ (.A1(_13388_),
    .A2(_13387_),
    .B1(_13395_),
    .X(_06170_));
 sky130_fd_sc_hd__a21oi_2 _17250_ (.A1(_06169_),
    .A2(_06170_),
    .B1(net351),
    .Y(_06171_));
 sky130_fd_sc_hd__nand2_8 _17251_ (.A(_06168_),
    .B(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__inv_4 _17252_ (.A(_06172_),
    .Y(\hash.CA1.S0.X[23] ));
 sky130_fd_sc_hd__nor2_2 _17253_ (.A(_06164_),
    .B(_06165_),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_1 _17254_ (.A(_06135_),
    .B(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__xnor2_1 _17255_ (.A(\hash.CA1.S0.X[23] ),
    .B(_06174_),
    .Y(_00673_));
 sky130_fd_sc_hd__inv_1 _17256_ (.A(_13387_),
    .Y(_06175_));
 sky130_fd_sc_hd__o211ai_1 _17257_ (.A1(_06141_),
    .A2(_06159_),
    .B1(_06162_),
    .C1(_13388_),
    .Y(_06176_));
 sky130_fd_sc_hd__a21boi_2 _17258_ (.A1(_06176_),
    .A2(_06175_),
    .B1_N(_13395_),
    .Y(_06177_));
 sky130_fd_sc_hd__o21ai_1 _17259_ (.A1(_13394_),
    .A2(_06177_),
    .B1(_13402_),
    .Y(_06178_));
 sky130_fd_sc_hd__o311a_4 _17260_ (.A1(_13402_),
    .A2(_13394_),
    .A3(_06177_),
    .B1(_06178_),
    .C1(_06002_),
    .X(_06179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1196 ();
 sky130_fd_sc_hd__nor4_2 _17262_ (.A(_06149_),
    .B(_06164_),
    .C(_06165_),
    .D(_06172_),
    .Y(_06180_));
 sky130_fd_sc_hd__xor2_1 _17263_ (.A(_06179_),
    .B(_06180_),
    .X(_00674_));
 sky130_fd_sc_hd__clkinv_1 _17264_ (.A(_13409_),
    .Y(_06181_));
 sky130_fd_sc_hd__a2111o_2 _17265_ (.A1(_06169_),
    .A2(_06170_),
    .B1(_06181_),
    .C1(_13394_),
    .D1(_13401_),
    .X(_06182_));
 sky130_fd_sc_hd__inv_1 _17266_ (.A(_13402_),
    .Y(_06183_));
 sky130_fd_sc_hd__nor2_2 _17267_ (.A(_06183_),
    .B(_13409_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand3_2 _17268_ (.A(_06169_),
    .B(_06170_),
    .C(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__nor3_1 _17269_ (.A(_13402_),
    .B(_06181_),
    .C(_13401_),
    .Y(_06186_));
 sky130_fd_sc_hd__a221oi_2 _17270_ (.A1(_06181_),
    .A2(_13401_),
    .B1(_06184_),
    .B2(_13394_),
    .C1(_06186_),
    .Y(_06187_));
 sky130_fd_sc_hd__nand4_1 _17271_ (.A(_06002_),
    .B(_06182_),
    .C(_06185_),
    .D(_06187_),
    .Y(\hash.CA1.S0.X[25] ));
 sky130_fd_sc_hd__and4_4 _17272_ (.A(_06135_),
    .B(\hash.CA1.S0.X[23] ),
    .C(_06173_),
    .D(_06179_),
    .X(_06188_));
 sky130_fd_sc_hd__xnor2_1 _17273_ (.A(net1056),
    .B(_06188_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand3_1 _17274_ (.A(_13388_),
    .B(_13395_),
    .C(_13402_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _17275_ (.A(_13381_),
    .B(_13409_),
    .Y(_06190_));
 sky130_fd_sc_hd__nor2_2 _17276_ (.A(_06189_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__o211a_4 _17277_ (.A1(_06141_),
    .A2(_06145_),
    .B1(_06191_),
    .C1(_13374_),
    .X(_06192_));
 sky130_fd_sc_hd__a21oi_1 _17278_ (.A1(_13395_),
    .A2(_13387_),
    .B1(_13394_),
    .Y(_06193_));
 sky130_fd_sc_hd__a41oi_1 _17279_ (.A1(_13388_),
    .A2(_13395_),
    .A3(_13402_),
    .A4(_13380_),
    .B1(_13401_),
    .Y(_06194_));
 sky130_fd_sc_hd__o21ai_0 _17280_ (.A1(_06183_),
    .A2(_06193_),
    .B1(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__a21oi_1 _17281_ (.A1(_13409_),
    .A2(_06195_),
    .B1(_13408_),
    .Y(_06196_));
 sky130_fd_sc_hd__nand2_1 _17282_ (.A(_13373_),
    .B(_06191_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_2 _17283_ (.A(_06196_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__nor3_2 _17284_ (.A(_13416_),
    .B(_06192_),
    .C(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__o21a_4 _17285_ (.A1(_06192_),
    .A2(_06198_),
    .B1(_13416_),
    .X(_06200_));
 sky130_fd_sc_hd__nor3_4 _17286_ (.A(net351),
    .B(_06200_),
    .C(_06199_),
    .Y(_06201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1195 ();
 sky130_fd_sc_hd__a21oi_1 _17288_ (.A1(_06179_),
    .A2(_06180_),
    .B1(net1056),
    .Y(_06202_));
 sky130_fd_sc_hd__xnor2_1 _17289_ (.A(net1096),
    .B(_06202_),
    .Y(_00676_));
 sky130_fd_sc_hd__and3_1 _17290_ (.A(_13374_),
    .B(_13416_),
    .C(_06191_),
    .X(_06203_));
 sky130_fd_sc_hd__nand3_2 _17291_ (.A(_06203_),
    .B(_06153_),
    .C(_06151_),
    .Y(_06204_));
 sky130_fd_sc_hd__inv_1 _17292_ (.A(_13416_),
    .Y(_06205_));
 sky130_fd_sc_hd__nand3_1 _17293_ (.A(_13416_),
    .B(_13373_),
    .C(_06191_),
    .Y(_06206_));
 sky130_fd_sc_hd__o21ai_0 _17294_ (.A1(_06205_),
    .A2(_06196_),
    .B1(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__inv_1 _17295_ (.A(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__nand3b_1 _17296_ (.A_N(_13415_),
    .B(_06204_),
    .C(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__xor2_1 _17297_ (.A(_13423_),
    .B(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__or2_4 _17298_ (.A(net350),
    .B(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1194 ();
 sky130_fd_sc_hd__nand3_4 _17300_ (.A(_06182_),
    .B(_06185_),
    .C(_06187_),
    .Y(_06212_));
 sky130_fd_sc_hd__o21ai_0 _17301_ (.A1(_06212_),
    .A2(_06188_),
    .B1(net1095),
    .Y(_06213_));
 sky130_fd_sc_hd__xor2_1 _17302_ (.A(_06211_),
    .B(_06213_),
    .X(_00677_));
 sky130_fd_sc_hd__o21a_1 _17303_ (.A1(_13415_),
    .A2(_06200_),
    .B1(_13423_),
    .X(_06214_));
 sky130_fd_sc_hd__nor3_1 _17304_ (.A(_13430_),
    .B(_13422_),
    .C(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__or2_0 _17305_ (.A(_13423_),
    .B(_13422_),
    .X(_06216_));
 sky130_fd_sc_hd__o311a_4 _17306_ (.A1(_13415_),
    .A2(_13422_),
    .A3(_06200_),
    .B1(_06216_),
    .C1(_13430_),
    .X(_06217_));
 sky130_fd_sc_hd__or3_4 _17307_ (.A(net351),
    .B(_06215_),
    .C(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1193 ();
 sky130_fd_sc_hd__a21o_1 _17309_ (.A1(_06212_),
    .A2(net1095),
    .B1(_06211_),
    .X(_06220_));
 sky130_fd_sc_hd__a31o_4 _17310_ (.A1(_06179_),
    .A2(_06180_),
    .A3(net1094),
    .B1(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__xnor2_1 _17311_ (.A(_06218_),
    .B(_06221_),
    .Y(_00678_));
 sky130_fd_sc_hd__nor3_1 _17312_ (.A(_13415_),
    .B(_13422_),
    .C(_13429_),
    .Y(_06222_));
 sky130_fd_sc_hd__a21oi_1 _17313_ (.A1(_13430_),
    .A2(_06216_),
    .B1(_13429_),
    .Y(_06223_));
 sky130_fd_sc_hd__a31oi_4 _17314_ (.A1(_06204_),
    .A2(_06208_),
    .A3(_06222_),
    .B1(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__xor2_1 _17315_ (.A(_13437_),
    .B(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__nor2_4 _17316_ (.A(net350),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__inv_6 _17317_ (.A(_06226_),
    .Y(\hash.CA1.S0.X[29] ));
 sky130_fd_sc_hd__and3b_1 _17318_ (.A_N(_06172_),
    .B(_06173_),
    .C(net1094),
    .X(_06227_));
 sky130_fd_sc_hd__nand3_1 _17319_ (.A(_06135_),
    .B(_06179_),
    .C(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21oi_1 _17320_ (.A1(_06212_),
    .A2(net1094),
    .B1(_06211_),
    .Y(_06229_));
 sky130_fd_sc_hd__a21oi_1 _17321_ (.A1(_06228_),
    .A2(_06229_),
    .B1(_06218_),
    .Y(_06230_));
 sky130_fd_sc_hd__xnor2_1 _17322_ (.A(\hash.CA1.S0.X[29] ),
    .B(_06230_),
    .Y(_00679_));
 sky130_fd_sc_hd__o21a_1 _17323_ (.A1(_13429_),
    .A2(_06217_),
    .B1(_13437_),
    .X(_06231_));
 sky130_fd_sc_hd__o21ai_1 _17324_ (.A1(_13436_),
    .A2(_06231_),
    .B1(_13444_),
    .Y(_06232_));
 sky130_fd_sc_hd__or3_4 _17325_ (.A(_13444_),
    .B(_13436_),
    .C(_06231_),
    .X(_06233_));
 sky130_fd_sc_hd__a21o_4 _17326_ (.A1(_06232_),
    .A2(_06233_),
    .B1(net351),
    .X(_06234_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1192 ();
 sky130_fd_sc_hd__inv_1 _17328_ (.A(_06218_),
    .Y(\hash.CA1.S0.X[28] ));
 sky130_fd_sc_hd__a21o_1 _17329_ (.A1(\hash.CA1.S0.X[28] ),
    .A2(_06221_),
    .B1(\hash.CA1.S0.X[29] ),
    .X(_06235_));
 sky130_fd_sc_hd__xnor2_1 _17330_ (.A(_06234_),
    .B(_06235_),
    .Y(_00681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1191 ();
 sky130_fd_sc_hd__maj3_1 _17332_ (.A(\hash.CA2.b_dash[31] ),
    .B(\hash.CA2.a_dash[31] ),
    .C(_04612_),
    .X(_06237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1190 ();
 sky130_fd_sc_hd__mux2i_1 _17334_ (.A0(\hash.CA2.f_dash[31] ),
    .A1(\hash.CA2.e_dash[31] ),
    .S(\hash.CA2.S1.X[31] ),
    .Y(_06239_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1187 ();
 sky130_fd_sc_hd__xor2_1 _17338_ (.A(\hash.CA2.S1.X[5] ),
    .B(\hash.CA2.S1.X[24] ),
    .X(_06243_));
 sky130_fd_sc_hd__xnor2_1 _17339_ (.A(\hash.CA2.S1.X[10] ),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__xnor2_2 _17340_ (.A(_06239_),
    .B(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__o211ai_1 _17341_ (.A1(_04723_),
    .A2(_04749_),
    .B1(_04775_),
    .C1(_04751_),
    .Y(_06246_));
 sky130_fd_sc_hd__a31o_4 _17342_ (.A1(_13441_),
    .A2(_04776_),
    .A3(_06246_),
    .B1(_13440_),
    .X(_06247_));
 sky130_fd_sc_hd__xor2_4 _17343_ (.A(_06245_),
    .B(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__and3_4 _17344_ (.A(_04457_),
    .B(net1091),
    .C(_04590_),
    .X(_06249_));
 sky130_fd_sc_hd__a21boi_0 _17345_ (.A1(_04457_),
    .A2(net1091),
    .B1_N(_04592_),
    .Y(_06250_));
 sky130_fd_sc_hd__inv_1 _17346_ (.A(_04595_),
    .Y(_06251_));
 sky130_fd_sc_hd__xnor2_1 _17347_ (.A(\hash.CA2.p4[31] ),
    .B(_12360_),
    .Y(_06252_));
 sky130_fd_sc_hd__xnor2_1 _17348_ (.A(_12082_),
    .B(_12356_),
    .Y(_06253_));
 sky130_fd_sc_hd__xnor2_2 _17349_ (.A(_06252_),
    .B(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__xnor3_1 _17350_ (.A(_12948_),
    .B(_04472_),
    .C(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__or4_4 _17351_ (.A(_06249_),
    .B(_06250_),
    .C(_06251_),
    .D(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__o31ai_1 _17352_ (.A1(_06249_),
    .A2(_06250_),
    .A3(_06251_),
    .B1(_06255_),
    .Y(_06257_));
 sky130_fd_sc_hd__nand2_2 _17353_ (.A(_06256_),
    .B(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__nand2_1 _17354_ (.A(_13444_),
    .B(_13436_),
    .Y(_06259_));
 sky130_fd_sc_hd__inv_1 _17355_ (.A(_13443_),
    .Y(_06260_));
 sky130_fd_sc_hd__a22oi_1 _17356_ (.A1(_06256_),
    .A2(_06257_),
    .B1(_06259_),
    .B2(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__a41o_1 _17357_ (.A1(_13437_),
    .A2(_13444_),
    .A3(_06224_),
    .A4(_06258_),
    .B1(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__nor4_2 _17358_ (.A(_13436_),
    .B(_13443_),
    .C(_06224_),
    .D(_06258_),
    .Y(_06263_));
 sky130_fd_sc_hd__nor4_1 _17359_ (.A(_13437_),
    .B(_13436_),
    .C(_13443_),
    .D(_06258_),
    .Y(_06264_));
 sky130_fd_sc_hd__nor3_1 _17360_ (.A(_13444_),
    .B(_13443_),
    .C(_06258_),
    .Y(_06265_));
 sky130_fd_sc_hd__or4_4 _17361_ (.A(_06262_),
    .B(_06263_),
    .C(_06264_),
    .D(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__xor2_2 _17362_ (.A(_06248_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__xnor2_2 _17363_ (.A(_06237_),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_8 _17364_ (.A(_06002_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__inv_1 _17365_ (.A(_06269_),
    .Y(\hash.CA1.S0.X[31] ));
 sky130_fd_sc_hd__nor3_1 _17366_ (.A(\hash.CA1.S0.X[29] ),
    .B(_06230_),
    .C(_06234_),
    .Y(_06270_));
 sky130_fd_sc_hd__xor2_1 _17367_ (.A(_06269_),
    .B(_06270_),
    .X(_00682_));
 sky130_fd_sc_hd__xor2_1 _17368_ (.A(\hash.CA1.S0.X[3] ),
    .B(\hash.CA1.S0.X[14] ),
    .X(_06271_));
 sky130_fd_sc_hd__xnor2_1 _17369_ (.A(_06172_),
    .B(_06271_),
    .Y(_13548_));
 sky130_fd_sc_hd__inv_1 _17370_ (.A(_13548_),
    .Y(_12881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1184 ();
 sky130_fd_sc_hd__nor2b_4 _17374_ (.A(net349),
    .B_N(_12082_),
    .Y(\hash.CA1.b[1] ));
 sky130_fd_sc_hd__a21oi_1 _17375_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_13241_),
    .B1(_12082_),
    .Y(_06275_));
 sky130_fd_sc_hd__nor2_1 _17376_ (.A(\hash.CA2.a_dash[1] ),
    .B(_13241_),
    .Y(_06276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1183 ();
 sky130_fd_sc_hd__o21ai_1 _17378_ (.A1(_06275_),
    .A2(_06276_),
    .B1(_06002_),
    .Y(_13547_));
 sky130_fd_sc_hd__inv_1 _17379_ (.A(_13547_),
    .Y(_12880_));
 sky130_fd_sc_hd__nor2b_4 _17380_ (.A(net349),
    .B_N(\hash.CA2.a_dash[0] ),
    .Y(\hash.CA1.c[0] ));
 sky130_fd_sc_hd__nand2b_2 _17381_ (.A_N(_04421_),
    .B(_06002_),
    .Y(\hash.CA1.b[2] ));
 sky130_fd_sc_hd__nor2b_4 _17382_ (.A(net349),
    .B_N(\hash.CA2.a_dash[2] ),
    .Y(_13673_));
 sky130_fd_sc_hd__and2_0 _17383_ (.A(_06002_),
    .B(_04470_),
    .X(\hash.CA1.b[3] ));
 sky130_fd_sc_hd__nor2b_2 _17384_ (.A(net349),
    .B_N(\hash.CA2.a_dash[3] ),
    .Y(_13679_));
 sky130_fd_sc_hd__and2_4 _17385_ (.A(_06002_),
    .B(_04487_),
    .X(\hash.CA1.b[4] ));
 sky130_fd_sc_hd__and2_4 _17386_ (.A(_06002_),
    .B(_04501_),
    .X(\hash.CA1.b[5] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1182 ();
 sky130_fd_sc_hd__or2_4 _17388_ (.A(net350),
    .B(\hash.CA2.a_dash[5] ),
    .X(_13691_));
 sky130_fd_sc_hd__and2_4 _17389_ (.A(_06002_),
    .B(_04522_),
    .X(\hash.CA1.b[6] ));
 sky130_fd_sc_hd__or2_4 _17390_ (.A(net350),
    .B(\hash.CA2.a_dash[6] ),
    .X(_13697_));
 sky130_fd_sc_hd__nand2_2 _17391_ (.A(_06002_),
    .B(_04543_),
    .Y(\hash.CA1.b[7] ));
 sky130_fd_sc_hd__and2_4 _17392_ (.A(_06002_),
    .B(_04562_),
    .X(_06279_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1181 ();
 sky130_fd_sc_hd__or2_4 _17394_ (.A(net350),
    .B(_04580_),
    .X(_06280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1180 ();
 sky130_fd_sc_hd__or2_4 _17396_ (.A(net350),
    .B(\hash.CA2.a_dash[9] ),
    .X(_13716_));
 sky130_fd_sc_hd__or2_4 _17397_ (.A(net349),
    .B(_04599_),
    .X(\hash.CA1.b[10] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1179 ();
 sky130_fd_sc_hd__nor2_4 _17399_ (.A(net350),
    .B(_04614_),
    .Y(_06282_));
 sky130_fd_sc_hd__inv_1 _17400_ (.A(_06282_),
    .Y(\hash.CA1.b[11] ));
 sky130_fd_sc_hd__and2_4 _17401_ (.A(_06002_),
    .B(_04623_),
    .X(_06283_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1178 ();
 sky130_fd_sc_hd__or2_0 _17403_ (.A(net350),
    .B(_04437_),
    .X(\hash.CA1.b[13] ));
 sky130_fd_sc_hd__or2_4 _17404_ (.A(net350),
    .B(\hash.CA2.a_dash[13] ),
    .X(_13740_));
 sky130_fd_sc_hd__nor2_1 _17405_ (.A(net350),
    .B(_04475_),
    .Y(\hash.CA1.b[14] ));
 sky130_fd_sc_hd__or2_4 _17406_ (.A(net350),
    .B(\hash.CA2.a_dash[14] ),
    .X(_13746_));
 sky130_fd_sc_hd__or2_4 _17407_ (.A(net350),
    .B(_04484_),
    .X(\hash.CA1.b[15] ));
 sky130_fd_sc_hd__or2_4 _17408_ (.A(net350),
    .B(\hash.CA2.a_dash[15] ),
    .X(_13753_));
 sky130_fd_sc_hd__nand2b_4 _17409_ (.A_N(_04503_),
    .B(_06002_),
    .Y(\hash.CA1.b[16] ));
 sky130_fd_sc_hd__or2_4 _17410_ (.A(net351),
    .B(_04520_),
    .X(\hash.CA1.b[17] ));
 sky130_fd_sc_hd__or2_4 _17411_ (.A(net351),
    .B(_04541_),
    .X(\hash.CA1.b[18] ));
 sky130_fd_sc_hd__and2_4 _17412_ (.A(_06002_),
    .B(_04559_),
    .X(_06284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1177 ();
 sky130_fd_sc_hd__or2_4 _17414_ (.A(net351),
    .B(\hash.CA2.a_dash[19] ),
    .X(_13778_));
 sky130_fd_sc_hd__nor2_1 _17415_ (.A(net350),
    .B(_04681_),
    .Y(\hash.CA1.b[20] ));
 sky130_fd_sc_hd__nand4_1 _17416_ (.A(_06002_),
    .B(_04591_),
    .C(_04593_),
    .D(_04595_),
    .Y(\hash.CA1.b[21] ));
 sky130_fd_sc_hd__or2_4 _17417_ (.A(net351),
    .B(_04420_),
    .X(\hash.CA1.b[22] ));
 sky130_fd_sc_hd__and2_4 _17418_ (.A(_06002_),
    .B(_04467_),
    .X(_06285_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1176 ();
 sky130_fd_sc_hd__nand2_1 _17420_ (.A(_06002_),
    .B(_04481_),
    .Y(\hash.CA1.b[24] ));
 sky130_fd_sc_hd__nand2_4 _17421_ (.A(_06002_),
    .B(_04499_),
    .Y(\hash.CA1.b[25] ));
 sky130_fd_sc_hd__clkinv_1 _17422_ (.A(_04517_),
    .Y(_06286_));
 sky130_fd_sc_hd__nor2_2 _17423_ (.A(net351),
    .B(_06286_),
    .Y(\hash.CA1.b[26] ));
 sky130_fd_sc_hd__or2_4 _17424_ (.A(net352),
    .B(\hash.CA2.a_dash[26] ),
    .X(_06287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1175 ();
 sky130_fd_sc_hd__nor2_2 _17426_ (.A(net351),
    .B(_04537_),
    .Y(_06288_));
 sky130_fd_sc_hd__inv_1 _17427_ (.A(_06288_),
    .Y(\hash.CA1.b[27] ));
 sky130_fd_sc_hd__or2_0 _17428_ (.A(net352),
    .B(\hash.CA2.a_dash[27] ),
    .X(_13827_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1174 ();
 sky130_fd_sc_hd__nand2_1 _17430_ (.A(_06002_),
    .B(_04662_),
    .Y(\hash.CA1.b[28] ));
 sky130_fd_sc_hd__or2_4 _17431_ (.A(net352),
    .B(\hash.CA2.a_dash[28] ),
    .X(_13834_));
 sky130_fd_sc_hd__or2_4 _17432_ (.A(net352),
    .B(\hash.CA2.a_dash[29] ),
    .X(_13840_));
 sky130_fd_sc_hd__nor2_1 _17433_ (.A(net351),
    .B(_04588_),
    .Y(\hash.CA1.b[30] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1173 ();
 sky130_fd_sc_hd__o21ai_0 _17435_ (.A1(_04608_),
    .A2(_04611_),
    .B1(_06002_),
    .Y(\hash.CA1.b[31] ));
 sky130_fd_sc_hd__nor2_4 _17436_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[1] ),
    .Y(_12368_));
 sky130_fd_sc_hd__nor2b_4 _17437_ (.A(\hash.reset ),
    .B_N(\hash.CA2.e_dash[2] ),
    .Y(_12375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1172 ();
 sky130_fd_sc_hd__nor2_4 _17439_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[3] ),
    .Y(_12383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1171 ();
 sky130_fd_sc_hd__nor2b_4 _17441_ (.A(\hash.reset ),
    .B_N(\hash.CA2.e_dash[4] ),
    .Y(_12386_));
 sky130_fd_sc_hd__nor2_4 _17442_ (.A(net355),
    .B(\hash.CA2.e_dash[5] ),
    .Y(_12391_));
 sky130_fd_sc_hd__nor2b_4 _17443_ (.A(net355),
    .B_N(\hash.CA2.e_dash[6] ),
    .Y(_12394_));
 sky130_fd_sc_hd__nor2_4 _17444_ (.A(net355),
    .B(\hash.CA2.e_dash[7] ),
    .Y(_12399_));
 sky130_fd_sc_hd__nor2_4 _17445_ (.A(net355),
    .B(\hash.CA2.e_dash[8] ),
    .Y(_12404_));
 sky130_fd_sc_hd__nor2b_4 _17446_ (.A(net355),
    .B_N(\hash.CA2.e_dash[9] ),
    .Y(_12407_));
 sky130_fd_sc_hd__nor2b_4 _17447_ (.A(net355),
    .B_N(\hash.CA2.e_dash[10] ),
    .Y(_12410_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1170 ();
 sky130_fd_sc_hd__nor2_4 _17449_ (.A(net350),
    .B(\hash.CA2.e_dash[11] ),
    .Y(_12415_));
 sky130_fd_sc_hd__nor2_4 _17450_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[12] ),
    .Y(_12420_));
 sky130_fd_sc_hd__nor2b_4 _17451_ (.A(net354),
    .B_N(\hash.CA2.e_dash[13] ),
    .Y(_12423_));
 sky130_fd_sc_hd__nor2_4 _17452_ (.A(net350),
    .B(\hash.CA2.e_dash[14] ),
    .Y(_12428_));
 sky130_fd_sc_hd__nor2_4 _17453_ (.A(net350),
    .B(\hash.CA2.e_dash[15] ),
    .Y(_12433_));
 sky130_fd_sc_hd__nor2_4 _17454_ (.A(net350),
    .B(\hash.CA2.e_dash[16] ),
    .Y(_12438_));
 sky130_fd_sc_hd__nor2_4 _17455_ (.A(net350),
    .B(\hash.CA2.e_dash[17] ),
    .Y(_12443_));
 sky130_fd_sc_hd__nor2b_4 _17456_ (.A(net350),
    .B_N(\hash.CA2.e_dash[18] ),
    .Y(_12446_));
 sky130_fd_sc_hd__clkinv_2 _17457_ (.A(\hash.CA2.e_dash[19] ),
    .Y(_06294_));
 sky130_fd_sc_hd__nor2_4 _17458_ (.A(net350),
    .B(_06294_),
    .Y(_12449_));
 sky130_fd_sc_hd__nor2b_4 _17459_ (.A(net350),
    .B_N(\hash.CA2.e_dash[20] ),
    .Y(_12452_));
 sky130_fd_sc_hd__nor2b_4 _17460_ (.A(net350),
    .B_N(\hash.CA2.e_dash[21] ),
    .Y(_12455_));
 sky130_fd_sc_hd__nor2b_4 _17461_ (.A(net350),
    .B_N(\hash.CA2.e_dash[22] ),
    .Y(_12458_));
 sky130_fd_sc_hd__nor2_4 _17462_ (.A(net353),
    .B(\hash.CA2.e_dash[23] ),
    .Y(_12463_));
 sky130_fd_sc_hd__nor2_1 _17463_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[24] ),
    .Y(_12468_));
 sky130_fd_sc_hd__nor2_2 _17464_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[25] ),
    .Y(_12473_));
 sky130_fd_sc_hd__nor2_1 _17465_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[26] ),
    .Y(_12478_));
 sky130_fd_sc_hd__nor2_2 _17466_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[27] ),
    .Y(_12483_));
 sky130_fd_sc_hd__nor2_2 _17467_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[28] ),
    .Y(_12488_));
 sky130_fd_sc_hd__nor2b_4 _17468_ (.A(\hash.reset ),
    .B_N(\hash.CA2.e_dash[29] ),
    .Y(_12491_));
 sky130_fd_sc_hd__nor2b_1 _17469_ (.A(\hash.reset ),
    .B_N(\hash.CA2.e_dash[30] ),
    .Y(_12494_));
 sky130_fd_sc_hd__nor2b_4 _17470_ (.A(\hash.reset ),
    .B_N(\hash.CA2.f_dash[1] ),
    .Y(_12505_));
 sky130_fd_sc_hd__nand2_2 _17471_ (.A(_06002_),
    .B(\hash.CA2.f_dash[2] ),
    .Y(_12667_));
 sky130_fd_sc_hd__inv_2 _17472_ (.A(_12667_),
    .Y(_12510_));
 sky130_fd_sc_hd__xor2_2 _17473_ (.A(_13848_),
    .B(_12510_),
    .X(_00896_));
 sky130_fd_sc_hd__nor2_2 _17474_ (.A(net355),
    .B(\hash.CA2.f_dash[3] ),
    .Y(_12515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1169 ();
 sky130_fd_sc_hd__nand3_2 _17476_ (.A(\hash.CA2.f_dash[0] ),
    .B(\hash.CA2.f_dash[1] ),
    .C(\hash.CA2.f_dash[2] ),
    .Y(_06296_));
 sky130_fd_sc_hd__xnor2_2 _17477_ (.A(\hash.CA2.f_dash[3] ),
    .B(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__nor2_1 _17478_ (.A(net352),
    .B(_06297_),
    .Y(_00899_));
 sky130_fd_sc_hd__nor2_4 _17479_ (.A(\hash.reset ),
    .B(\hash.CA2.f_dash[4] ),
    .Y(_12520_));
 sky130_fd_sc_hd__a21oi_4 _17480_ (.A1(\hash.CA2.f_dash[2] ),
    .A2(_13848_),
    .B1(\hash.CA2.f_dash[3] ),
    .Y(_06298_));
 sky130_fd_sc_hd__xnor2_2 _17481_ (.A(\hash.CA2.f_dash[4] ),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2_1 _17482_ (.A(_06002_),
    .B(_06299_),
    .Y(_00900_));
 sky130_fd_sc_hd__nor2b_4 _17483_ (.A(net355),
    .B_N(\hash.CA2.f_dash[5] ),
    .Y(_12525_));
 sky130_fd_sc_hd__nand3b_1 _17484_ (.A_N(\hash.CA2.f_dash[3] ),
    .B(_06296_),
    .C(_12520_),
    .Y(_06300_));
 sky130_fd_sc_hd__xor2_2 _17485_ (.A(_12525_),
    .B(_06300_),
    .X(_00901_));
 sky130_fd_sc_hd__nand2_4 _17486_ (.A(_06002_),
    .B(\hash.CA2.f_dash[6] ),
    .Y(_12693_));
 sky130_fd_sc_hd__inv_1 _17487_ (.A(_12693_),
    .Y(_12530_));
 sky130_fd_sc_hd__a21boi_4 _17488_ (.A1(_12520_),
    .A2(_06298_),
    .B1_N(_12525_),
    .Y(_06301_));
 sky130_fd_sc_hd__mux2i_4 _17489_ (.A0(_12693_),
    .A1(\hash.CA2.f_dash[6] ),
    .S(_06301_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_8 _17490_ (.A(_06002_),
    .B(\hash.CA2.f_dash[7] ),
    .Y(_12702_));
 sky130_fd_sc_hd__inv_4 _17491_ (.A(_12702_),
    .Y(_12535_));
 sky130_fd_sc_hd__nand3_4 _17492_ (.A(\hash.CA2.f_dash[6] ),
    .B(_12525_),
    .C(_06300_),
    .Y(_06302_));
 sky130_fd_sc_hd__xnor2_2 _17493_ (.A(_12535_),
    .B(_06302_),
    .Y(_00903_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1168 ();
 sky130_fd_sc_hd__nor2_4 _17495_ (.A(net354),
    .B(\hash.CA2.f_dash[8] ),
    .Y(_12540_));
 sky130_fd_sc_hd__and3_4 _17496_ (.A(\hash.CA2.f_dash[6] ),
    .B(_06301_),
    .C(_12535_),
    .X(_06304_));
 sky130_fd_sc_hd__xor2_2 _17497_ (.A(_12540_),
    .B(_06304_),
    .X(_00904_));
 sky130_fd_sc_hd__nand2_4 _17498_ (.A(_06002_),
    .B(\hash.CA2.f_dash[9] ),
    .Y(_12715_));
 sky130_fd_sc_hd__inv_4 _17499_ (.A(_12715_),
    .Y(_12545_));
 sky130_fd_sc_hd__nor2_1 _17500_ (.A(_12702_),
    .B(_06302_),
    .Y(_06305_));
 sky130_fd_sc_hd__o21a_4 _17501_ (.A1(\hash.CA2.f_dash[8] ),
    .A2(_06305_),
    .B1(\hash.CA2.f_dash[9] ),
    .X(_06306_));
 sky130_fd_sc_hd__nor3_2 _17502_ (.A(\hash.CA2.f_dash[8] ),
    .B(\hash.CA2.f_dash[9] ),
    .C(_06305_),
    .Y(_06307_));
 sky130_fd_sc_hd__o21ai_1 _17503_ (.A1(_06306_),
    .A2(_06307_),
    .B1(_06002_),
    .Y(_00905_));
 sky130_fd_sc_hd__nor2_4 _17504_ (.A(net354),
    .B(\hash.CA2.f_dash[10] ),
    .Y(_12550_));
 sky130_fd_sc_hd__o21ai_4 _17505_ (.A1(\hash.CA2.f_dash[8] ),
    .A2(_06304_),
    .B1(_12545_),
    .Y(_06308_));
 sky130_fd_sc_hd__mux2_1 _17506_ (.A0(\hash.CA2.f_dash[10] ),
    .A1(_12550_),
    .S(_06308_),
    .X(_00876_));
 sky130_fd_sc_hd__or2_4 _17507_ (.A(net354),
    .B(\hash.CA2.f_dash[11] ),
    .X(_12733_));
 sky130_fd_sc_hd__inv_1 _17508_ (.A(_12733_),
    .Y(_12555_));
 sky130_fd_sc_hd__or3_1 _17509_ (.A(\hash.CA2.f_dash[10] ),
    .B(\hash.CA2.f_dash[11] ),
    .C(_06306_),
    .X(_06309_));
 sky130_fd_sc_hd__o21ai_0 _17510_ (.A1(\hash.CA2.f_dash[10] ),
    .A2(_06306_),
    .B1(\hash.CA2.f_dash[11] ),
    .Y(_06310_));
 sky130_fd_sc_hd__nand3_1 _17511_ (.A(_06002_),
    .B(_06309_),
    .C(_06310_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_8 _17512_ (.A(_06002_),
    .B(\hash.CA2.f_dash[12] ),
    .Y(_06311_));
 sky130_fd_sc_hd__clkinv_2 _17513_ (.A(_06311_),
    .Y(_12560_));
 sky130_fd_sc_hd__nor3_2 _17514_ (.A(net352),
    .B(\hash.CA2.f_dash[10] ),
    .C(\hash.CA2.f_dash[11] ),
    .Y(_06312_));
 sky130_fd_sc_hd__nand2_1 _17515_ (.A(_06308_),
    .B(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__xnor2_1 _17516_ (.A(_06311_),
    .B(_06313_),
    .Y(_00878_));
 sky130_fd_sc_hd__inv_4 _17517_ (.A(\hash.CA2.f_dash[13] ),
    .Y(_06314_));
 sky130_fd_sc_hd__nor2_4 _17518_ (.A(net354),
    .B(_06314_),
    .Y(_12565_));
 sky130_fd_sc_hd__nor3_1 _17519_ (.A(\hash.CA2.f_dash[10] ),
    .B(_12702_),
    .C(_06302_),
    .Y(_06315_));
 sky130_fd_sc_hd__o21ai_4 _17520_ (.A1(\hash.CA2.f_dash[8] ),
    .A2(_06315_),
    .B1(\hash.CA2.f_dash[9] ),
    .Y(_06316_));
 sky130_fd_sc_hd__a21oi_4 _17521_ (.A1(_06312_),
    .A2(_06316_),
    .B1(_06311_),
    .Y(_06317_));
 sky130_fd_sc_hd__mux2_1 _17522_ (.A0(_12565_),
    .A1(_06314_),
    .S(_06317_),
    .X(_00879_));
 sky130_fd_sc_hd__nor2_4 _17523_ (.A(net354),
    .B(\hash.CA2.f_dash[14] ),
    .Y(_12570_));
 sky130_fd_sc_hd__and3_4 _17524_ (.A(\hash.CA2.f_dash[12] ),
    .B(_06313_),
    .C(_12565_),
    .X(_06318_));
 sky130_fd_sc_hd__xor2_1 _17525_ (.A(_12570_),
    .B(_06318_),
    .X(_00880_));
 sky130_fd_sc_hd__nor2_4 _17526_ (.A(net353),
    .B(\hash.CA2.f_dash[15] ),
    .Y(_12575_));
 sky130_fd_sc_hd__a21oi_1 _17527_ (.A1(\hash.CA2.f_dash[13] ),
    .A2(_06317_),
    .B1(\hash.CA2.f_dash[14] ),
    .Y(_06319_));
 sky130_fd_sc_hd__xnor2_1 _17528_ (.A(\hash.CA2.f_dash[15] ),
    .B(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_06002_),
    .B(_06320_),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2b_4 _17530_ (.A(net354),
    .B_N(\hash.CA2.f_dash[16] ),
    .Y(_12580_));
 sky130_fd_sc_hd__nor3_4 _17531_ (.A(net354),
    .B(\hash.CA2.f_dash[14] ),
    .C(\hash.CA2.f_dash[15] ),
    .Y(_06321_));
 sky130_fd_sc_hd__nand2b_2 _17532_ (.A_N(_06318_),
    .B(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__xor2_1 _17533_ (.A(_12580_),
    .B(_06322_),
    .X(_00882_));
 sky130_fd_sc_hd__nor2b_4 _17534_ (.A(net354),
    .B_N(\hash.CA2.f_dash[17] ),
    .Y(_12585_));
 sky130_fd_sc_hd__a21boi_4 _17535_ (.A1(\hash.CA2.f_dash[13] ),
    .A2(_06317_),
    .B1_N(_06321_),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2b_1 _17536_ (.A_N(_06323_),
    .B(_12580_),
    .Y(_06324_));
 sky130_fd_sc_hd__xnor2_1 _17537_ (.A(_12585_),
    .B(_06324_),
    .Y(_00883_));
 sky130_fd_sc_hd__nor2b_4 _17538_ (.A(net354),
    .B_N(\hash.CA2.f_dash[18] ),
    .Y(_06325_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1167 ();
 sky130_fd_sc_hd__nand2_4 _17540_ (.A(\hash.CA2.f_dash[17] ),
    .B(_12580_),
    .Y(_06326_));
 sky130_fd_sc_hd__nor2b_4 _17541_ (.A(_06326_),
    .B_N(_06322_),
    .Y(_06327_));
 sky130_fd_sc_hd__xor2_1 _17542_ (.A(_06325_),
    .B(_06327_),
    .X(_00884_));
 sky130_fd_sc_hd__nor2b_4 _17543_ (.A(net354),
    .B_N(\hash.CA2.f_dash[19] ),
    .Y(_12595_));
 sky130_fd_sc_hd__nor2_1 _17544_ (.A(_06323_),
    .B(_06326_),
    .Y(_06328_));
 sky130_fd_sc_hd__nand2_1 _17545_ (.A(\hash.CA2.f_dash[18] ),
    .B(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__xnor2_1 _17546_ (.A(_12595_),
    .B(_06329_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_2 _17547_ (.A(_06002_),
    .B(\hash.CA2.f_dash[20] ),
    .Y(_12794_));
 sky130_fd_sc_hd__inv_2 _17548_ (.A(_12794_),
    .Y(_12600_));
 sky130_fd_sc_hd__nand3_1 _17549_ (.A(\hash.CA2.f_dash[19] ),
    .B(_06325_),
    .C(_06327_),
    .Y(_06330_));
 sky130_fd_sc_hd__xnor2_1 _17550_ (.A(_12600_),
    .B(_06330_),
    .Y(_00886_));
 sky130_fd_sc_hd__nor2_4 _17551_ (.A(net354),
    .B(\hash.CA2.f_dash[21] ),
    .Y(_12605_));
 sky130_fd_sc_hd__clkinvlp_2 _17552_ (.A(_12605_),
    .Y(_12803_));
 sky130_fd_sc_hd__nand3_1 _17553_ (.A(\hash.CA2.f_dash[19] ),
    .B(\hash.CA2.f_dash[20] ),
    .C(_06325_),
    .Y(_06331_));
 sky130_fd_sc_hd__or3_4 _17554_ (.A(_06323_),
    .B(_06326_),
    .C(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__xnor2_1 _17555_ (.A(_12605_),
    .B(_06332_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_4 _17556_ (.A(net353),
    .B(\hash.CA2.f_dash[22] ),
    .Y(_12610_));
 sky130_fd_sc_hd__nand2_1 _17557_ (.A(\hash.CA2.f_dash[19] ),
    .B(_06325_),
    .Y(_06333_));
 sky130_fd_sc_hd__nor3_1 _17558_ (.A(\hash.CA2.f_dash[21] ),
    .B(_12794_),
    .C(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__nor2_1 _17559_ (.A(_06321_),
    .B(_06331_),
    .Y(_06335_));
 sky130_fd_sc_hd__a31oi_1 _17560_ (.A1(_06318_),
    .A2(_06321_),
    .A3(_06334_),
    .B1(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__o21ai_0 _17561_ (.A1(_06326_),
    .A2(_06336_),
    .B1(_12605_),
    .Y(_06337_));
 sky130_fd_sc_hd__xor2_1 _17562_ (.A(_12610_),
    .B(_06337_),
    .X(_00888_));
 sky130_fd_sc_hd__nor2_2 _17563_ (.A(net353),
    .B(\hash.CA2.f_dash[23] ),
    .Y(_12615_));
 sky130_fd_sc_hd__clkinvlp_2 _17564_ (.A(_12615_),
    .Y(_12819_));
 sky130_fd_sc_hd__nor2_2 _17565_ (.A(\hash.CA2.f_dash[22] ),
    .B(_12803_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _17566_ (.A(_06332_),
    .B(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__xnor2_1 _17567_ (.A(_12819_),
    .B(_06339_),
    .Y(_00889_));
 sky130_fd_sc_hd__nor2_2 _17568_ (.A(net353),
    .B(\hash.CA2.f_dash[24] ),
    .Y(_12620_));
 sky130_fd_sc_hd__nand4_1 _17569_ (.A(\hash.CA2.f_dash[19] ),
    .B(\hash.CA2.f_dash[20] ),
    .C(_06325_),
    .D(_06327_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand3b_1 _17570_ (.A_N(\hash.CA2.f_dash[23] ),
    .B(_06338_),
    .C(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__xor2_1 _17571_ (.A(\hash.CA2.f_dash[24] ),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__nand2_1 _17572_ (.A(_06002_),
    .B(_06342_),
    .Y(_00890_));
 sky130_fd_sc_hd__nor2_4 _17573_ (.A(net353),
    .B(\hash.CA2.f_dash[25] ),
    .Y(_12625_));
 sky130_fd_sc_hd__inv_2 _17574_ (.A(_12625_),
    .Y(_12835_));
 sky130_fd_sc_hd__nor2_1 _17575_ (.A(\hash.CA2.f_dash[24] ),
    .B(_12819_),
    .Y(_06343_));
 sky130_fd_sc_hd__nand3_1 _17576_ (.A(_06332_),
    .B(_06338_),
    .C(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__xnor2_1 _17577_ (.A(_12835_),
    .B(_06344_),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2b_4 _17578_ (.A(net353),
    .B_N(\hash.CA2.f_dash[26] ),
    .Y(_12630_));
 sky130_fd_sc_hd__nand2_1 _17579_ (.A(_06327_),
    .B(_06334_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand4_1 _17580_ (.A(_06338_),
    .B(_12625_),
    .C(_06343_),
    .D(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__xor2_1 _17581_ (.A(_12630_),
    .B(_06346_),
    .X(_00892_));
 sky130_fd_sc_hd__nor2_2 _17582_ (.A(net353),
    .B(\hash.CA2.f_dash[27] ),
    .Y(_12635_));
 sky130_fd_sc_hd__inv_1 _17583_ (.A(_12635_),
    .Y(_12850_));
 sky130_fd_sc_hd__nand4_1 _17584_ (.A(_06332_),
    .B(_06338_),
    .C(_12625_),
    .D(_06343_),
    .Y(_06347_));
 sky130_fd_sc_hd__nand2_1 _17585_ (.A(_12630_),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__mux2_1 _17586_ (.A0(\hash.CA2.f_dash[27] ),
    .A1(_12635_),
    .S(_06348_),
    .X(_00893_));
 sky130_fd_sc_hd__or2_4 _17587_ (.A(net353),
    .B(\hash.CA2.f_dash[28] ),
    .X(_12858_));
 sky130_fd_sc_hd__inv_1 _17588_ (.A(_12858_),
    .Y(_12640_));
 sky130_fd_sc_hd__a21oi_1 _17589_ (.A1(\hash.CA2.f_dash[26] ),
    .A2(_06346_),
    .B1(\hash.CA2.f_dash[27] ),
    .Y(_06349_));
 sky130_fd_sc_hd__xnor2_1 _17590_ (.A(\hash.CA2.f_dash[28] ),
    .B(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__nand2_1 _17591_ (.A(_06002_),
    .B(_06350_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_2 _17592_ (.A(_06002_),
    .B(\hash.CA2.f_dash[29] ),
    .Y(_06351_));
 sky130_fd_sc_hd__inv_2 _17593_ (.A(_06351_),
    .Y(_12645_));
 sky130_fd_sc_hd__nor2_1 _17594_ (.A(\hash.CA2.f_dash[27] ),
    .B(_12858_),
    .Y(_06352_));
 sky130_fd_sc_hd__nand2_1 _17595_ (.A(_06348_),
    .B(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__xnor2_1 _17596_ (.A(_06351_),
    .B(_06353_),
    .Y(_00895_));
 sky130_fd_sc_hd__nor2_4 _17597_ (.A(net353),
    .B(\hash.CA2.f_dash[30] ),
    .Y(_12650_));
 sky130_fd_sc_hd__inv_1 _17598_ (.A(_12650_),
    .Y(_12872_));
 sky130_fd_sc_hd__and3_1 _17599_ (.A(\hash.CA2.f_dash[26] ),
    .B(\hash.CA2.f_dash[29] ),
    .C(_06352_),
    .X(_06354_));
 sky130_fd_sc_hd__nor2_1 _17600_ (.A(_06351_),
    .B(_06352_),
    .Y(_06355_));
 sky130_fd_sc_hd__a21oi_1 _17601_ (.A1(_06346_),
    .A2(_06354_),
    .B1(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__xnor2_1 _17602_ (.A(_12650_),
    .B(_06356_),
    .Y(_00897_));
 sky130_fd_sc_hd__a211oi_1 _17603_ (.A1(_06347_),
    .A2(_06354_),
    .B1(_06355_),
    .C1(\hash.CA2.f_dash[30] ),
    .Y(_06357_));
 sky130_fd_sc_hd__xor2_1 _17604_ (.A(\hash.CA2.f_dash[31] ),
    .B(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__nand2_1 _17605_ (.A(_06002_),
    .B(_06358_),
    .Y(_00898_));
 sky130_fd_sc_hd__xnor2_1 _17606_ (.A(_13849_),
    .B(_12375_),
    .Y(_00865_));
 sky130_fd_sc_hd__o21ai_1 _17607_ (.A1(\hash.CA2.e_dash[0] ),
    .A2(\hash.CA2.e_dash[1] ),
    .B1(\hash.CA2.e_dash[2] ),
    .Y(_06359_));
 sky130_fd_sc_hd__xnor2_1 _17608_ (.A(\hash.CA2.e_dash[3] ),
    .B(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__nor2_1 _17609_ (.A(net349),
    .B(_06360_),
    .Y(_00868_));
 sky130_fd_sc_hd__nor2b_2 _17610_ (.A(_13849_),
    .B_N(\hash.CA2.e_dash[2] ),
    .Y(_06361_));
 sky130_fd_sc_hd__o21a_4 _17611_ (.A1(\hash.CA2.e_dash[3] ),
    .A2(_06361_),
    .B1(\hash.CA2.e_dash[4] ),
    .X(_06362_));
 sky130_fd_sc_hd__nor3_2 _17612_ (.A(\hash.CA2.e_dash[3] ),
    .B(\hash.CA2.e_dash[4] ),
    .C(_06361_),
    .Y(_06363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1166 ();
 sky130_fd_sc_hd__o21ai_4 _17614_ (.A1(_06362_),
    .A2(_06363_),
    .B1(_06002_),
    .Y(_00869_));
 sky130_fd_sc_hd__o21a_1 _17615_ (.A1(\hash.CA2.e_dash[0] ),
    .A2(\hash.CA2.e_dash[1] ),
    .B1(_12375_),
    .X(_06365_));
 sky130_fd_sc_hd__o21a_4 _17616_ (.A1(\hash.CA2.e_dash[3] ),
    .A2(_06365_),
    .B1(\hash.CA2.e_dash[4] ),
    .X(_06366_));
 sky130_fd_sc_hd__xor2_2 _17617_ (.A(\hash.CA2.e_dash[5] ),
    .B(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nor2_1 _17618_ (.A(net352),
    .B(_06367_),
    .Y(_00870_));
 sky130_fd_sc_hd__nor3_2 _17619_ (.A(net355),
    .B(\hash.CA2.e_dash[5] ),
    .C(_06362_),
    .Y(_06368_));
 sky130_fd_sc_hd__xnor2_2 _17620_ (.A(_12394_),
    .B(_06368_),
    .Y(_00871_));
 sky130_fd_sc_hd__o21ai_2 _17621_ (.A1(\hash.CA2.e_dash[5] ),
    .A2(_06366_),
    .B1(\hash.CA2.e_dash[6] ),
    .Y(_06369_));
 sky130_fd_sc_hd__xnor2_2 _17622_ (.A(\hash.CA2.e_dash[7] ),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_1 _17623_ (.A(net352),
    .B(_06370_),
    .Y(_00872_));
 sky130_fd_sc_hd__o21ai_2 _17624_ (.A1(\hash.CA2.e_dash[5] ),
    .A2(_06362_),
    .B1(\hash.CA2.e_dash[6] ),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2b_1 _17625_ (.A_N(\hash.CA2.e_dash[7] ),
    .B(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__xor2_1 _17626_ (.A(\hash.CA2.e_dash[8] ),
    .B(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__nand2_1 _17627_ (.A(_06002_),
    .B(_06373_),
    .Y(_00873_));
 sky130_fd_sc_hd__nor3_2 _17628_ (.A(net355),
    .B(\hash.CA2.e_dash[7] ),
    .C(\hash.CA2.e_dash[8] ),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_2 _17629_ (.A(_06369_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__xor2_2 _17630_ (.A(_12407_),
    .B(_06375_),
    .X(_00874_));
 sky130_fd_sc_hd__o21ai_0 _17631_ (.A1(\hash.CA2.e_dash[8] ),
    .A2(_06372_),
    .B1(\hash.CA2.e_dash[9] ),
    .Y(_06376_));
 sky130_fd_sc_hd__xor2_1 _17632_ (.A(\hash.CA2.e_dash[10] ),
    .B(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__nor2_1 _17633_ (.A(net352),
    .B(_06377_),
    .Y(_00844_));
 sky130_fd_sc_hd__and2_4 _17634_ (.A(\hash.CA2.e_dash[9] ),
    .B(_06375_),
    .X(_06378_));
 sky130_fd_sc_hd__nand2_2 _17635_ (.A(\hash.CA2.e_dash[10] ),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__xnor2_2 _17636_ (.A(\hash.CA2.e_dash[11] ),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__nor2_1 _17637_ (.A(net349),
    .B(_06380_),
    .Y(_00845_));
 sky130_fd_sc_hd__nand2_1 _17638_ (.A(\hash.CA2.e_dash[10] ),
    .B(_12407_),
    .Y(_06381_));
 sky130_fd_sc_hd__a21oi_2 _17639_ (.A1(_06371_),
    .A2(_06374_),
    .B1(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__or3_4 _17640_ (.A(\hash.CA2.e_dash[11] ),
    .B(\hash.CA2.e_dash[12] ),
    .C(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__o21ai_2 _17641_ (.A1(\hash.CA2.e_dash[11] ),
    .A2(_06382_),
    .B1(\hash.CA2.e_dash[12] ),
    .Y(_06384_));
 sky130_fd_sc_hd__nand3_4 _17642_ (.A(_06002_),
    .B(_06383_),
    .C(_06384_),
    .Y(_00846_));
 sky130_fd_sc_hd__a211o_1 _17643_ (.A1(_12410_),
    .A2(_06378_),
    .B1(\hash.CA2.e_dash[11] ),
    .C1(\hash.CA2.e_dash[12] ),
    .X(_06385_));
 sky130_fd_sc_hd__or2_4 _17644_ (.A(\hash.CA2.e_dash[13] ),
    .B(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__nand2_2 _17645_ (.A(\hash.CA2.e_dash[13] ),
    .B(_06385_),
    .Y(_06387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1165 ();
 sky130_fd_sc_hd__a21o_4 _17647_ (.A1(_06386_),
    .A2(_06387_),
    .B1(net350),
    .X(_00847_));
 sky130_fd_sc_hd__o311a_4 _17648_ (.A1(\hash.CA2.e_dash[11] ),
    .A2(\hash.CA2.e_dash[12] ),
    .A3(_06382_),
    .B1(\hash.CA2.e_dash[13] ),
    .C1(_06002_),
    .X(_06389_));
 sky130_fd_sc_hd__xor2_2 _17649_ (.A(_12428_),
    .B(_06389_),
    .X(_00848_));
 sky130_fd_sc_hd__nand2_1 _17650_ (.A(_12428_),
    .B(_06387_),
    .Y(_06390_));
 sky130_fd_sc_hd__xor2_2 _17651_ (.A(_12433_),
    .B(_06390_),
    .X(_00849_));
 sky130_fd_sc_hd__nor4_1 _17652_ (.A(net350),
    .B(\hash.CA2.e_dash[14] ),
    .C(\hash.CA2.e_dash[15] ),
    .D(_06389_),
    .Y(_06391_));
 sky130_fd_sc_hd__xnor2_1 _17653_ (.A(_12438_),
    .B(_06391_),
    .Y(_00850_));
 sky130_fd_sc_hd__nor4_1 _17654_ (.A(net350),
    .B(\hash.CA2.e_dash[14] ),
    .C(\hash.CA2.e_dash[15] ),
    .D(\hash.CA2.e_dash[16] ),
    .Y(_06392_));
 sky130_fd_sc_hd__nand2_1 _17655_ (.A(_06387_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__xor2_1 _17656_ (.A(_12443_),
    .B(_06393_),
    .X(_00851_));
 sky130_fd_sc_hd__or3b_4 _17657_ (.A(\hash.CA2.e_dash[17] ),
    .B(_06389_),
    .C_N(_06392_),
    .X(_06394_));
 sky130_fd_sc_hd__xor2_2 _17658_ (.A(_12446_),
    .B(_06394_),
    .X(_00852_));
 sky130_fd_sc_hd__o31a_1 _17659_ (.A1(net350),
    .A2(\hash.CA2.e_dash[17] ),
    .A3(_06393_),
    .B1(_12446_),
    .X(_06395_));
 sky130_fd_sc_hd__mux2_1 _17660_ (.A0(_12449_),
    .A1(_06294_),
    .S(_06395_),
    .X(_00853_));
 sky130_fd_sc_hd__and3_4 _17661_ (.A(\hash.CA2.e_dash[19] ),
    .B(_12446_),
    .C(_06394_),
    .X(_06396_));
 sky130_fd_sc_hd__xor2_1 _17662_ (.A(_12452_),
    .B(_06396_),
    .X(_00855_));
 sky130_fd_sc_hd__and3_4 _17663_ (.A(\hash.CA2.e_dash[19] ),
    .B(\hash.CA2.e_dash[20] ),
    .C(_06395_),
    .X(_06397_));
 sky130_fd_sc_hd__xor2_1 _17664_ (.A(_12455_),
    .B(_06397_),
    .X(_00856_));
 sky130_fd_sc_hd__nand3_1 _17665_ (.A(\hash.CA2.e_dash[20] ),
    .B(\hash.CA2.e_dash[21] ),
    .C(_06396_),
    .Y(_06398_));
 sky130_fd_sc_hd__xor2_1 _17666_ (.A(\hash.CA2.e_dash[22] ),
    .B(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__nor2_1 _17667_ (.A(net349),
    .B(_06399_),
    .Y(_00857_));
 sky130_fd_sc_hd__and3_4 _17668_ (.A(\hash.CA2.e_dash[21] ),
    .B(\hash.CA2.e_dash[22] ),
    .C(_12452_),
    .X(_06400_));
 sky130_fd_sc_hd__and3_4 _17669_ (.A(_12449_),
    .B(_06395_),
    .C(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__xor2_1 _17670_ (.A(_12463_),
    .B(_06401_),
    .X(_00858_));
 sky130_fd_sc_hd__and3_4 _17671_ (.A(_12463_),
    .B(_06396_),
    .C(_06400_),
    .X(_06402_));
 sky130_fd_sc_hd__or3_1 _17672_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .C(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__o21ai_0 _17673_ (.A1(\hash.CA2.e_dash[23] ),
    .A2(_06402_),
    .B1(\hash.CA2.e_dash[24] ),
    .Y(_06404_));
 sky130_fd_sc_hd__nand3_1 _17674_ (.A(_06002_),
    .B(_06403_),
    .C(_06404_),
    .Y(_00859_));
 sky130_fd_sc_hd__nor3_1 _17675_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .C(_06401_),
    .Y(_06405_));
 sky130_fd_sc_hd__xnor2_1 _17676_ (.A(\hash.CA2.e_dash[25] ),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand2_2 _17677_ (.A(_06002_),
    .B(_06406_),
    .Y(_00860_));
 sky130_fd_sc_hd__nor4_1 _17678_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .C(\hash.CA2.e_dash[25] ),
    .D(_06402_),
    .Y(_06407_));
 sky130_fd_sc_hd__xnor2_1 _17679_ (.A(\hash.CA2.e_dash[26] ),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand2_1 _17680_ (.A(_06002_),
    .B(_06408_),
    .Y(_00861_));
 sky130_fd_sc_hd__nor2_2 _17681_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .Y(_06409_));
 sky130_fd_sc_hd__nor4b_1 _17682_ (.A(\hash.CA2.e_dash[25] ),
    .B(\hash.CA2.e_dash[26] ),
    .C(_06401_),
    .D_N(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__xnor2_1 _17683_ (.A(\hash.CA2.e_dash[27] ),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_1 _17684_ (.A(_06002_),
    .B(_06411_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand4_1 _17685_ (.A(_12473_),
    .B(_12478_),
    .C(_12483_),
    .D(_06409_),
    .Y(_06412_));
 sky130_fd_sc_hd__nor2_1 _17686_ (.A(_06402_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__xnor2_1 _17687_ (.A(_12488_),
    .B(_06413_),
    .Y(_00863_));
 sky130_fd_sc_hd__or2_4 _17688_ (.A(\hash.CA2.e_dash[28] ),
    .B(_06412_),
    .X(_06414_));
 sky130_fd_sc_hd__a41oi_2 _17689_ (.A1(_12455_),
    .A2(_12458_),
    .A3(_06397_),
    .A4(_06409_),
    .B1(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__xnor2_1 _17690_ (.A(_12491_),
    .B(_06415_),
    .Y(_00864_));
 sky130_fd_sc_hd__o21ai_0 _17691_ (.A1(_06402_),
    .A2(_06414_),
    .B1(\hash.CA2.e_dash[29] ),
    .Y(_06416_));
 sky130_fd_sc_hd__xor2_1 _17692_ (.A(\hash.CA2.e_dash[30] ),
    .B(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__nor2_1 _17693_ (.A(net350),
    .B(_06417_),
    .Y(_00866_));
 sky130_fd_sc_hd__nor2b_4 _17694_ (.A(net352),
    .B_N(\hash.CA2.e_dash[31] ),
    .Y(_06418_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(\hash.CA2.e_dash[30] ),
    .B(_12491_),
    .Y(_06419_));
 sky130_fd_sc_hd__nor2_2 _17696_ (.A(_06415_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__xor2_1 _17697_ (.A(_06418_),
    .B(_06420_),
    .X(_00867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1164 ();
 sky130_fd_sc_hd__nor2b_1 _17699_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[4] ),
    .Y(\hash.CA1.f[4] ));
 sky130_fd_sc_hd__xnor2_2 _17700_ (.A(_13852_),
    .B(\hash.CA1.f[4] ),
    .Y(_00835_));
 sky130_fd_sc_hd__nor2b_1 _17701_ (.A(net355),
    .B_N(\hash.CA2.S1.X[5] ),
    .Y(\hash.CA1.f[5] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1163 ();
 sky130_fd_sc_hd__o21ai_0 _17703_ (.A1(\hash.CA2.S1.X[2] ),
    .A2(\hash.CA2.S1.X[3] ),
    .B1(\hash.CA2.S1.X[4] ),
    .Y(_06423_));
 sky130_fd_sc_hd__xor2_1 _17704_ (.A(\hash.CA2.S1.X[5] ),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__nor2_1 _17705_ (.A(net352),
    .B(_06424_),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2b_4 _17706_ (.A(net351),
    .B_N(\hash.CA2.S1.X[6] ),
    .Y(\hash.CA1.f[6] ));
 sky130_fd_sc_hd__nor2b_4 _17707_ (.A(_13852_),
    .B_N(\hash.CA2.S1.X[5] ),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _17708_ (.A(\hash.CA2.S1.X[4] ),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__xor2_1 _17709_ (.A(\hash.CA2.S1.X[6] ),
    .B(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__nor2_1 _17710_ (.A(net352),
    .B(_06427_),
    .Y(_00837_));
 sky130_fd_sc_hd__inv_2 _17711_ (.A(\hash.CA2.S1.X[7] ),
    .Y(_06428_));
 sky130_fd_sc_hd__nand2_4 _17712_ (.A(_06002_),
    .B(_06428_),
    .Y(\hash.CA1.f[7] ));
 sky130_fd_sc_hd__o2111ai_4 _17713_ (.A1(\hash.CA2.S1.X[2] ),
    .A2(\hash.CA2.S1.X[3] ),
    .B1(\hash.CA2.S1.X[5] ),
    .C1(\hash.CA1.f[4] ),
    .D1(\hash.CA1.f[6] ),
    .Y(_06429_));
 sky130_fd_sc_hd__inv_2 _17714_ (.A(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__nand2_1 _17715_ (.A(net1061),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__o21ai_2 _17716_ (.A1(\hash.CA1.f[7] ),
    .A2(_06430_),
    .B1(_06431_),
    .Y(_00838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1162 ();
 sky130_fd_sc_hd__inv_6 _17718_ (.A(\hash.CA2.S1.X[8] ),
    .Y(_06433_));
 sky130_fd_sc_hd__nor2_4 _17719_ (.A(net352),
    .B(_06433_),
    .Y(\hash.CA1.f[8] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1161 ();
 sky130_fd_sc_hd__a31oi_4 _17721_ (.A1(\hash.CA2.S1.X[6] ),
    .A2(\hash.CA1.f[4] ),
    .A3(_06425_),
    .B1(\hash.CA2.S1.X[7] ),
    .Y(_06435_));
 sky130_fd_sc_hd__xnor2_1 _17722_ (.A(_06433_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _17723_ (.A(_06002_),
    .B(_06436_),
    .Y(_00839_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1160 ();
 sky130_fd_sc_hd__nor2b_4 _17725_ (.A(net352),
    .B_N(\hash.CA2.S1.X[9] ),
    .Y(_06438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1159 ();
 sky130_fd_sc_hd__o21ai_2 _17727_ (.A1(net1059),
    .A2(_06430_),
    .B1(\hash.CA1.f[8] ),
    .Y(_06439_));
 sky130_fd_sc_hd__xnor2_1 _17728_ (.A(_06438_),
    .B(_06439_),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2b_4 _17729_ (.A(net352),
    .B_N(\hash.CA2.S1.X[10] ),
    .Y(\hash.CA1.f[10] ));
 sky130_fd_sc_hd__nand2_2 _17730_ (.A(\hash.CA2.S1.X[8] ),
    .B(_06438_),
    .Y(_06440_));
 sky130_fd_sc_hd__nor2_1 _17731_ (.A(_06435_),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__xor2_1 _17732_ (.A(\hash.CA1.f[10] ),
    .B(_06441_),
    .X(_00841_));
 sky130_fd_sc_hd__nor2_2 _17733_ (.A(net352),
    .B(\hash.CA2.S1.X[11] ),
    .Y(_06442_));
 sky130_fd_sc_hd__inv_4 _17734_ (.A(_06442_),
    .Y(\hash.CA1.f[11] ));
 sky130_fd_sc_hd__nand2_2 _17735_ (.A(\hash.CA2.S1.X[10] ),
    .B(_06438_),
    .Y(_06443_));
 sky130_fd_sc_hd__nor2_1 _17736_ (.A(_06439_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__xnor2_1 _17737_ (.A(\hash.CA1.f[11] ),
    .B(_06444_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2b_4 _17738_ (.A(net352),
    .B_N(\hash.CA2.S1.X[12] ),
    .Y(\hash.CA1.f[12] ));
 sky130_fd_sc_hd__nand4_1 _17739_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[9] ),
    .C(\hash.CA2.S1.X[10] ),
    .D(_06442_),
    .Y(_06445_));
 sky130_fd_sc_hd__nor2_1 _17740_ (.A(_06435_),
    .B(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__o21ai_2 _17741_ (.A1(\hash.CA1.f[11] ),
    .A2(_06446_),
    .B1(\hash.CA1.f[12] ),
    .Y(_06447_));
 sky130_fd_sc_hd__o31a_1 _17742_ (.A1(\hash.CA2.S1.X[12] ),
    .A2(\hash.CA1.f[11] ),
    .A3(_06446_),
    .B1(_06447_),
    .X(_00814_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1158 ();
 sky130_fd_sc_hd__or2_0 _17744_ (.A(net354),
    .B(\hash.CA2.S1.X[13] ),
    .X(\hash.CA1.f[13] ));
 sky130_fd_sc_hd__nand2_1 _17745_ (.A(net1059),
    .B(\hash.CA1.f[8] ),
    .Y(_06449_));
 sky130_fd_sc_hd__o32ai_2 _17746_ (.A1(net1060),
    .A2(_06429_),
    .A3(_06445_),
    .B1(_06449_),
    .B2(_06443_),
    .Y(_06450_));
 sky130_fd_sc_hd__o21ai_4 _17747_ (.A1(\hash.CA2.S1.X[11] ),
    .A2(_06450_),
    .B1(\hash.CA1.f[12] ),
    .Y(_06451_));
 sky130_fd_sc_hd__xor2_1 _17748_ (.A(\hash.CA1.f[13] ),
    .B(_06451_),
    .X(_00815_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1157 ();
 sky130_fd_sc_hd__or2_0 _17750_ (.A(net354),
    .B(\hash.CA2.S1.X[14] ),
    .X(\hash.CA1.f[14] ));
 sky130_fd_sc_hd__inv_2 _17751_ (.A(\hash.CA2.S1.X[11] ),
    .Y(_06453_));
 sky130_fd_sc_hd__o21ai_0 _17752_ (.A1(_06435_),
    .A2(_06445_),
    .B1(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__a21oi_2 _17753_ (.A1(\hash.CA2.S1.X[12] ),
    .A2(_06454_),
    .B1(\hash.CA2.S1.X[13] ),
    .Y(_06455_));
 sky130_fd_sc_hd__xnor2_2 _17754_ (.A(\hash.CA2.S1.X[14] ),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand2_1 _17755_ (.A(_06002_),
    .B(_06456_),
    .Y(_00816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1156 ();
 sky130_fd_sc_hd__nand2_2 _17757_ (.A(_06002_),
    .B(\hash.CA2.S1.X[15] ),
    .Y(_06458_));
 sky130_fd_sc_hd__inv_1 _17758_ (.A(_06458_),
    .Y(\hash.CA1.f[15] ));
 sky130_fd_sc_hd__nor2_2 _17759_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA1.f[14] ),
    .Y(_06459_));
 sky130_fd_sc_hd__nand2_2 _17760_ (.A(_06451_),
    .B(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__xnor2_1 _17761_ (.A(_06458_),
    .B(_06460_),
    .Y(_00817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1155 ();
 sky130_fd_sc_hd__clkinv_2 _17763_ (.A(\hash.CA2.S1.X[16] ),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_2 _17764_ (.A(_06002_),
    .B(_06462_),
    .Y(\hash.CA1.f[16] ));
 sky130_fd_sc_hd__a21oi_2 _17765_ (.A1(_06447_),
    .A2(_06459_),
    .B1(_06458_),
    .Y(_06463_));
 sky130_fd_sc_hd__xnor2_1 _17766_ (.A(\hash.CA1.f[16] ),
    .B(_06463_),
    .Y(_00818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1154 ();
 sky130_fd_sc_hd__nor2b_4 _17768_ (.A(net353),
    .B_N(\hash.CA2.S1.X[17] ),
    .Y(\hash.CA1.f[17] ));
 sky130_fd_sc_hd__a21o_4 _17769_ (.A1(\hash.CA2.S1.X[15] ),
    .A2(_06460_),
    .B1(\hash.CA1.f[16] ),
    .X(_06465_));
 sky130_fd_sc_hd__xor2_1 _17770_ (.A(\hash.CA1.f[17] ),
    .B(_06465_),
    .X(_00819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1153 ();
 sky130_fd_sc_hd__or2_4 _17772_ (.A(net353),
    .B(\hash.CA2.S1.X[18] ),
    .X(_06467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1152 ();
 sky130_fd_sc_hd__o21a_4 _17774_ (.A1(\hash.CA2.S1.X[16] ),
    .A2(_06463_),
    .B1(\hash.CA1.f[17] ),
    .X(_06468_));
 sky130_fd_sc_hd__xnor2_1 _17775_ (.A(_06467_),
    .B(_06468_),
    .Y(_00820_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1151 ();
 sky130_fd_sc_hd__nor2b_4 _17777_ (.A(net353),
    .B_N(\hash.CA2.S1.X[19] ),
    .Y(\hash.CA1.f[19] ));
 sky130_fd_sc_hd__nand2_1 _17778_ (.A(\hash.CA1.f[15] ),
    .B(_06460_),
    .Y(_06470_));
 sky130_fd_sc_hd__nand2_2 _17779_ (.A(_06462_),
    .B(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__a21oi_4 _17780_ (.A1(\hash.CA2.S1.X[17] ),
    .A2(_06471_),
    .B1(_06467_),
    .Y(_06472_));
 sky130_fd_sc_hd__xnor2_1 _17781_ (.A(\hash.CA1.f[19] ),
    .B(_06472_),
    .Y(_00821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1150 ();
 sky130_fd_sc_hd__nor2b_1 _17783_ (.A(net351),
    .B_N(\hash.CA2.S1.X[20] ),
    .Y(\hash.CA1.f[20] ));
 sky130_fd_sc_hd__o21ai_0 _17784_ (.A1(\hash.CA2.S1.X[18] ),
    .A2(_06468_),
    .B1(\hash.CA2.S1.X[19] ),
    .Y(_06474_));
 sky130_fd_sc_hd__xor2_1 _17785_ (.A(\hash.CA2.S1.X[20] ),
    .B(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__nor2_1 _17786_ (.A(net354),
    .B(_06475_),
    .Y(_00822_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1149 ();
 sky130_fd_sc_hd__nor2b_4 _17788_ (.A(net353),
    .B_N(\hash.CA2.S1.X[21] ),
    .Y(\hash.CA1.f[21] ));
 sky130_fd_sc_hd__nand2_2 _17789_ (.A(\hash.CA2.S1.X[20] ),
    .B(\hash.CA1.f[19] ),
    .Y(_06477_));
 sky130_fd_sc_hd__a21oi_1 _17790_ (.A1(\hash.CA1.f[17] ),
    .A2(_06465_),
    .B1(\hash.CA2.S1.X[18] ),
    .Y(_06478_));
 sky130_fd_sc_hd__nor2_2 _17791_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__xor2_1 _17792_ (.A(\hash.CA1.f[21] ),
    .B(_06479_),
    .X(_00823_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1148 ();
 sky130_fd_sc_hd__nor2b_1 _17794_ (.A(net354),
    .B_N(\hash.CA2.S1.X[22] ),
    .Y(\hash.CA1.f[22] ));
 sky130_fd_sc_hd__o2111ai_1 _17795_ (.A1(\hash.CA2.S1.X[18] ),
    .A2(_06468_),
    .B1(\hash.CA1.f[19] ),
    .C1(\hash.CA2.S1.X[20] ),
    .D1(\hash.CA2.S1.X[21] ),
    .Y(_06481_));
 sky130_fd_sc_hd__xor2_1 _17796_ (.A(\hash.CA2.S1.X[22] ),
    .B(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__nor2_1 _17797_ (.A(net354),
    .B(_06482_),
    .Y(_00825_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1147 ();
 sky130_fd_sc_hd__clkinv_1 _17799_ (.A(\hash.CA2.S1.X[23] ),
    .Y(_06484_));
 sky130_fd_sc_hd__nor2_1 _17800_ (.A(net353),
    .B(_06484_),
    .Y(\hash.CA1.f[23] ));
 sky130_fd_sc_hd__nand2_2 _17801_ (.A(\hash.CA2.S1.X[22] ),
    .B(\hash.CA1.f[21] ),
    .Y(_06485_));
 sky130_fd_sc_hd__nor3_2 _17802_ (.A(_06472_),
    .B(_06477_),
    .C(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__xor2_1 _17803_ (.A(\hash.CA1.f[23] ),
    .B(_06486_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_4 _17804_ (.A(net353),
    .B(\hash.CA2.S1.X[24] ),
    .X(_06487_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1146 ();
 sky130_fd_sc_hd__nor4_1 _17806_ (.A(net353),
    .B(_06484_),
    .C(_06477_),
    .D(_06485_),
    .Y(_06488_));
 sky130_fd_sc_hd__o21ai_2 _17807_ (.A1(_06467_),
    .A2(_06468_),
    .B1(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__xor2_1 _17808_ (.A(_06487_),
    .B(_06489_),
    .X(_00827_));
 sky130_fd_sc_hd__clkinv_1 _17809_ (.A(net1071),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_1 _17810_ (.A(_06002_),
    .B(_06490_),
    .Y(\hash.CA1.f[25] ));
 sky130_fd_sc_hd__a21oi_1 _17811_ (.A1(\hash.CA2.S1.X[23] ),
    .A2(_06486_),
    .B1(\hash.CA2.S1.X[24] ),
    .Y(_06491_));
 sky130_fd_sc_hd__xnor2_1 _17812_ (.A(net1070),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__nand2_1 _17813_ (.A(_06002_),
    .B(_06492_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_4 _17814_ (.A(_06002_),
    .B(net1065),
    .Y(_06493_));
 sky130_fd_sc_hd__inv_1 _17815_ (.A(_06493_),
    .Y(\hash.CA1.f[26] ));
 sky130_fd_sc_hd__nor2_2 _17816_ (.A(\hash.CA2.S1.X[25] ),
    .B(_06487_),
    .Y(_06494_));
 sky130_fd_sc_hd__nand2_2 _17817_ (.A(_06489_),
    .B(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__xnor2_1 _17818_ (.A(_06493_),
    .B(_06495_),
    .Y(_00829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1145 ();
 sky130_fd_sc_hd__clkinvlp_4 _17820_ (.A(\hash.CA2.S1.X[27] ),
    .Y(_06497_));
 sky130_fd_sc_hd__nand2_1 _17821_ (.A(_06002_),
    .B(_06497_),
    .Y(\hash.CA1.f[27] ));
 sky130_fd_sc_hd__nand2_1 _17822_ (.A(\hash.CA2.S1.X[23] ),
    .B(_06486_),
    .Y(_06498_));
 sky130_fd_sc_hd__a21oi_1 _17823_ (.A1(_06498_),
    .A2(_06494_),
    .B1(_06493_),
    .Y(_06499_));
 sky130_fd_sc_hd__xnor2_1 _17824_ (.A(\hash.CA1.f[27] ),
    .B(_06499_),
    .Y(_00830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1144 ();
 sky130_fd_sc_hd__inv_2 _17826_ (.A(\hash.CA2.S1.X[28] ),
    .Y(_06501_));
 sky130_fd_sc_hd__nand2_1 _17827_ (.A(_06002_),
    .B(_06501_),
    .Y(\hash.CA1.f[28] ));
 sky130_fd_sc_hd__a21oi_1 _17828_ (.A1(net1066),
    .A2(_06495_),
    .B1(\hash.CA2.S1.X[27] ),
    .Y(_06502_));
 sky130_fd_sc_hd__xnor2_1 _17829_ (.A(\hash.CA2.S1.X[28] ),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(_06002_),
    .B(_06503_),
    .Y(_00831_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1143 ();
 sky130_fd_sc_hd__nand2_2 _17832_ (.A(_06002_),
    .B(\hash.CA2.S1.X[29] ),
    .Y(_06505_));
 sky130_fd_sc_hd__inv_1 _17833_ (.A(_06505_),
    .Y(\hash.CA1.f[29] ));
 sky130_fd_sc_hd__nor3_1 _17834_ (.A(_06485_),
    .B(_06487_),
    .C(_06493_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand3_1 _17835_ (.A(\hash.CA2.S1.X[23] ),
    .B(_06479_),
    .C(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__nor2_1 _17836_ (.A(\hash.CA2.S1.X[27] ),
    .B(\hash.CA1.f[28] ),
    .Y(_06508_));
 sky130_fd_sc_hd__o211ai_1 _17837_ (.A1(_06493_),
    .A2(_06494_),
    .B1(_06507_),
    .C1(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__xnor2_1 _17838_ (.A(_06505_),
    .B(_06509_),
    .Y(_00832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1142 ();
 sky130_fd_sc_hd__nor2b_4 _17840_ (.A(net353),
    .B_N(\hash.CA2.S1.X[30] ),
    .Y(\hash.CA1.f[30] ));
 sky130_fd_sc_hd__a21oi_1 _17841_ (.A1(_06501_),
    .A2(_06502_),
    .B1(_06505_),
    .Y(_06511_));
 sky130_fd_sc_hd__xor2_1 _17842_ (.A(\hash.CA1.f[30] ),
    .B(_06511_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_4 _17843_ (.A(net353),
    .B(\hash.CA2.S1.X[31] ),
    .X(\hash.CA1.f[31] ));
 sky130_fd_sc_hd__nand3_2 _17844_ (.A(\hash.CA2.S1.X[29] ),
    .B(_06509_),
    .C(\hash.CA1.f[30] ),
    .Y(_06512_));
 sky130_fd_sc_hd__xor2_1 _17845_ (.A(\hash.CA1.f[31] ),
    .B(_06512_),
    .X(_00834_));
 sky130_fd_sc_hd__xor2_4 _17846_ (.A(_12364_),
    .B(_13449_),
    .X(_06513_));
 sky130_fd_sc_hd__nor2_4 _17847_ (.A(net353),
    .B(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__inv_4 _17848_ (.A(_06514_),
    .Y(\hash.CA1.S1.X[2] ));
 sky130_fd_sc_hd__xnor2_1 _17849_ (.A(_13855_),
    .B(_06514_),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_4 _17850_ (.A(net353),
    .B(_12365_),
    .Y(_13854_));
 sky130_fd_sc_hd__inv_4 _17851_ (.A(_13854_),
    .Y(\hash.CA1.S1.X[1] ));
 sky130_fd_sc_hd__inv_6 _17852_ (.A(_00781_),
    .Y(\hash.CA1.S1.X[0] ));
 sky130_fd_sc_hd__a211oi_2 _17853_ (.A1(_12362_),
    .A2(_13447_),
    .B1(_13446_),
    .C1(_13448_),
    .Y(_06515_));
 sky130_fd_sc_hd__o21ai_2 _17854_ (.A1(_13449_),
    .A2(_13448_),
    .B1(_13451_),
    .Y(_06516_));
 sky130_fd_sc_hd__nor2_4 _17855_ (.A(_06515_),
    .B(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__a21o_1 _17856_ (.A1(_12362_),
    .A2(_13447_),
    .B1(_13446_),
    .X(_06518_));
 sky130_fd_sc_hd__a211oi_2 _17857_ (.A1(_13449_),
    .A2(_06518_),
    .B1(_13448_),
    .C1(_13451_),
    .Y(_06519_));
 sky130_fd_sc_hd__o21ai_4 _17858_ (.A1(_06517_),
    .A2(_06519_),
    .B1(_06002_),
    .Y(\hash.CA1.S1.X[3] ));
 sky130_fd_sc_hd__or3_4 _17859_ (.A(_12365_),
    .B(\hash.CA1.S1.X[0] ),
    .C(_06513_),
    .X(_06520_));
 sky130_fd_sc_hd__xnor2_1 _17860_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06520_),
    .Y(_00806_));
 sky130_fd_sc_hd__a21o_1 _17861_ (.A1(_12364_),
    .A2(_13449_),
    .B1(_13448_),
    .X(_06521_));
 sky130_fd_sc_hd__a21oi_2 _17862_ (.A1(_13451_),
    .A2(_06521_),
    .B1(_13450_),
    .Y(_06522_));
 sky130_fd_sc_hd__xnor2_4 _17863_ (.A(_13453_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__nor2_4 _17864_ (.A(net353),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__inv_1 _17865_ (.A(_06524_),
    .Y(\hash.CA1.S1.X[4] ));
 sky130_fd_sc_hd__nand2_1 _17866_ (.A(_13855_),
    .B(_06514_),
    .Y(_06525_));
 sky130_fd_sc_hd__nor2_1 _17867_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__xnor2_1 _17868_ (.A(_06524_),
    .B(_06526_),
    .Y(_00807_));
 sky130_fd_sc_hd__o21a_4 _17869_ (.A1(_13453_),
    .A2(_13452_),
    .B1(_13455_),
    .X(_06527_));
 sky130_fd_sc_hd__o31ai_4 _17870_ (.A1(_13450_),
    .A2(_13452_),
    .A3(_06517_),
    .B1(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__o21bai_1 _17871_ (.A1(_06515_),
    .A2(_06516_),
    .B1_N(_13450_),
    .Y(_06529_));
 sky130_fd_sc_hd__a211o_4 _17872_ (.A1(_13453_),
    .A2(_06529_),
    .B1(_13452_),
    .C1(_13455_),
    .X(_06530_));
 sky130_fd_sc_hd__a21oi_4 _17873_ (.A1(_06528_),
    .A2(_06530_),
    .B1(net355),
    .Y(_06531_));
 sky130_fd_sc_hd__inv_4 _17874_ (.A(_06531_),
    .Y(\hash.CA1.S1.X[5] ));
 sky130_fd_sc_hd__or3_4 _17875_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06520_),
    .C(_06523_),
    .X(_06532_));
 sky130_fd_sc_hd__xor2_2 _17876_ (.A(_06531_),
    .B(_06532_),
    .X(_00808_));
 sky130_fd_sc_hd__a211oi_1 _17877_ (.A1(_12364_),
    .A2(_13449_),
    .B1(_13448_),
    .C1(_13450_),
    .Y(_06533_));
 sky130_fd_sc_hd__o21ai_1 _17878_ (.A1(_13451_),
    .A2(_13450_),
    .B1(_13453_),
    .Y(_06534_));
 sky130_fd_sc_hd__o21bai_1 _17879_ (.A1(_06533_),
    .A2(_06534_),
    .B1_N(_13452_),
    .Y(_06535_));
 sky130_fd_sc_hd__a21oi_1 _17880_ (.A1(_13455_),
    .A2(_06535_),
    .B1(_13454_),
    .Y(_06536_));
 sky130_fd_sc_hd__xor2_2 _17881_ (.A(_13457_),
    .B(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__nand2_8 _17882_ (.A(_06002_),
    .B(_06537_),
    .Y(\hash.CA1.S1.X[6] ));
 sky130_fd_sc_hd__nor2_1 _17883_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06523_),
    .Y(_06538_));
 sky130_fd_sc_hd__nand4_1 _17884_ (.A(_13855_),
    .B(_06514_),
    .C(_06531_),
    .D(_06538_),
    .Y(_06539_));
 sky130_fd_sc_hd__xnor2_2 _17885_ (.A(\hash.CA1.S1.X[6] ),
    .B(_06539_),
    .Y(_00809_));
 sky130_fd_sc_hd__nor3_1 _17886_ (.A(_13450_),
    .B(_13452_),
    .C(_13454_),
    .Y(_06540_));
 sky130_fd_sc_hd__o21ai_1 _17887_ (.A1(_06515_),
    .A2(_06516_),
    .B1(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__o21a_1 _17888_ (.A1(_13454_),
    .A2(_06527_),
    .B1(_13457_),
    .X(_06542_));
 sky130_fd_sc_hd__a21oi_1 _17889_ (.A1(_06541_),
    .A2(_06542_),
    .B1(_13456_),
    .Y(_06543_));
 sky130_fd_sc_hd__xor2_1 _17890_ (.A(_13459_),
    .B(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__nor2_4 _17891_ (.A(net355),
    .B(_06544_),
    .Y(\hash.CA1.S1.X[7] ));
 sky130_fd_sc_hd__nor3_1 _17892_ (.A(\hash.CA1.S1.X[5] ),
    .B(_06532_),
    .C(\hash.CA1.S1.X[6] ),
    .Y(_06545_));
 sky130_fd_sc_hd__xnor2_1 _17893_ (.A(\hash.CA1.S1.X[7] ),
    .B(_06545_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor3_1 _17894_ (.A(_13452_),
    .B(_13454_),
    .C(_13456_),
    .Y(_06546_));
 sky130_fd_sc_hd__o21ai_1 _17895_ (.A1(_06533_),
    .A2(_06534_),
    .B1(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__o21a_1 _17896_ (.A1(_13455_),
    .A2(_13454_),
    .B1(_13457_),
    .X(_06548_));
 sky130_fd_sc_hd__o21a_1 _17897_ (.A1(_13456_),
    .A2(_06548_),
    .B1(_13459_),
    .X(_06549_));
 sky130_fd_sc_hd__a21oi_1 _17898_ (.A1(_06547_),
    .A2(_06549_),
    .B1(_13458_),
    .Y(_06550_));
 sky130_fd_sc_hd__xnor2_2 _17899_ (.A(net1105),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__and2_4 _17900_ (.A(_06002_),
    .B(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1141 ();
 sky130_fd_sc_hd__o21ai_0 _17902_ (.A1(\hash.CA1.S1.X[6] ),
    .A2(_06539_),
    .B1(\hash.CA1.S1.X[7] ),
    .Y(_06553_));
 sky130_fd_sc_hd__xnor2_1 _17903_ (.A(_06552_),
    .B(_06553_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand4_1 _17904_ (.A(_13459_),
    .B(net1105),
    .C(_06541_),
    .D(_06542_),
    .Y(_06554_));
 sky130_fd_sc_hd__a21o_1 _17905_ (.A1(_13459_),
    .A2(_13456_),
    .B1(_13458_),
    .X(_06555_));
 sky130_fd_sc_hd__a21oi_2 _17906_ (.A1(net1105),
    .A2(_06555_),
    .B1(_13460_),
    .Y(_06556_));
 sky130_fd_sc_hd__nand2_4 _17907_ (.A(_06554_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__xor2_1 _17908_ (.A(_13463_),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__nor2_4 _17909_ (.A(net355),
    .B(_06558_),
    .Y(_06559_));
 sky130_fd_sc_hd__clkinv_2 _17910_ (.A(_06559_),
    .Y(\hash.CA1.S1.X[9] ));
 sky130_fd_sc_hd__o311ai_2 _17911_ (.A1(\hash.CA1.S1.X[5] ),
    .A2(_06532_),
    .A3(\hash.CA1.S1.X[6] ),
    .B1(\hash.CA1.S1.X[7] ),
    .C1(_06551_),
    .Y(_06560_));
 sky130_fd_sc_hd__xnor2_1 _17912_ (.A(_06559_),
    .B(_06560_),
    .Y(_00812_));
 sky130_fd_sc_hd__o211ai_1 _17913_ (.A1(\hash.CA1.S1.X[6] ),
    .A2(_06539_),
    .B1(\hash.CA1.S1.X[7] ),
    .C1(_06551_),
    .Y(_06561_));
 sky130_fd_sc_hd__and4_4 _17914_ (.A(_13463_),
    .B(_13461_),
    .C(_06547_),
    .D(_06549_),
    .X(_06562_));
 sky130_fd_sc_hd__a21o_1 _17915_ (.A1(_13461_),
    .A2(_13458_),
    .B1(_13460_),
    .X(_06563_));
 sky130_fd_sc_hd__a21oi_2 _17916_ (.A1(_06563_),
    .A2(_13463_),
    .B1(_13462_),
    .Y(_06564_));
 sky130_fd_sc_hd__clkinv_2 _17917_ (.A(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__nor2_1 _17918_ (.A(_06562_),
    .B(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__xnor2_2 _17919_ (.A(_13465_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__nand2_8 _17920_ (.A(_06002_),
    .B(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__a21oi_2 _17921_ (.A1(_06559_),
    .A2(_06561_),
    .B1(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__and3_1 _17922_ (.A(_06559_),
    .B(_06568_),
    .C(_06561_),
    .X(_06570_));
 sky130_fd_sc_hd__nor2_1 _17923_ (.A(_06569_),
    .B(_06570_),
    .Y(_00782_));
 sky130_fd_sc_hd__nor2_1 _17924_ (.A(net355),
    .B(_13467_),
    .Y(_06571_));
 sky130_fd_sc_hd__nor2b_1 _17925_ (.A(net355),
    .B_N(_13467_),
    .Y(_06572_));
 sky130_fd_sc_hd__a21o_1 _17926_ (.A1(_13463_),
    .A2(_06557_),
    .B1(_13462_),
    .X(_06573_));
 sky130_fd_sc_hd__a21oi_2 _17927_ (.A1(_13465_),
    .A2(_06573_),
    .B1(_13464_),
    .Y(_06574_));
 sky130_fd_sc_hd__mux2_8 _17928_ (.A0(_06571_),
    .A1(_06572_),
    .S(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1140 ();
 sky130_fd_sc_hd__a21oi_2 _17930_ (.A1(_06559_),
    .A2(_06560_),
    .B1(_06568_),
    .Y(_06576_));
 sky130_fd_sc_hd__xor2_1 _17931_ (.A(_06575_),
    .B(_06576_),
    .X(_00783_));
 sky130_fd_sc_hd__a21o_4 _17932_ (.A1(_13467_),
    .A2(_13464_),
    .B1(_13466_),
    .X(_06577_));
 sky130_fd_sc_hd__o211a_1 _17933_ (.A1(_06562_),
    .A2(_06565_),
    .B1(_13465_),
    .C1(_13467_),
    .X(_06578_));
 sky130_fd_sc_hd__nor2_1 _17934_ (.A(_06577_),
    .B(_06578_),
    .Y(_06579_));
 sky130_fd_sc_hd__xnor2_1 _17935_ (.A(_13469_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__nor2_4 _17936_ (.A(net352),
    .B(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__clkinvlp_2 _17937_ (.A(_06581_),
    .Y(\hash.CA1.S1.X[12] ));
 sky130_fd_sc_hd__nand2_1 _17938_ (.A(_06569_),
    .B(_06575_),
    .Y(_06582_));
 sky130_fd_sc_hd__xnor2_1 _17939_ (.A(_06581_),
    .B(_06582_),
    .Y(_00784_));
 sky130_fd_sc_hd__nor2_1 _17940_ (.A(net355),
    .B(_13471_),
    .Y(_06583_));
 sky130_fd_sc_hd__nor2b_2 _17941_ (.A(net355),
    .B_N(_13471_),
    .Y(_06584_));
 sky130_fd_sc_hd__a21oi_1 _17942_ (.A1(_13463_),
    .A2(_06557_),
    .B1(_13462_),
    .Y(_06585_));
 sky130_fd_sc_hd__nand3_2 _17943_ (.A(_13469_),
    .B(_13465_),
    .C(_13467_),
    .Y(_06586_));
 sky130_fd_sc_hd__a21oi_4 _17944_ (.A1(_13469_),
    .A2(_06577_),
    .B1(_13468_),
    .Y(_06587_));
 sky130_fd_sc_hd__o21a_4 _17945_ (.A1(_06585_),
    .A2(_06586_),
    .B1(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__mux2i_4 _17946_ (.A0(_06583_),
    .A1(_06584_),
    .S(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__inv_6 _17947_ (.A(_06589_),
    .Y(\hash.CA1.S1.X[13] ));
 sky130_fd_sc_hd__nand2_1 _17948_ (.A(_06575_),
    .B(_06576_),
    .Y(_06590_));
 sky130_fd_sc_hd__nand2_1 _17949_ (.A(_06581_),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__xnor2_1 _17950_ (.A(_06589_),
    .B(_06591_),
    .Y(_00785_));
 sky130_fd_sc_hd__o211a_2 _17951_ (.A1(_06577_),
    .A2(_06578_),
    .B1(_13469_),
    .C1(_13471_),
    .X(_06592_));
 sky130_fd_sc_hd__a21oi_1 _17952_ (.A1(_13471_),
    .A2(_13468_),
    .B1(_13470_),
    .Y(_06593_));
 sky130_fd_sc_hd__inv_1 _17953_ (.A(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__o21ai_2 _17954_ (.A1(_06592_),
    .A2(_06594_),
    .B1(_13473_),
    .Y(_06595_));
 sky130_fd_sc_hd__or3_4 _17955_ (.A(_13473_),
    .B(_06592_),
    .C(_06594_),
    .X(_06596_));
 sky130_fd_sc_hd__a21oi_4 _17956_ (.A1(_06595_),
    .A2(_06596_),
    .B1(net355),
    .Y(_06597_));
 sky130_fd_sc_hd__clkinvlp_2 _17957_ (.A(_06597_),
    .Y(\hash.CA1.S1.X[14] ));
 sky130_fd_sc_hd__a21boi_4 _17958_ (.A1(_06569_),
    .A2(_06575_),
    .B1_N(_06581_),
    .Y(_06598_));
 sky130_fd_sc_hd__nand2_1 _17959_ (.A(\hash.CA1.S1.X[13] ),
    .B(\hash.CA1.S1.X[14] ),
    .Y(_06599_));
 sky130_fd_sc_hd__o21ai_4 _17960_ (.A1(_06598_),
    .A2(_06589_),
    .B1(_06597_),
    .Y(_06600_));
 sky130_fd_sc_hd__o21ai_2 _17961_ (.A1(_06598_),
    .A2(_06599_),
    .B1(_06600_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand2_2 _17962_ (.A(_13473_),
    .B(_13471_),
    .Y(_06601_));
 sky130_fd_sc_hd__a21oi_4 _17963_ (.A1(_13473_),
    .A2(_13470_),
    .B1(_13472_),
    .Y(_06602_));
 sky130_fd_sc_hd__o21ai_2 _17964_ (.A1(_06587_),
    .A2(_06601_),
    .B1(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__o21a_1 _17965_ (.A1(_06587_),
    .A2(_06601_),
    .B1(_06602_),
    .X(_06604_));
 sky130_fd_sc_hd__nor2_1 _17966_ (.A(_06586_),
    .B(_06601_),
    .Y(_06605_));
 sky130_fd_sc_hd__o21ai_0 _17967_ (.A1(_13463_),
    .A2(_13462_),
    .B1(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__nand2_1 _17968_ (.A(_06604_),
    .B(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__o31a_1 _17969_ (.A1(_13462_),
    .A2(_06557_),
    .A3(_06603_),
    .B1(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__xnor2_1 _17970_ (.A(_13475_),
    .B(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__nor2_4 _17971_ (.A(net351),
    .B(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1139 ();
 sky130_fd_sc_hd__o21a_4 _17973_ (.A1(_06581_),
    .A2(_06589_),
    .B1(_06597_),
    .X(_06611_));
 sky130_fd_sc_hd__nand3_2 _17974_ (.A(_06575_),
    .B(_06576_),
    .C(\hash.CA1.S1.X[13] ),
    .Y(_06612_));
 sky130_fd_sc_hd__nand2_1 _17975_ (.A(_06611_),
    .B(_06612_),
    .Y(_06613_));
 sky130_fd_sc_hd__xor2_1 _17976_ (.A(_06610_),
    .B(_06613_),
    .X(_00787_));
 sky130_fd_sc_hd__nor2_1 _17977_ (.A(_13474_),
    .B(_06605_),
    .Y(_06614_));
 sky130_fd_sc_hd__nor2_1 _17978_ (.A(_13475_),
    .B(_13474_),
    .Y(_06615_));
 sky130_fd_sc_hd__a21oi_2 _17979_ (.A1(_06604_),
    .A2(_06614_),
    .B1(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__or4_4 _17980_ (.A(_13474_),
    .B(_06562_),
    .C(_06565_),
    .D(_06603_),
    .X(_06617_));
 sky130_fd_sc_hd__and2_4 _17981_ (.A(_06616_),
    .B(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__xnor2_1 _17982_ (.A(_13477_),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__nor2_4 _17983_ (.A(net351),
    .B(_06619_),
    .Y(\hash.CA1.S1.X[16] ));
 sky130_fd_sc_hd__nand2_1 _17984_ (.A(_06600_),
    .B(_06610_),
    .Y(_06620_));
 sky130_fd_sc_hd__xnor2_1 _17985_ (.A(\hash.CA1.S1.X[16] ),
    .B(_06620_),
    .Y(_00788_));
 sky130_fd_sc_hd__a21o_1 _17986_ (.A1(_13477_),
    .A2(_13474_),
    .B1(_13476_),
    .X(_06621_));
 sky130_fd_sc_hd__a31oi_1 _17987_ (.A1(_13475_),
    .A2(_13481_),
    .A3(_06608_),
    .B1(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__xnor2_2 _17988_ (.A(_13479_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__nor2_4 _17989_ (.A(net354),
    .B(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__inv_1 _17990_ (.A(_06624_),
    .Y(\hash.CA1.S1.X[17] ));
 sky130_fd_sc_hd__nand2_1 _17991_ (.A(_06610_),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_06625_));
 sky130_fd_sc_hd__a21o_4 _17992_ (.A1(_06611_),
    .A2(_06612_),
    .B1(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__xnor2_1 _17993_ (.A(_06624_),
    .B(_06626_),
    .Y(_00789_));
 sky130_fd_sc_hd__a211oi_4 _17994_ (.A1(_06616_),
    .A2(_06617_),
    .B1(_13476_),
    .C1(_13478_),
    .Y(_06627_));
 sky130_fd_sc_hd__o21a_1 _17995_ (.A1(_13481_),
    .A2(_13476_),
    .B1(_13479_),
    .X(_06628_));
 sky130_fd_sc_hd__o21ai_1 _17996_ (.A1(_13478_),
    .A2(_06628_),
    .B1(_13483_),
    .Y(_06629_));
 sky130_fd_sc_hd__or2_4 _17997_ (.A(_06627_),
    .B(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__o21ai_0 _17998_ (.A1(_13476_),
    .A2(_06618_),
    .B1(_06628_),
    .Y(_06631_));
 sky130_fd_sc_hd__nor2_1 _17999_ (.A(_13483_),
    .B(_13478_),
    .Y(_06632_));
 sky130_fd_sc_hd__nand2_2 _18000_ (.A(_06631_),
    .B(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__a21oi_4 _18001_ (.A1(_06630_),
    .A2(_06633_),
    .B1(net351),
    .Y(_06634_));
 sky130_fd_sc_hd__inv_1 _18002_ (.A(_06634_),
    .Y(\hash.CA1.S1.X[18] ));
 sky130_fd_sc_hd__a31oi_2 _18003_ (.A1(_06600_),
    .A2(_06610_),
    .A3(\hash.CA1.S1.X[16] ),
    .B1(\hash.CA1.S1.X[17] ),
    .Y(_06635_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_06634_),
    .B(_06635_),
    .Y(_00790_));
 sky130_fd_sc_hd__a21o_1 _18005_ (.A1(_13479_),
    .A2(_06621_),
    .B1(_13478_),
    .X(_06636_));
 sky130_fd_sc_hd__a21oi_2 _18006_ (.A1(_06636_),
    .A2(_13483_),
    .B1(_13482_),
    .Y(_06637_));
 sky130_fd_sc_hd__and4_4 _18007_ (.A(_13475_),
    .B(_13479_),
    .C(_13481_),
    .D(_13483_),
    .X(_06638_));
 sky130_fd_sc_hd__o311ai_2 _18008_ (.A1(_13462_),
    .A2(_06557_),
    .A3(_06603_),
    .B1(_06607_),
    .C1(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__and2_4 _18009_ (.A(_06637_),
    .B(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__xnor2_1 _18010_ (.A(_13485_),
    .B(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nor2_4 _18011_ (.A(net351),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__inv_1 _18012_ (.A(_06642_),
    .Y(\hash.CA1.S1.X[19] ));
 sky130_fd_sc_hd__nand3_1 _18013_ (.A(_06624_),
    .B(_06626_),
    .C(_06634_),
    .Y(_06643_));
 sky130_fd_sc_hd__xnor2_1 _18014_ (.A(\hash.CA1.S1.X[19] ),
    .B(_06643_),
    .Y(_00791_));
 sky130_fd_sc_hd__nor2_1 _18015_ (.A(_13482_),
    .B(_13484_),
    .Y(_06644_));
 sky130_fd_sc_hd__or2_0 _18016_ (.A(_13485_),
    .B(_13484_),
    .X(_06645_));
 sky130_fd_sc_hd__a21boi_0 _18017_ (.A1(_06630_),
    .A2(_06644_),
    .B1_N(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__xnor2_1 _18018_ (.A(_13487_),
    .B(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__nor2_4 _18019_ (.A(net351),
    .B(_06647_),
    .Y(\hash.CA1.S1.X[20] ));
 sky130_fd_sc_hd__nand3_4 _18020_ (.A(_06624_),
    .B(_06634_),
    .C(_06642_),
    .Y(_06648_));
 sky130_fd_sc_hd__a31oi_4 _18021_ (.A1(_06600_),
    .A2(_06610_),
    .A3(\hash.CA1.S1.X[16] ),
    .B1(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__xnor2_1 _18022_ (.A(\hash.CA1.S1.X[20] ),
    .B(_06649_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_2 _18023_ (.A(_13485_),
    .B(_13491_),
    .Y(_06650_));
 sky130_fd_sc_hd__a21oi_1 _18024_ (.A1(_13487_),
    .A2(_13484_),
    .B1(_13486_),
    .Y(_06651_));
 sky130_fd_sc_hd__o21ai_2 _18025_ (.A1(_06640_),
    .A2(_06650_),
    .B1(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__xnor2_1 _18026_ (.A(_13489_),
    .B(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__nor2_4 _18027_ (.A(net351),
    .B(_06653_),
    .Y(\hash.CA1.S1.X[21] ));
 sky130_fd_sc_hd__nor2b_4 _18028_ (.A(_06648_),
    .B_N(_06626_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2b_2 _18029_ (.A_N(_06654_),
    .B(\hash.CA1.S1.X[20] ),
    .Y(_06655_));
 sky130_fd_sc_hd__xnor2_1 _18030_ (.A(\hash.CA1.S1.X[21] ),
    .B(_06655_),
    .Y(_00794_));
 sky130_fd_sc_hd__a21o_1 _18031_ (.A1(_13489_),
    .A2(_13486_),
    .B1(_13488_),
    .X(_06656_));
 sky130_fd_sc_hd__nor3_2 _18032_ (.A(_13482_),
    .B(_13484_),
    .C(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__a31oi_4 _18033_ (.A1(_13491_),
    .A2(_13495_),
    .A3(_06645_),
    .B1(_06656_),
    .Y(_06658_));
 sky130_fd_sc_hd__a21oi_1 _18034_ (.A1(_06630_),
    .A2(_06657_),
    .B1(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__xnor2_1 _18035_ (.A(_13493_),
    .B(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__nor2_4 _18036_ (.A(net351),
    .B(_06660_),
    .Y(\hash.CA1.S1.X[22] ));
 sky130_fd_sc_hd__nor4_1 _18037_ (.A(net351),
    .B(_06647_),
    .C(_06649_),
    .D(_06653_),
    .Y(_06661_));
 sky130_fd_sc_hd__xor2_1 _18038_ (.A(\hash.CA1.S1.X[22] ),
    .B(_06661_),
    .X(_00795_));
 sky130_fd_sc_hd__a21o_1 _18039_ (.A1(_13493_),
    .A2(_13488_),
    .B1(_13492_),
    .X(_06662_));
 sky130_fd_sc_hd__a31oi_2 _18040_ (.A1(_13495_),
    .A2(_13499_),
    .A3(_06652_),
    .B1(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__xnor2_2 _18041_ (.A(_13497_),
    .B(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand2_8 _18042_ (.A(_06002_),
    .B(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__inv_4 _18043_ (.A(_06665_),
    .Y(\hash.CA1.S1.X[23] ));
 sky130_fd_sc_hd__nand3_2 _18044_ (.A(\hash.CA1.S1.X[20] ),
    .B(\hash.CA1.S1.X[21] ),
    .C(\hash.CA1.S1.X[22] ),
    .Y(_06666_));
 sky130_fd_sc_hd__nor2_1 _18045_ (.A(_06654_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__xnor2_1 _18046_ (.A(_06665_),
    .B(_06667_),
    .Y(_00796_));
 sky130_fd_sc_hd__o21ai_2 _18047_ (.A1(_06627_),
    .A2(_06629_),
    .B1(_06657_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_1 _18048_ (.A(_13499_),
    .B(_13503_),
    .Y(_06669_));
 sky130_fd_sc_hd__nor2_2 _18049_ (.A(_06658_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__a221oi_4 _18050_ (.A1(_13497_),
    .A2(_13492_),
    .B1(_06668_),
    .B2(_06670_),
    .C1(_13496_),
    .Y(_06671_));
 sky130_fd_sc_hd__xnor2_1 _18051_ (.A(_13501_),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__nor2_4 _18052_ (.A(net354),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__inv_1 _18053_ (.A(_06673_),
    .Y(\hash.CA1.S1.X[24] ));
 sky130_fd_sc_hd__o31ai_2 _18054_ (.A1(_06649_),
    .A2(_06665_),
    .A3(_06666_),
    .B1(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__or4_1 _18055_ (.A(_06649_),
    .B(_06665_),
    .C(_06666_),
    .D(_06673_),
    .X(_06675_));
 sky130_fd_sc_hd__nand2_1 _18056_ (.A(_06674_),
    .B(_06675_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand3_2 _18057_ (.A(_13495_),
    .B(_13499_),
    .C(_13503_),
    .Y(_06676_));
 sky130_fd_sc_hd__a211oi_2 _18058_ (.A1(_06639_),
    .A2(_06637_),
    .B1(_06650_),
    .C1(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand2_1 _18059_ (.A(_13503_),
    .B(_06662_),
    .Y(_06678_));
 sky130_fd_sc_hd__o21ai_1 _18060_ (.A1(_06651_),
    .A2(_06676_),
    .B1(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__or3_1 _18061_ (.A(_13496_),
    .B(_06677_),
    .C(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__a21oi_2 _18062_ (.A1(_06680_),
    .A2(_13501_),
    .B1(_13500_),
    .Y(_06681_));
 sky130_fd_sc_hd__xor2_2 _18063_ (.A(_06681_),
    .B(_13505_),
    .X(_06682_));
 sky130_fd_sc_hd__nor2_4 _18064_ (.A(net351),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1138 ();
 sky130_fd_sc_hd__o31ai_2 _18066_ (.A1(_06654_),
    .A2(_06665_),
    .A3(_06666_),
    .B1(_06673_),
    .Y(_06684_));
 sky130_fd_sc_hd__xor2_1 _18067_ (.A(net1052),
    .B(_06684_),
    .X(_00798_));
 sky130_fd_sc_hd__nand2_1 _18068_ (.A(_13501_),
    .B(_13509_),
    .Y(_06685_));
 sky130_fd_sc_hd__a21oi_1 _18069_ (.A1(_13505_),
    .A2(_13500_),
    .B1(_13504_),
    .Y(_06686_));
 sky130_fd_sc_hd__o21ai_1 _18070_ (.A1(_06671_),
    .A2(_06685_),
    .B1(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__xnor2_2 _18071_ (.A(_13507_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__nor2_4 _18072_ (.A(_06688_),
    .B(net352),
    .Y(_06689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1137 ();
 sky130_fd_sc_hd__nand2_1 _18074_ (.A(_06674_),
    .B(net1052),
    .Y(_06690_));
 sky130_fd_sc_hd__xnor2_1 _18075_ (.A(net1054),
    .B(_06690_),
    .Y(_00799_));
 sky130_fd_sc_hd__a21o_1 _18076_ (.A1(_13507_),
    .A2(_13504_),
    .B1(_13506_),
    .X(_06691_));
 sky130_fd_sc_hd__or3_1 _18077_ (.A(_13496_),
    .B(_13500_),
    .C(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__or3_4 _18078_ (.A(_06677_),
    .B(_06679_),
    .C(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__a21oi_1 _18079_ (.A1(_13509_),
    .A2(_13513_),
    .B1(_06691_),
    .Y(_06694_));
 sky130_fd_sc_hd__nor3_1 _18080_ (.A(_13501_),
    .B(_13500_),
    .C(_06691_),
    .Y(_06695_));
 sky130_fd_sc_hd__nor2_1 _18081_ (.A(_06694_),
    .B(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(_06693_),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__xor2_1 _18083_ (.A(_13511_),
    .B(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__nor2_4 _18084_ (.A(net352),
    .B(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1136 ();
 sky130_fd_sc_hd__nand3_1 _18086_ (.A(net1052),
    .B(_06684_),
    .C(net1054),
    .Y(_06700_));
 sky130_fd_sc_hd__xnor2_1 _18087_ (.A(_06699_),
    .B(_06700_),
    .Y(_00800_));
 sky130_fd_sc_hd__nor2b_1 _18088_ (.A(_06686_),
    .B_N(_13507_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand3_1 _18089_ (.A(_13507_),
    .B(_13501_),
    .C(_13509_),
    .Y(_06702_));
 sky130_fd_sc_hd__nor2_1 _18090_ (.A(_06671_),
    .B(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__o31a_1 _18091_ (.A1(_13506_),
    .A2(_06701_),
    .A3(_06703_),
    .B1(_13511_),
    .X(_06704_));
 sky130_fd_sc_hd__o21ai_2 _18092_ (.A1(_13510_),
    .A2(_06704_),
    .B1(_13515_),
    .Y(_06705_));
 sky130_fd_sc_hd__or3_1 _18093_ (.A(net352),
    .B(_13515_),
    .C(_13510_),
    .X(_06706_));
 sky130_fd_sc_hd__o22a_4 _18094_ (.A1(net352),
    .A2(_06705_),
    .B1(_06706_),
    .B2(_06704_),
    .X(_06707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1135 ();
 sky130_fd_sc_hd__nand4_1 _18096_ (.A(_06674_),
    .B(net1052),
    .C(net1054),
    .D(_06699_),
    .Y(_06708_));
 sky130_fd_sc_hd__xor2_1 _18097_ (.A(_06707_),
    .B(_06708_),
    .X(_00801_));
 sky130_fd_sc_hd__a31o_1 _18098_ (.A1(_13511_),
    .A2(_06693_),
    .A3(_06696_),
    .B1(_13510_),
    .X(_06709_));
 sky130_fd_sc_hd__a21oi_4 _18099_ (.A1(_06709_),
    .A2(_13515_),
    .B1(_13514_),
    .Y(_06710_));
 sky130_fd_sc_hd__xnor2_2 _18100_ (.A(_13517_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_4 _18101_ (.A(_06002_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__inv_6 _18102_ (.A(_06712_),
    .Y(\hash.CA1.S1.X[29] ));
 sky130_fd_sc_hd__a41oi_1 _18103_ (.A1(net1053),
    .A2(_06684_),
    .A3(_06689_),
    .A4(_06699_),
    .B1(_06707_),
    .Y(_06713_));
 sky130_fd_sc_hd__xnor2_1 _18104_ (.A(\hash.CA1.S1.X[29] ),
    .B(_06713_),
    .Y(_00802_));
 sky130_fd_sc_hd__nor4_2 _18105_ (.A(net352),
    .B(_13519_),
    .C(_13514_),
    .D(_13516_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand3_1 _18106_ (.A(_06002_),
    .B(_13517_),
    .C(_13519_),
    .Y(_06715_));
 sky130_fd_sc_hd__nor2_2 _18107_ (.A(_06705_),
    .B(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__nor4_1 _18108_ (.A(net352),
    .B(_13517_),
    .C(_13519_),
    .D(_13516_),
    .Y(_06717_));
 sky130_fd_sc_hd__a31oi_1 _18109_ (.A1(_06002_),
    .A2(_13519_),
    .A3(_13516_),
    .B1(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__nand4_1 _18110_ (.A(_06002_),
    .B(_13517_),
    .C(_13519_),
    .D(_13514_),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_2 _18111_ (.A(_06718_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__a211oi_4 _18112_ (.A1(net1050),
    .A2(_06714_),
    .B1(_06720_),
    .C1(_06716_),
    .Y(\hash.CA1.S1.X[30] ));
 sky130_fd_sc_hd__a41o_1 _18113_ (.A1(_06674_),
    .A2(net1053),
    .A3(net1054),
    .A4(_06699_),
    .B1(_06707_),
    .X(_06721_));
 sky130_fd_sc_hd__nand2_1 _18114_ (.A(_06721_),
    .B(\hash.CA1.S1.X[29] ),
    .Y(_06722_));
 sky130_fd_sc_hd__xor2_1 _18115_ (.A(\hash.CA1.S1.X[30] ),
    .B(_06722_),
    .X(_00804_));
 sky130_fd_sc_hd__nand2_1 _18116_ (.A(_13517_),
    .B(_13519_),
    .Y(_06723_));
 sky130_fd_sc_hd__a21oi_1 _18117_ (.A1(_13519_),
    .A2(_13516_),
    .B1(_13518_),
    .Y(_06724_));
 sky130_fd_sc_hd__o21ai_2 _18118_ (.A1(_06723_),
    .A2(_06710_),
    .B1(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__xnor2_2 _18119_ (.A(\hash.CA2.p5[31] ),
    .B(_06248_),
    .Y(_06726_));
 sky130_fd_sc_hd__xnor2_2 _18120_ (.A(_06725_),
    .B(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__nor2_4 _18121_ (.A(net352),
    .B(_06727_),
    .Y(\hash.CA1.S1.X[31] ));
 sky130_fd_sc_hd__o21ba_1 _18122_ (.A1(_06712_),
    .A2(_06713_),
    .B1_N(\hash.CA1.S1.X[30] ),
    .X(_06728_));
 sky130_fd_sc_hd__xnor2_1 _18123_ (.A(\hash.CA1.S1.X[31] ),
    .B(_06728_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand2_4 _18124_ (.A(_06002_),
    .B(\hash.CA2.b_dash[2] ),
    .Y(_12666_));
 sky130_fd_sc_hd__clkinv_1 _18125_ (.A(_12666_),
    .Y(_13857_));
 sky130_fd_sc_hd__nor2_4 _18126_ (.A(net355),
    .B(\hash.CA2.b_dash[3] ),
    .Y(_12674_));
 sky130_fd_sc_hd__xor2_1 _18127_ (.A(_13858_),
    .B(_12674_),
    .X(_00772_));
 sky130_fd_sc_hd__nor2_2 _18128_ (.A(net355),
    .B(\hash.CA2.b_dash[4] ),
    .Y(_12679_));
 sky130_fd_sc_hd__a21oi_1 _18129_ (.A1(\hash.CA2.b_dash[1] ),
    .A2(\hash.CA2.b_dash[2] ),
    .B1(\hash.CA2.b_dash[3] ),
    .Y(_06729_));
 sky130_fd_sc_hd__xnor2_1 _18130_ (.A(\hash.CA2.b_dash[4] ),
    .B(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__nand2_1 _18131_ (.A(_06002_),
    .B(_06730_),
    .Y(_00774_));
 sky130_fd_sc_hd__or2_4 _18132_ (.A(net355),
    .B(\hash.CA2.b_dash[5] ),
    .X(_12684_));
 sky130_fd_sc_hd__nor4_1 _18133_ (.A(net355),
    .B(\hash.CA2.b_dash[3] ),
    .C(\hash.CA2.b_dash[4] ),
    .D(_13858_),
    .Y(_06731_));
 sky130_fd_sc_hd__xor2_2 _18134_ (.A(_12684_),
    .B(_06731_),
    .X(_00775_));
 sky130_fd_sc_hd__nand2b_4 _18135_ (.A_N(net355),
    .B(\hash.CA2.b_dash[6] ),
    .Y(_12692_));
 sky130_fd_sc_hd__nor3_2 _18136_ (.A(net355),
    .B(\hash.CA2.b_dash[3] ),
    .C(\hash.CA2.b_dash[4] ),
    .Y(_06732_));
 sky130_fd_sc_hd__a21oi_2 _18137_ (.A1(\hash.CA2.b_dash[1] ),
    .A2(\hash.CA2.b_dash[2] ),
    .B1(\hash.CA2.b_dash[5] ),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_1 _18138_ (.A(_06732_),
    .B(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__xnor2_1 _18139_ (.A(_12692_),
    .B(_06734_),
    .Y(_00776_));
 sky130_fd_sc_hd__nor4_2 _18140_ (.A(\hash.CA2.b_dash[3] ),
    .B(\hash.CA2.b_dash[4] ),
    .C(\hash.CA2.b_dash[5] ),
    .D(_13858_),
    .Y(_06735_));
 sky130_fd_sc_hd__nor2_4 _18141_ (.A(_12692_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_8 _18142_ (.A(_06002_),
    .B(\hash.CA2.b_dash[7] ),
    .Y(_12701_));
 sky130_fd_sc_hd__inv_2 _18143_ (.A(\hash.CA2.b_dash[7] ),
    .Y(_06737_));
 sky130_fd_sc_hd__nand2_1 _18144_ (.A(_06737_),
    .B(_06736_),
    .Y(_06738_));
 sky130_fd_sc_hd__o21ai_1 _18145_ (.A1(_06736_),
    .A2(_12701_),
    .B1(_06738_),
    .Y(_00777_));
 sky130_fd_sc_hd__nor2_4 _18146_ (.A(net351),
    .B(\hash.CA2.b_dash[8] ),
    .Y(_12708_));
 sky130_fd_sc_hd__a211oi_4 _18147_ (.A1(_06732_),
    .A2(_06733_),
    .B1(_12692_),
    .C1(_06737_),
    .Y(_06739_));
 sky130_fd_sc_hd__xor2_2 _18148_ (.A(_12708_),
    .B(_06739_),
    .X(_00778_));
 sky130_fd_sc_hd__clkinv_1 _18149_ (.A(\hash.CA2.b_dash[9] ),
    .Y(_06740_));
 sky130_fd_sc_hd__a21oi_4 _18150_ (.A1(\hash.CA2.b_dash[7] ),
    .A2(_06736_),
    .B1(\hash.CA2.b_dash[8] ),
    .Y(_06741_));
 sky130_fd_sc_hd__xnor2_1 _18151_ (.A(_06740_),
    .B(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_1 _18152_ (.A(_06002_),
    .B(_06742_),
    .Y(_00779_));
 sky130_fd_sc_hd__nor2_4 _18153_ (.A(net352),
    .B(\hash.CA2.b_dash[10] ),
    .Y(_12723_));
 sky130_fd_sc_hd__nand2_8 _18154_ (.A(_06002_),
    .B(\hash.CA2.b_dash[9] ),
    .Y(_12714_));
 sky130_fd_sc_hd__nor2_2 _18155_ (.A(\hash.CA2.b_dash[8] ),
    .B(_06739_),
    .Y(_06743_));
 sky130_fd_sc_hd__nor2_4 _18156_ (.A(_12714_),
    .B(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__mux2_1 _18157_ (.A0(_12723_),
    .A1(\hash.CA2.b_dash[10] ),
    .S(_06744_),
    .X(_00780_));
 sky130_fd_sc_hd__nand2_4 _18158_ (.A(_06002_),
    .B(\hash.CA2.b_dash[11] ),
    .Y(_06745_));
 sky130_fd_sc_hd__inv_8 _18159_ (.A(_06745_),
    .Y(_12732_));
 sky130_fd_sc_hd__o21ai_2 _18160_ (.A1(_06740_),
    .A2(_06741_),
    .B1(_12723_),
    .Y(_06746_));
 sky130_fd_sc_hd__xnor2_1 _18161_ (.A(_06745_),
    .B(_06746_),
    .Y(_00752_));
 sky130_fd_sc_hd__or2_4 _18162_ (.A(net352),
    .B(\hash.CA2.b_dash[12] ),
    .X(_06747_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1134 ();
 sky130_fd_sc_hd__inv_1 _18164_ (.A(\hash.CA2.b_dash[10] ),
    .Y(_06748_));
 sky130_fd_sc_hd__o21ai_4 _18165_ (.A1(\hash.CA2.b_dash[8] ),
    .A2(_06739_),
    .B1(\hash.CA2.b_dash[9] ),
    .Y(_06749_));
 sky130_fd_sc_hd__a21oi_1 _18166_ (.A1(_06748_),
    .A2(_06749_),
    .B1(_06745_),
    .Y(_06750_));
 sky130_fd_sc_hd__xnor2_1 _18167_ (.A(_06747_),
    .B(_06750_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_2 _18168_ (.A(\hash.CA2.b_dash[7] ),
    .B(_06736_),
    .Y(_06751_));
 sky130_fd_sc_hd__a21oi_4 _18169_ (.A1(_12708_),
    .A2(_06751_),
    .B1(_12714_),
    .Y(_06752_));
 sky130_fd_sc_hd__o21a_1 _18170_ (.A1(\hash.CA2.b_dash[10] ),
    .A2(_06752_),
    .B1(\hash.CA2.b_dash[11] ),
    .X(_06753_));
 sky130_fd_sc_hd__nor2_1 _18171_ (.A(_06747_),
    .B(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__or2_4 _18172_ (.A(net352),
    .B(\hash.CA2.b_dash[13] ),
    .X(_12746_));
 sky130_fd_sc_hd__nor2_1 _18173_ (.A(_06754_),
    .B(_12746_),
    .Y(_06755_));
 sky130_fd_sc_hd__a21oi_1 _18174_ (.A1(\hash.CA2.b_dash[13] ),
    .A2(_06754_),
    .B1(_06755_),
    .Y(_00754_));
 sky130_fd_sc_hd__nor2_4 _18175_ (.A(net352),
    .B(\hash.CA2.b_dash[14] ),
    .Y(_12752_));
 sky130_fd_sc_hd__o21ai_0 _18176_ (.A1(\hash.CA2.b_dash[10] ),
    .A2(_06744_),
    .B1(\hash.CA2.b_dash[11] ),
    .Y(_06756_));
 sky130_fd_sc_hd__nor2_1 _18177_ (.A(\hash.CA2.b_dash[13] ),
    .B(_06747_),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_1 _18178_ (.A(_06756_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__xor2_1 _18179_ (.A(_12752_),
    .B(_06758_),
    .X(_00755_));
 sky130_fd_sc_hd__nor2_2 _18180_ (.A(net353),
    .B(\hash.CA2.b_dash[15] ),
    .Y(_12759_));
 sky130_fd_sc_hd__nor2_1 _18181_ (.A(\hash.CA2.b_dash[12] ),
    .B(\hash.CA2.b_dash[13] ),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_1 _18182_ (.A(_12752_),
    .B(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__a21oi_2 _18183_ (.A1(_12732_),
    .A2(_06746_),
    .B1(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nor3_1 _18184_ (.A(net352),
    .B(\hash.CA2.b_dash[15] ),
    .C(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__a21oi_1 _18185_ (.A1(\hash.CA2.b_dash[15] ),
    .A2(_06761_),
    .B1(_06762_),
    .Y(_00756_));
 sky130_fd_sc_hd__or2_4 _18186_ (.A(net352),
    .B(\hash.CA2.b_dash[16] ),
    .X(_12767_));
 sky130_fd_sc_hd__or2_4 _18187_ (.A(_06750_),
    .B(_06760_),
    .X(_06763_));
 sky130_fd_sc_hd__nor2_1 _18188_ (.A(\hash.CA2.b_dash[15] ),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__xor2_1 _18189_ (.A(_12767_),
    .B(_06764_),
    .X(_00757_));
 sky130_fd_sc_hd__nor2_4 _18190_ (.A(net352),
    .B(\hash.CA2.b_dash[17] ),
    .Y(_06765_));
 sky130_fd_sc_hd__inv_8 _18191_ (.A(_06765_),
    .Y(_12774_));
 sky130_fd_sc_hd__nor4_1 _18192_ (.A(net352),
    .B(\hash.CA2.b_dash[14] ),
    .C(\hash.CA2.b_dash[15] ),
    .D(\hash.CA2.b_dash[16] ),
    .Y(_06766_));
 sky130_fd_sc_hd__nand3b_1 _18193_ (.A_N(\hash.CA2.b_dash[13] ),
    .B(_06754_),
    .C(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__xnor2_1 _18194_ (.A(_12774_),
    .B(_06767_),
    .Y(_00758_));
 sky130_fd_sc_hd__or2_4 _18195_ (.A(net352),
    .B(\hash.CA2.b_dash[18] ),
    .X(_12780_));
 sky130_fd_sc_hd__nor3b_1 _18196_ (.A(\hash.CA2.b_dash[17] ),
    .B(_06758_),
    .C_N(_06766_),
    .Y(_06768_));
 sky130_fd_sc_hd__xor2_1 _18197_ (.A(_12780_),
    .B(_06768_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_4 _18198_ (.A(net352),
    .B(\hash.CA2.b_dash[19] ),
    .X(_12786_));
 sky130_fd_sc_hd__nor4_1 _18199_ (.A(net352),
    .B(\hash.CA2.b_dash[15] ),
    .C(\hash.CA2.b_dash[16] ),
    .D(\hash.CA2.b_dash[18] ),
    .Y(_06769_));
 sky130_fd_sc_hd__nand3_2 _18200_ (.A(_06761_),
    .B(_06765_),
    .C(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__xnor2_1 _18201_ (.A(_12786_),
    .B(_06770_),
    .Y(_00760_));
 sky130_fd_sc_hd__nor2b_4 _18202_ (.A(net352),
    .B_N(\hash.CA2.b_dash[20] ),
    .Y(_06771_));
 sky130_fd_sc_hd__nor4b_4 _18203_ (.A(\hash.CA2.b_dash[17] ),
    .B(_06763_),
    .C(_12786_),
    .D_N(_06769_),
    .Y(_06772_));
 sky130_fd_sc_hd__xnor2_1 _18204_ (.A(_06771_),
    .B(_06772_),
    .Y(_00761_));
 sky130_fd_sc_hd__nor2b_2 _18205_ (.A(net353),
    .B_N(\hash.CA2.b_dash[21] ),
    .Y(_12802_));
 sky130_fd_sc_hd__o21a_4 _18206_ (.A1(\hash.CA2.b_dash[19] ),
    .A2(_06770_),
    .B1(\hash.CA2.b_dash[20] ),
    .X(_06773_));
 sky130_fd_sc_hd__xnor2_1 _18207_ (.A(\hash.CA2.b_dash[21] ),
    .B(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__nor2_1 _18208_ (.A(net352),
    .B(_06774_),
    .Y(_00762_));
 sky130_fd_sc_hd__nor2_4 _18209_ (.A(net353),
    .B(\hash.CA2.b_dash[22] ),
    .Y(_12810_));
 sky130_fd_sc_hd__nand3b_1 _18210_ (.A_N(_06772_),
    .B(_06771_),
    .C(\hash.CA2.b_dash[21] ),
    .Y(_06775_));
 sky130_fd_sc_hd__xnor2_1 _18211_ (.A(_12810_),
    .B(_06775_),
    .Y(_00763_));
 sky130_fd_sc_hd__nor2b_4 _18212_ (.A(net353),
    .B_N(\hash.CA2.b_dash[23] ),
    .Y(_12818_));
 sky130_fd_sc_hd__a211o_4 _18213_ (.A1(\hash.CA2.b_dash[21] ),
    .A2(_06773_),
    .B1(\hash.CA2.b_dash[22] ),
    .C1(net354),
    .X(_06776_));
 sky130_fd_sc_hd__xor2_1 _18214_ (.A(_12818_),
    .B(_06776_),
    .X(_00764_));
 sky130_fd_sc_hd__nor2_4 _18215_ (.A(net353),
    .B(\hash.CA2.b_dash[24] ),
    .Y(_12826_));
 sky130_fd_sc_hd__nand2b_1 _18216_ (.A_N(\hash.CA2.b_dash[22] ),
    .B(_06775_),
    .Y(_06777_));
 sky130_fd_sc_hd__nand2_1 _18217_ (.A(_12818_),
    .B(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__xnor2_1 _18218_ (.A(_12826_),
    .B(_06778_),
    .Y(_00765_));
 sky130_fd_sc_hd__nor2_4 _18219_ (.A(net353),
    .B(_04733_),
    .Y(_12834_));
 sky130_fd_sc_hd__a21boi_0 _18220_ (.A1(_12818_),
    .A2(_06776_),
    .B1_N(_12826_),
    .Y(_06779_));
 sky130_fd_sc_hd__xnor2_1 _18221_ (.A(_12834_),
    .B(_06779_),
    .Y(_00766_));
 sky130_fd_sc_hd__a21o_1 _18222_ (.A1(\hash.CA2.b_dash[23] ),
    .A2(_06777_),
    .B1(\hash.CA2.b_dash[24] ),
    .X(_06780_));
 sky130_fd_sc_hd__nand2_2 _18223_ (.A(_12834_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__nor2_4 _18224_ (.A(net354),
    .B(\hash.CA2.b_dash[26] ),
    .Y(_06782_));
 sky130_fd_sc_hd__xnor2_1 _18225_ (.A(_06781_),
    .B(_06782_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2b_4 _18226_ (.A(net353),
    .B_N(\hash.CA2.b_dash[27] ),
    .Y(_12849_));
 sky130_fd_sc_hd__a21oi_1 _18227_ (.A1(\hash.CA2.b_dash[23] ),
    .A2(_06776_),
    .B1(\hash.CA2.b_dash[24] ),
    .Y(_06783_));
 sky130_fd_sc_hd__o21ai_2 _18228_ (.A1(_04733_),
    .A2(_06783_),
    .B1(_06782_),
    .Y(_06784_));
 sky130_fd_sc_hd__xor2_1 _18229_ (.A(_12849_),
    .B(_06784_),
    .X(_00768_));
 sky130_fd_sc_hd__inv_1 _18230_ (.A(\hash.CA2.b_dash[28] ),
    .Y(_06785_));
 sky130_fd_sc_hd__nor2_2 _18231_ (.A(net353),
    .B(_06785_),
    .Y(_12857_));
 sky130_fd_sc_hd__a21boi_2 _18232_ (.A1(_06781_),
    .A2(_06782_),
    .B1_N(_12849_),
    .Y(_06786_));
 sky130_fd_sc_hd__mux2_1 _18233_ (.A0(_12857_),
    .A1(_06785_),
    .S(_06786_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_4 _18234_ (.A(net353),
    .B(\hash.CA2.b_dash[29] ),
    .X(_12864_));
 sky130_fd_sc_hd__and3_4 _18235_ (.A(\hash.CA2.b_dash[28] ),
    .B(_12849_),
    .C(_06784_),
    .X(_06787_));
 sky130_fd_sc_hd__xnor2_1 _18236_ (.A(_12864_),
    .B(_06787_),
    .Y(_00770_));
 sky130_fd_sc_hd__nor2b_4 _18237_ (.A(net353),
    .B_N(\hash.CA2.b_dash[30] ),
    .Y(_12871_));
 sky130_fd_sc_hd__a21oi_1 _18238_ (.A1(\hash.CA2.b_dash[28] ),
    .A2(_06786_),
    .B1(\hash.CA2.b_dash[29] ),
    .Y(_06788_));
 sky130_fd_sc_hd__xor2_1 _18239_ (.A(\hash.CA2.b_dash[30] ),
    .B(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__nand2_1 _18240_ (.A(_06002_),
    .B(_06789_),
    .Y(_00771_));
 sky130_fd_sc_hd__o21ai_0 _18241_ (.A1(\hash.CA2.b_dash[29] ),
    .A2(_06787_),
    .B1(\hash.CA2.b_dash[30] ),
    .Y(_06790_));
 sky130_fd_sc_hd__xnor2_1 _18242_ (.A(\hash.CA2.b_dash[31] ),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__nor2_1 _18243_ (.A(net353),
    .B(_06791_),
    .Y(_00773_));
 sky130_fd_sc_hd__xor2_1 _18244_ (.A(_13859_),
    .B(_13679_),
    .X(_00742_));
 sky130_fd_sc_hd__nand3_4 _18245_ (.A(\hash.CA2.a_dash[1] ),
    .B(\hash.CA2.a_dash[2] ),
    .C(\hash.CA2.a_dash[3] ),
    .Y(_06792_));
 sky130_fd_sc_hd__xnor2_1 _18246_ (.A(\hash.CA2.a_dash[4] ),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__nor2_1 _18247_ (.A(net349),
    .B(_06793_),
    .Y(_00744_));
 sky130_fd_sc_hd__or2_4 _18248_ (.A(net349),
    .B(\hash.CA2.a_dash[4] ),
    .X(_13685_));
 sky130_fd_sc_hd__a21oi_1 _18249_ (.A1(\hash.CA2.a_dash[3] ),
    .A2(_13859_),
    .B1(\hash.CA2.a_dash[4] ),
    .Y(_06794_));
 sky130_fd_sc_hd__xnor2_1 _18250_ (.A(\hash.CA2.a_dash[5] ),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand2_1 _18251_ (.A(_06002_),
    .B(_06795_),
    .Y(_00745_));
 sky130_fd_sc_hd__nor2_4 _18252_ (.A(\hash.CA2.a_dash[5] ),
    .B(_13685_),
    .Y(_06796_));
 sky130_fd_sc_hd__nand2_4 _18253_ (.A(_06792_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__xnor2_2 _18254_ (.A(_13697_),
    .B(_06797_),
    .Y(_00746_));
 sky130_fd_sc_hd__a21oi_1 _18255_ (.A1(\hash.CA2.a_dash[3] ),
    .A2(_13859_),
    .B1(\hash.CA2.a_dash[6] ),
    .Y(_06798_));
 sky130_fd_sc_hd__nand2_4 _18256_ (.A(_06796_),
    .B(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__nand2_4 _18257_ (.A(_06002_),
    .B(\hash.CA2.a_dash[7] ),
    .Y(_06800_));
 sky130_fd_sc_hd__xnor2_2 _18258_ (.A(_06799_),
    .B(_06800_),
    .Y(_00747_));
 sky130_fd_sc_hd__or2_0 _18259_ (.A(net350),
    .B(\hash.CA2.a_dash[8] ),
    .X(_13710_));
 sky130_fd_sc_hd__o21ai_0 _18260_ (.A1(\hash.CA2.a_dash[6] ),
    .A2(_06797_),
    .B1(\hash.CA2.a_dash[7] ),
    .Y(_06801_));
 sky130_fd_sc_hd__xnor2_1 _18261_ (.A(\hash.CA2.a_dash[8] ),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__nor2_1 _18262_ (.A(net349),
    .B(_06802_),
    .Y(_00748_));
 sky130_fd_sc_hd__a21oi_2 _18263_ (.A1(\hash.CA2.a_dash[7] ),
    .A2(_06799_),
    .B1(\hash.CA2.a_dash[8] ),
    .Y(_06803_));
 sky130_fd_sc_hd__xnor2_2 _18264_ (.A(\hash.CA2.a_dash[9] ),
    .B(_06803_),
    .Y(_06804_));
 sky130_fd_sc_hd__nand2_1 _18265_ (.A(_06002_),
    .B(_06804_),
    .Y(_00749_));
 sky130_fd_sc_hd__nor2b_4 _18266_ (.A(net350),
    .B_N(\hash.CA2.a_dash[10] ),
    .Y(_13721_));
 sky130_fd_sc_hd__nor2_1 _18267_ (.A(\hash.CA2.a_dash[6] ),
    .B(_06797_),
    .Y(_06805_));
 sky130_fd_sc_hd__nor2_1 _18268_ (.A(\hash.CA2.a_dash[8] ),
    .B(_13716_),
    .Y(_06806_));
 sky130_fd_sc_hd__o21ai_2 _18269_ (.A1(_06800_),
    .A2(_06805_),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__xor2_2 _18270_ (.A(_13721_),
    .B(_06807_),
    .X(_00750_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1133 ();
 sky130_fd_sc_hd__clkinv_2 _18272_ (.A(_06803_),
    .Y(_06809_));
 sky130_fd_sc_hd__o21ai_2 _18273_ (.A1(\hash.CA2.a_dash[9] ),
    .A2(_06809_),
    .B1(\hash.CA2.a_dash[10] ),
    .Y(_06810_));
 sky130_fd_sc_hd__xor2_2 _18274_ (.A(\hash.CA2.a_dash[11] ),
    .B(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__nor2_1 _18275_ (.A(net351),
    .B(_06811_),
    .Y(_00722_));
 sky130_fd_sc_hd__or2_4 _18276_ (.A(net350),
    .B(\hash.CA2.a_dash[12] ),
    .X(_13734_));
 sky130_fd_sc_hd__and3_4 _18277_ (.A(\hash.CA2.a_dash[11] ),
    .B(_13721_),
    .C(_06807_),
    .X(_06812_));
 sky130_fd_sc_hd__xnor2_1 _18278_ (.A(_13734_),
    .B(_06812_),
    .Y(_00723_));
 sky130_fd_sc_hd__o211a_4 _18279_ (.A1(_13716_),
    .A2(_06809_),
    .B1(_13721_),
    .C1(\hash.CA2.a_dash[11] ),
    .X(_06813_));
 sky130_fd_sc_hd__or3_4 _18280_ (.A(\hash.CA2.a_dash[12] ),
    .B(\hash.CA2.a_dash[13] ),
    .C(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__o21ai_2 _18281_ (.A1(\hash.CA2.a_dash[12] ),
    .A2(_06813_),
    .B1(\hash.CA2.a_dash[13] ),
    .Y(_06815_));
 sky130_fd_sc_hd__nand3_4 _18282_ (.A(_06002_),
    .B(_06814_),
    .C(_06815_),
    .Y(_00724_));
 sky130_fd_sc_hd__or3_4 _18283_ (.A(net350),
    .B(\hash.CA2.a_dash[12] ),
    .C(\hash.CA2.a_dash[13] ),
    .X(_06816_));
 sky130_fd_sc_hd__nor2_1 _18284_ (.A(_06812_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__xor2_1 _18285_ (.A(_13746_),
    .B(_06817_),
    .X(_00725_));
 sky130_fd_sc_hd__or3_4 _18286_ (.A(\hash.CA2.a_dash[14] ),
    .B(_06813_),
    .C(_06816_),
    .X(_06818_));
 sky130_fd_sc_hd__xnor2_1 _18287_ (.A(_13753_),
    .B(_06818_),
    .Y(_00726_));
 sky130_fd_sc_hd__nor2b_4 _18288_ (.A(net350),
    .B_N(\hash.CA2.a_dash[16] ),
    .Y(_13760_));
 sky130_fd_sc_hd__or4_4 _18289_ (.A(\hash.CA2.a_dash[15] ),
    .B(_13746_),
    .C(_06812_),
    .D(_06816_),
    .X(_06819_));
 sky130_fd_sc_hd__xor2_1 _18290_ (.A(_13760_),
    .B(_06819_),
    .X(_00727_));
 sky130_fd_sc_hd__nor2_1 _18291_ (.A(net351),
    .B(\hash.CA2.a_dash[17] ),
    .Y(_06820_));
 sky130_fd_sc_hd__clkinv_1 _18292_ (.A(_06820_),
    .Y(_13767_));
 sky130_fd_sc_hd__o21ai_2 _18293_ (.A1(\hash.CA2.a_dash[15] ),
    .A2(_06818_),
    .B1(_13760_),
    .Y(_06821_));
 sky130_fd_sc_hd__mux2_1 _18294_ (.A0(\hash.CA2.a_dash[17] ),
    .A1(_06820_),
    .S(_06821_),
    .X(_00728_));
 sky130_fd_sc_hd__or2_0 _18295_ (.A(net350),
    .B(\hash.CA2.a_dash[18] ),
    .X(_13773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1132 ();
 sky130_fd_sc_hd__a21oi_1 _18297_ (.A1(\hash.CA2.a_dash[16] ),
    .A2(_06819_),
    .B1(\hash.CA2.a_dash[17] ),
    .Y(_06823_));
 sky130_fd_sc_hd__xnor2_1 _18298_ (.A(\hash.CA2.a_dash[18] ),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__nand2_1 _18299_ (.A(_06002_),
    .B(_06824_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand3b_1 _18300_ (.A_N(\hash.CA2.a_dash[18] ),
    .B(_06820_),
    .C(_06821_),
    .Y(_06825_));
 sky130_fd_sc_hd__xnor2_1 _18301_ (.A(_13778_),
    .B(_06825_),
    .Y(_00730_));
 sky130_fd_sc_hd__nor2b_2 _18302_ (.A(net351),
    .B_N(\hash.CA2.a_dash[20] ),
    .Y(_13783_));
 sky130_fd_sc_hd__nand2_1 _18303_ (.A(\hash.CA2.a_dash[16] ),
    .B(_06819_),
    .Y(_06826_));
 sky130_fd_sc_hd__nor3_1 _18304_ (.A(\hash.CA2.a_dash[18] ),
    .B(\hash.CA2.a_dash[19] ),
    .C(_13767_),
    .Y(_06827_));
 sky130_fd_sc_hd__nand2_2 _18305_ (.A(_06826_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__xor2_1 _18306_ (.A(_13783_),
    .B(_06828_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_0 _18307_ (.A(net351),
    .B(\hash.CA2.a_dash[21] ),
    .X(_13788_));
 sky130_fd_sc_hd__a21boi_2 _18308_ (.A1(_06821_),
    .A2(_06827_),
    .B1_N(\hash.CA2.a_dash[20] ),
    .Y(_06829_));
 sky130_fd_sc_hd__xor2_1 _18309_ (.A(\hash.CA2.a_dash[21] ),
    .B(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__nor2_1 _18310_ (.A(net352),
    .B(_06830_),
    .Y(_00732_));
 sky130_fd_sc_hd__or2_4 _18311_ (.A(net351),
    .B(\hash.CA2.a_dash[22] ),
    .X(_13793_));
 sky130_fd_sc_hd__a21oi_2 _18312_ (.A1(\hash.CA2.a_dash[20] ),
    .A2(_06828_),
    .B1(\hash.CA2.a_dash[21] ),
    .Y(_06831_));
 sky130_fd_sc_hd__xnor2_1 _18313_ (.A(\hash.CA2.a_dash[22] ),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2_1 _18314_ (.A(_06002_),
    .B(_06832_),
    .Y(_00733_));
 sky130_fd_sc_hd__nor2b_4 _18315_ (.A(net351),
    .B_N(\hash.CA2.a_dash[23] ),
    .Y(_13799_));
 sky130_fd_sc_hd__or3_4 _18316_ (.A(\hash.CA2.a_dash[21] ),
    .B(_06829_),
    .C(_13793_),
    .X(_06833_));
 sky130_fd_sc_hd__xor2_1 _18317_ (.A(_13799_),
    .B(_06833_),
    .X(_00734_));
 sky130_fd_sc_hd__nand2b_2 _18318_ (.A_N(_13793_),
    .B(_06831_),
    .Y(_06834_));
 sky130_fd_sc_hd__nand2_1 _18319_ (.A(\hash.CA2.a_dash[23] ),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__xor2_1 _18320_ (.A(\hash.CA2.a_dash[24] ),
    .B(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__nor2_1 _18321_ (.A(net352),
    .B(_06836_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand3_1 _18322_ (.A(\hash.CA2.a_dash[23] ),
    .B(\hash.CA2.a_dash[24] ),
    .C(_06833_),
    .Y(_06837_));
 sky130_fd_sc_hd__xnor2_1 _18323_ (.A(_04734_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_1 _18324_ (.A(net352),
    .B(_06838_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand4_1 _18325_ (.A(\hash.CA2.a_dash[24] ),
    .B(\hash.CA2.a_dash[25] ),
    .C(_13799_),
    .D(_06834_),
    .Y(_06839_));
 sky130_fd_sc_hd__xor2_1 _18326_ (.A(_06287_),
    .B(_06839_),
    .X(_00737_));
 sky130_fd_sc_hd__and4_4 _18327_ (.A(\hash.CA2.a_dash[24] ),
    .B(\hash.CA2.a_dash[25] ),
    .C(_13799_),
    .D(_06833_),
    .X(_06840_));
 sky130_fd_sc_hd__or3_1 _18328_ (.A(\hash.CA2.a_dash[26] ),
    .B(\hash.CA2.a_dash[27] ),
    .C(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__o21ai_0 _18329_ (.A1(\hash.CA2.a_dash[26] ),
    .A2(_06840_),
    .B1(\hash.CA2.a_dash[27] ),
    .Y(_06842_));
 sky130_fd_sc_hd__nand3_1 _18330_ (.A(_06002_),
    .B(_06841_),
    .C(_06842_),
    .Y(_00738_));
 sky130_fd_sc_hd__nor2_1 _18331_ (.A(\hash.CA2.a_dash[27] ),
    .B(_06287_),
    .Y(_06843_));
 sky130_fd_sc_hd__nand2_1 _18332_ (.A(_06839_),
    .B(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__xnor2_1 _18333_ (.A(_13834_),
    .B(_06844_),
    .Y(_00739_));
 sky130_fd_sc_hd__or3_4 _18334_ (.A(\hash.CA2.a_dash[27] ),
    .B(\hash.CA2.a_dash[28] ),
    .C(_06287_),
    .X(_06845_));
 sky130_fd_sc_hd__nor2_1 _18335_ (.A(_06840_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__xor2_1 _18336_ (.A(_13840_),
    .B(_06846_),
    .X(_00740_));
 sky130_fd_sc_hd__nor2_2 _18337_ (.A(net352),
    .B(_04769_),
    .Y(_13845_));
 sky130_fd_sc_hd__nor2_1 _18338_ (.A(\hash.CA2.a_dash[29] ),
    .B(_06845_),
    .Y(_06847_));
 sky130_fd_sc_hd__nand2_1 _18339_ (.A(_06839_),
    .B(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__xor2_1 _18340_ (.A(_13845_),
    .B(_06848_),
    .X(_00741_));
 sky130_fd_sc_hd__o31ai_1 _18341_ (.A1(\hash.CA2.a_dash[29] ),
    .A2(_06840_),
    .A3(_06845_),
    .B1(\hash.CA2.a_dash[30] ),
    .Y(_06849_));
 sky130_fd_sc_hd__xor2_1 _18342_ (.A(\hash.CA2.a_dash[31] ),
    .B(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__nor2_1 _18343_ (.A(net352),
    .B(_06850_),
    .Y(_00743_));
 sky130_fd_sc_hd__xnor2_1 _18344_ (.A(_13860_),
    .B(\hash.CA1.b[2] ),
    .Y(_00711_));
 sky130_fd_sc_hd__a21oi_2 _18345_ (.A1(_12922_),
    .A2(_12082_),
    .B1(_04421_),
    .Y(_06851_));
 sky130_fd_sc_hd__xor2_1 _18346_ (.A(_04470_),
    .B(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__nand2_1 _18347_ (.A(_06002_),
    .B(_06852_),
    .Y(_00714_));
 sky130_fd_sc_hd__o21ai_0 _18348_ (.A1(_13860_),
    .A2(_04421_),
    .B1(_04470_),
    .Y(_06853_));
 sky130_fd_sc_hd__xor2_1 _18349_ (.A(_04487_),
    .B(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__nor2_1 _18350_ (.A(net349),
    .B(_06854_),
    .Y(_00715_));
 sky130_fd_sc_hd__and4bb_4 _18351_ (.A_N(net349),
    .B_N(_06851_),
    .C(_04487_),
    .D(_04470_),
    .X(_06855_));
 sky130_fd_sc_hd__xor2_1 _18352_ (.A(\hash.CA1.b[5] ),
    .B(_06855_),
    .X(_00716_));
 sky130_fd_sc_hd__o211a_4 _18353_ (.A1(_13860_),
    .A2(_04421_),
    .B1(_04470_),
    .C1(_04501_),
    .X(_06856_));
 sky130_fd_sc_hd__nand2_1 _18354_ (.A(\hash.CA1.b[4] ),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__xnor2_1 _18355_ (.A(\hash.CA1.b[6] ),
    .B(_06857_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand3_1 _18356_ (.A(_04501_),
    .B(_04522_),
    .C(_06855_),
    .Y(_06858_));
 sky130_fd_sc_hd__xor2_1 _18357_ (.A(\hash.CA1.b[7] ),
    .B(_06858_),
    .X(_00718_));
 sky130_fd_sc_hd__xnor2_1 _18358_ (.A(_12930_),
    .B(_04400_),
    .Y(_06859_));
 sky130_fd_sc_hd__nand3_2 _18359_ (.A(_04487_),
    .B(_06856_),
    .C(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__nand3_2 _18360_ (.A(_06002_),
    .B(_04543_),
    .C(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__nor2_1 _18361_ (.A(_04562_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21oi_2 _18362_ (.A1(_06279_),
    .A2(_06861_),
    .B1(_06862_),
    .Y(_00719_));
 sky130_fd_sc_hd__a31o_1 _18363_ (.A1(_04501_),
    .A2(_04522_),
    .A3(_06855_),
    .B1(_04542_),
    .X(_06863_));
 sky130_fd_sc_hd__and2_4 _18364_ (.A(_06279_),
    .B(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__nand2_1 _18365_ (.A(_04580_),
    .B(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__o21ai_2 _18366_ (.A1(_06280_),
    .A2(_06864_),
    .B1(_06865_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand3_1 _18367_ (.A(\hash.CA1.b[4] ),
    .B(\hash.CA1.b[6] ),
    .C(_06856_),
    .Y(_06866_));
 sky130_fd_sc_hd__nand2_1 _18368_ (.A(_04543_),
    .B(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__a21oi_1 _18369_ (.A1(_04562_),
    .A2(_06867_),
    .B1(_04580_),
    .Y(_06868_));
 sky130_fd_sc_hd__xnor2_2 _18370_ (.A(_04599_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand2_1 _18371_ (.A(_06002_),
    .B(_06869_),
    .Y(_00691_));
 sky130_fd_sc_hd__nor3_1 _18372_ (.A(_04580_),
    .B(\hash.CA1.b[10] ),
    .C(_06864_),
    .Y(_06870_));
 sky130_fd_sc_hd__xnor2_2 _18373_ (.A(_06282_),
    .B(_06870_),
    .Y(_00692_));
 sky130_fd_sc_hd__a2111o_2 _18374_ (.A1(_04562_),
    .A2(_06861_),
    .B1(_06280_),
    .C1(_04614_),
    .D1(_04599_),
    .X(_06871_));
 sky130_fd_sc_hd__xor2_1 _18375_ (.A(_06283_),
    .B(_06871_),
    .X(_00693_));
 sky130_fd_sc_hd__a2111o_2 _18376_ (.A1(_06279_),
    .A2(_06863_),
    .B1(_06280_),
    .C1(_04599_),
    .D1(_04614_),
    .X(_06872_));
 sky130_fd_sc_hd__nand2_1 _18377_ (.A(_04623_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__xnor2_1 _18378_ (.A(_04437_),
    .B(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__nor2_1 _18379_ (.A(net351),
    .B(_06874_),
    .Y(_00694_));
 sky130_fd_sc_hd__a21oi_2 _18380_ (.A1(_04623_),
    .A2(_06871_),
    .B1(_04437_),
    .Y(_06875_));
 sky130_fd_sc_hd__xnor2_1 _18381_ (.A(net1093),
    .B(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__nand2_1 _18382_ (.A(_06002_),
    .B(_06876_),
    .Y(_00695_));
 sky130_fd_sc_hd__a21oi_2 _18383_ (.A1(_06283_),
    .A2(_06872_),
    .B1(_04437_),
    .Y(_06877_));
 sky130_fd_sc_hd__nor3_1 _18384_ (.A(_04475_),
    .B(_04484_),
    .C(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__o21a_1 _18385_ (.A1(_04475_),
    .A2(_06877_),
    .B1(_04484_),
    .X(_06879_));
 sky130_fd_sc_hd__nor3_2 _18386_ (.A(net350),
    .B(_06878_),
    .C(_06879_),
    .Y(_00696_));
 sky130_fd_sc_hd__a21oi_1 _18387_ (.A1(_06283_),
    .A2(_06871_),
    .B1(_04437_),
    .Y(_06880_));
 sky130_fd_sc_hd__nor2_1 _18388_ (.A(_04475_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__nor2_1 _18389_ (.A(_04484_),
    .B(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__xnor2_1 _18390_ (.A(_04503_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_1 _18391_ (.A(_06002_),
    .B(_06883_),
    .Y(_00697_));
 sky130_fd_sc_hd__nor3_2 _18392_ (.A(net350),
    .B(_04484_),
    .C(_04503_),
    .Y(_06884_));
 sky130_fd_sc_hd__o21ai_4 _18393_ (.A1(net1092),
    .A2(_06877_),
    .B1(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__xnor2_1 _18394_ (.A(\hash.CA1.b[17] ),
    .B(_06885_),
    .Y(_00698_));
 sky130_fd_sc_hd__o21ai_2 _18395_ (.A1(net1093),
    .A2(_06875_),
    .B1(_06884_),
    .Y(_06886_));
 sky130_fd_sc_hd__or2_4 _18396_ (.A(_04520_),
    .B(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__xnor2_1 _18397_ (.A(\hash.CA1.b[18] ),
    .B(_06887_),
    .Y(_00699_));
 sky130_fd_sc_hd__nor4_2 _18398_ (.A(net351),
    .B(_04520_),
    .C(_04541_),
    .D(_06885_),
    .Y(_06888_));
 sky130_fd_sc_hd__xnor2_1 _18399_ (.A(_06284_),
    .B(_06888_),
    .Y(_00700_));
 sky130_fd_sc_hd__o21ai_0 _18400_ (.A1(_04541_),
    .A2(_06887_),
    .B1(_04559_),
    .Y(_06889_));
 sky130_fd_sc_hd__xnor2_1 _18401_ (.A(_04681_),
    .B(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__nor2_1 _18402_ (.A(net351),
    .B(_06890_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand2_1 _18403_ (.A(_04577_),
    .B(_06284_),
    .Y(_06891_));
 sky130_fd_sc_hd__nor2_1 _18404_ (.A(_06888_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__xnor2_1 _18405_ (.A(\hash.CA1.b[21] ),
    .B(_06892_),
    .Y(_00702_));
 sky130_fd_sc_hd__o311a_4 _18406_ (.A1(_04520_),
    .A2(_04541_),
    .A3(_06886_),
    .B1(_06284_),
    .C1(_04577_),
    .X(_06893_));
 sky130_fd_sc_hd__nor2_1 _18407_ (.A(\hash.CA1.b[21] ),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__xor2_1 _18408_ (.A(\hash.CA1.b[22] ),
    .B(_06894_),
    .X(_00703_));
 sky130_fd_sc_hd__clkinv_1 _18409_ (.A(_06285_),
    .Y(_06895_));
 sky130_fd_sc_hd__o21ai_2 _18410_ (.A1(_04420_),
    .A2(\hash.CA1.b[21] ),
    .B1(_06285_),
    .Y(_06896_));
 sky130_fd_sc_hd__o31ai_1 _18411_ (.A1(_06895_),
    .A2(_06888_),
    .A3(_06891_),
    .B1(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__or3_4 _18412_ (.A(_04420_),
    .B(\hash.CA1.b[21] ),
    .C(_06892_),
    .X(_06898_));
 sky130_fd_sc_hd__nor2_1 _18413_ (.A(_06285_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__nor2_1 _18414_ (.A(_06897_),
    .B(_06899_),
    .Y(_00704_));
 sky130_fd_sc_hd__o31ai_1 _18415_ (.A1(_04420_),
    .A2(\hash.CA1.b[21] ),
    .A3(_06893_),
    .B1(_04467_),
    .Y(_06900_));
 sky130_fd_sc_hd__xnor2_1 _18416_ (.A(_04726_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__nor2_1 _18417_ (.A(net351),
    .B(_06901_),
    .Y(_00705_));
 sky130_fd_sc_hd__a21oi_1 _18418_ (.A1(_04467_),
    .A2(_06898_),
    .B1(\hash.CA1.b[24] ),
    .Y(_06902_));
 sky130_fd_sc_hd__xor2_1 _18419_ (.A(\hash.CA1.b[25] ),
    .B(_06902_),
    .X(_00706_));
 sky130_fd_sc_hd__nand2_1 _18420_ (.A(_06285_),
    .B(_06893_),
    .Y(_06903_));
 sky130_fd_sc_hd__nor2_1 _18421_ (.A(_04726_),
    .B(\hash.CA1.b[25] ),
    .Y(_06904_));
 sky130_fd_sc_hd__nand3_1 _18422_ (.A(_06896_),
    .B(_06903_),
    .C(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__xor2_1 _18423_ (.A(\hash.CA1.b[26] ),
    .B(_06905_),
    .X(_00707_));
 sky130_fd_sc_hd__a21oi_1 _18424_ (.A1(_04481_),
    .A2(_04499_),
    .B1(net351),
    .Y(_06906_));
 sky130_fd_sc_hd__o21ai_2 _18425_ (.A1(_06897_),
    .A2(_06906_),
    .B1(_04517_),
    .Y(_06907_));
 sky130_fd_sc_hd__xnor2_1 _18426_ (.A(_06288_),
    .B(_06907_),
    .Y(_00708_));
 sky130_fd_sc_hd__a31oi_1 _18427_ (.A1(_06896_),
    .A2(_06903_),
    .A3(_06904_),
    .B1(_06286_),
    .Y(_06908_));
 sky130_fd_sc_hd__or3_1 _18428_ (.A(_04537_),
    .B(_04554_),
    .C(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__o21ai_0 _18429_ (.A1(_04537_),
    .A2(_06908_),
    .B1(_04554_),
    .Y(_06910_));
 sky130_fd_sc_hd__nand3_1 _18430_ (.A(_06002_),
    .B(_06909_),
    .C(_06910_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _18431_ (.A(_06002_),
    .B(_04574_),
    .Y(\hash.CA1.b[29] ));
 sky130_fd_sc_hd__nor3b_1 _18432_ (.A(_04537_),
    .B(_04554_),
    .C_N(_06907_),
    .Y(_06911_));
 sky130_fd_sc_hd__xnor2_1 _18433_ (.A(_04754_),
    .B(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__nand2_1 _18434_ (.A(_06002_),
    .B(_06912_),
    .Y(_00710_));
 sky130_fd_sc_hd__nor4_1 _18435_ (.A(_04554_),
    .B(_04754_),
    .C(\hash.CA1.b[27] ),
    .D(_06908_),
    .Y(_06913_));
 sky130_fd_sc_hd__xnor2_1 _18436_ (.A(\hash.CA1.b[30] ),
    .B(_06913_),
    .Y(_00712_));
 sky130_fd_sc_hd__a41oi_1 _18437_ (.A1(_04662_),
    .A2(_04574_),
    .A3(_06288_),
    .A4(_06907_),
    .B1(_04588_),
    .Y(_06914_));
 sky130_fd_sc_hd__xor2_1 _18438_ (.A(_04612_),
    .B(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__nor2_1 _18439_ (.A(net352),
    .B(_06915_),
    .Y(_00713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1131 ();
 sky130_fd_sc_hd__nor2b_1 _18441_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[0] ),
    .Y(\hash.CA1.f[0] ));
 sky130_fd_sc_hd__mux2i_1 _18442_ (.A0(\hash.CA2.e_dash[0] ),
    .A1(\hash.CA2.S1.X[0] ),
    .S(_13445_),
    .Y(_06917_));
 sky130_fd_sc_hd__nor2_1 _18443_ (.A(net355),
    .B(_06917_),
    .Y(_13862_));
 sky130_fd_sc_hd__nor2b_1 _18444_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[1] ),
    .Y(\hash.CA1.f[1] ));
 sky130_fd_sc_hd__mux2i_1 _18445_ (.A0(\hash.CA2.e_dash[1] ),
    .A1(\hash.CA2.S1.X[1] ),
    .S(_12365_),
    .Y(_06918_));
 sky130_fd_sc_hd__nor2_1 _18446_ (.A(net355),
    .B(_06918_),
    .Y(_12502_));
 sky130_fd_sc_hd__xor2_2 _18447_ (.A(_12498_),
    .B(_13868_),
    .X(_12509_));
 sky130_fd_sc_hd__inv_1 _18448_ (.A(_12509_),
    .Y(_12665_));
 sky130_fd_sc_hd__xor2_1 _18449_ (.A(_12503_),
    .B(_13872_),
    .X(_12508_));
 sky130_fd_sc_hd__inv_1 _18450_ (.A(_12508_),
    .Y(_12671_));
 sky130_fd_sc_hd__a21oi_1 _18451_ (.A1(_12497_),
    .A2(_13864_),
    .B1(_13863_),
    .Y(_06919_));
 sky130_fd_sc_hd__nor2b_1 _18452_ (.A(_06919_),
    .B_N(_13868_),
    .Y(_06920_));
 sky130_fd_sc_hd__nor2_1 _18453_ (.A(_13867_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__xor2_2 _18454_ (.A(_13876_),
    .B(_06921_),
    .X(_12514_));
 sky130_fd_sc_hd__inv_1 _18455_ (.A(_13851_),
    .Y(\hash.CA1.f[3] ));
 sky130_fd_sc_hd__nor2_1 _18456_ (.A(\hash.CA2.e_dash[3] ),
    .B(\hash.CA1.S1.X[3] ),
    .Y(_06922_));
 sky130_fd_sc_hd__a21oi_1 _18457_ (.A1(_13851_),
    .A2(\hash.CA1.S1.X[3] ),
    .B1(_06922_),
    .Y(_13878_));
 sky130_fd_sc_hd__a21oi_2 _18458_ (.A1(_12500_),
    .A2(_13866_),
    .B1(_13865_),
    .Y(_06923_));
 sky130_fd_sc_hd__nor2b_4 _18459_ (.A(_06923_),
    .B_N(_13872_),
    .Y(_06924_));
 sky130_fd_sc_hd__nor2_1 _18460_ (.A(_13871_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__xor2_2 _18461_ (.A(_13880_),
    .B(_06925_),
    .X(_12513_));
 sky130_fd_sc_hd__inv_2 _18462_ (.A(_13885_),
    .Y(_06926_));
 sky130_fd_sc_hd__a21o_1 _18463_ (.A1(_12498_),
    .A2(_13868_),
    .B1(_13867_),
    .X(_06927_));
 sky130_fd_sc_hd__a21oi_2 _18464_ (.A1(_13876_),
    .A2(_06927_),
    .B1(_13875_),
    .Y(_06928_));
 sky130_fd_sc_hd__xnor2_2 _18465_ (.A(_06926_),
    .B(_06928_),
    .Y(_12519_));
 sky130_fd_sc_hd__clkinv_1 _18466_ (.A(_13889_),
    .Y(_06929_));
 sky130_fd_sc_hd__a21o_1 _18467_ (.A1(_12503_),
    .A2(_13872_),
    .B1(_13871_),
    .X(_06930_));
 sky130_fd_sc_hd__a21oi_2 _18468_ (.A1(_06930_),
    .A2(_13880_),
    .B1(_13879_),
    .Y(_06931_));
 sky130_fd_sc_hd__xnor2_1 _18469_ (.A(_06929_),
    .B(_06931_),
    .Y(_12518_));
 sky130_fd_sc_hd__a21oi_1 _18470_ (.A1(_13880_),
    .A2(_13871_),
    .B1(_13879_),
    .Y(_06932_));
 sky130_fd_sc_hd__nor2_2 _18471_ (.A(_06929_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__a311oi_1 _18472_ (.A1(_13880_),
    .A2(_13889_),
    .A3(_06924_),
    .B1(_06933_),
    .C1(_13888_),
    .Y(_06934_));
 sky130_fd_sc_hd__xnor2_1 _18473_ (.A(_13899_),
    .B(_06934_),
    .Y(_12523_));
 sky130_fd_sc_hd__inv_1 _18474_ (.A(_12523_),
    .Y(_12688_));
 sky130_fd_sc_hd__o21bai_1 _18475_ (.A1(_06926_),
    .A2(_06928_),
    .B1_N(_13884_),
    .Y(_06935_));
 sky130_fd_sc_hd__a21oi_2 _18476_ (.A1(_13895_),
    .A2(_06935_),
    .B1(_13894_),
    .Y(_06936_));
 sky130_fd_sc_hd__xnor2_1 _18477_ (.A(_13904_),
    .B(_06936_),
    .Y(_12529_));
 sky130_fd_sc_hd__inv_1 _18478_ (.A(_12529_),
    .Y(_12691_));
 sky130_fd_sc_hd__mux2_8 _18479_ (.A0(\hash.CA2.e_dash[6] ),
    .A1(\hash.CA1.f[6] ),
    .S(\hash.CA1.S1.X[6] ),
    .X(_13906_));
 sky130_fd_sc_hd__o21bai_1 _18480_ (.A1(_06929_),
    .A2(_06931_),
    .B1_N(_13888_),
    .Y(_06937_));
 sky130_fd_sc_hd__a21oi_2 _18481_ (.A1(_06937_),
    .A2(_13899_),
    .B1(_13898_),
    .Y(_06938_));
 sky130_fd_sc_hd__xnor2_1 _18482_ (.A(_13908_),
    .B(_06938_),
    .Y(_12528_));
 sky130_fd_sc_hd__inv_1 _18483_ (.A(_12528_),
    .Y(_12697_));
 sky130_fd_sc_hd__o21ai_2 _18484_ (.A1(_13895_),
    .A2(_13894_),
    .B1(_13904_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand2b_4 _18485_ (.A_N(_13903_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__a21o_1 _18486_ (.A1(_13876_),
    .A2(_13867_),
    .B1(_13875_),
    .X(_06941_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_13885_),
    .B(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__nand4b_1 _18488_ (.A_N(_06919_),
    .B(_13885_),
    .C(_13876_),
    .D(_13868_),
    .Y(_06943_));
 sky130_fd_sc_hd__nor3_1 _18489_ (.A(_13884_),
    .B(_13894_),
    .C(_13903_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand3_2 _18490_ (.A(_06942_),
    .B(_06943_),
    .C(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__and2_4 _18491_ (.A(_06940_),
    .B(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__xor2_1 _18492_ (.A(_13912_),
    .B(_06946_),
    .X(_12534_));
 sky130_fd_sc_hd__inv_1 _18493_ (.A(_12534_),
    .Y(_12700_));
 sky130_fd_sc_hd__inv_1 _18494_ (.A(_13908_),
    .Y(_06947_));
 sky130_fd_sc_hd__nor2_1 _18495_ (.A(_13899_),
    .B(_13898_),
    .Y(_06948_));
 sky130_fd_sc_hd__nor2_1 _18496_ (.A(_06947_),
    .B(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__nor2_2 _18497_ (.A(_13907_),
    .B(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__or3_4 _18498_ (.A(_13888_),
    .B(_13898_),
    .C(_13907_),
    .X(_06951_));
 sky130_fd_sc_hd__a311oi_2 _18499_ (.A1(_13880_),
    .A2(_13889_),
    .A3(_06924_),
    .B1(_06933_),
    .C1(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__or2_4 _18500_ (.A(_06950_),
    .B(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__xnor2_1 _18501_ (.A(_13916_),
    .B(_06953_),
    .Y(_12533_));
 sky130_fd_sc_hd__inv_1 _18502_ (.A(_12533_),
    .Y(_12705_));
 sky130_fd_sc_hd__clkinv_2 _18503_ (.A(_13920_),
    .Y(_06954_));
 sky130_fd_sc_hd__clkinv_1 _18504_ (.A(_13904_),
    .Y(_06955_));
 sky130_fd_sc_hd__o21bai_4 _18505_ (.A1(_06955_),
    .A2(_06936_),
    .B1_N(_13903_),
    .Y(_06956_));
 sky130_fd_sc_hd__a21oi_1 _18506_ (.A1(_13912_),
    .A2(_06956_),
    .B1(_13911_),
    .Y(_06957_));
 sky130_fd_sc_hd__xnor2_1 _18507_ (.A(_06954_),
    .B(_06957_),
    .Y(_12539_));
 sky130_fd_sc_hd__o21bai_2 _18508_ (.A1(_06947_),
    .A2(_06938_),
    .B1_N(_13907_),
    .Y(_06958_));
 sky130_fd_sc_hd__a21oi_4 _18509_ (.A1(_06958_),
    .A2(_13916_),
    .B1(_13915_),
    .Y(_06959_));
 sky130_fd_sc_hd__xor2_2 _18510_ (.A(_13924_),
    .B(_06959_),
    .X(_12538_));
 sky130_fd_sc_hd__a21oi_1 _18511_ (.A1(_13912_),
    .A2(_06946_),
    .B1(_13911_),
    .Y(_06960_));
 sky130_fd_sc_hd__o21bai_2 _18512_ (.A1(_06954_),
    .A2(_06960_),
    .B1_N(_13919_),
    .Y(_06961_));
 sky130_fd_sc_hd__xor2_2 _18513_ (.A(_13929_),
    .B(_06961_),
    .X(_12544_));
 sky130_fd_sc_hd__inv_1 _18514_ (.A(_12544_),
    .Y(_12713_));
 sky130_fd_sc_hd__nor2_1 _18515_ (.A(_06954_),
    .B(_06957_),
    .Y(_06962_));
 sky130_fd_sc_hd__o21ai_0 _18516_ (.A1(_13919_),
    .A2(_06962_),
    .B1(_13929_),
    .Y(_06963_));
 sky130_fd_sc_hd__nand2b_2 _18517_ (.A_N(_13928_),
    .B(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__xnor2_2 _18518_ (.A(_13938_),
    .B(_06964_),
    .Y(_12549_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1130 ();
 sky130_fd_sc_hd__nand2_1 _18520_ (.A(_13924_),
    .B(_13933_),
    .Y(_06966_));
 sky130_fd_sc_hd__a21oi_1 _18521_ (.A1(_13933_),
    .A2(_13923_),
    .B1(_13932_),
    .Y(_06967_));
 sky130_fd_sc_hd__o21ai_2 _18522_ (.A1(_06959_),
    .A2(_06966_),
    .B1(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__xor2_2 _18523_ (.A(_13942_),
    .B(_06968_),
    .X(_12728_));
 sky130_fd_sc_hd__inv_1 _18524_ (.A(_12728_),
    .Y(_12548_));
 sky130_fd_sc_hd__inv_4 _18525_ (.A(_13947_),
    .Y(_06969_));
 sky130_fd_sc_hd__nand4_1 _18526_ (.A(_13912_),
    .B(_13920_),
    .C(_13929_),
    .D(_13938_),
    .Y(_06970_));
 sky130_fd_sc_hd__inv_1 _18527_ (.A(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__a21o_1 _18528_ (.A1(_13920_),
    .A2(_13911_),
    .B1(_13919_),
    .X(_06972_));
 sky130_fd_sc_hd__a21o_1 _18529_ (.A1(_13929_),
    .A2(_06972_),
    .B1(_13928_),
    .X(_06973_));
 sky130_fd_sc_hd__a21o_4 _18530_ (.A1(_13938_),
    .A2(_06973_),
    .B1(_13937_),
    .X(_06974_));
 sky130_fd_sc_hd__a21o_1 _18531_ (.A1(_06946_),
    .A2(_06971_),
    .B1(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__xnor2_1 _18532_ (.A(_06969_),
    .B(_06975_),
    .Y(_12731_));
 sky130_fd_sc_hd__inv_1 _18533_ (.A(_12731_),
    .Y(_12554_));
 sky130_fd_sc_hd__nor3_2 _18534_ (.A(net351),
    .B(\hash.CA2.e_dash[11] ),
    .C(_06575_),
    .Y(_06976_));
 sky130_fd_sc_hd__a21oi_4 _18535_ (.A1(_06453_),
    .A2(_06575_),
    .B1(_06976_),
    .Y(_13949_));
 sky130_fd_sc_hd__nand4_1 _18536_ (.A(_13924_),
    .B(_13916_),
    .C(_13933_),
    .D(_13942_),
    .Y(_06977_));
 sky130_fd_sc_hd__a21o_1 _18537_ (.A1(_13924_),
    .A2(_13915_),
    .B1(_13923_),
    .X(_06978_));
 sky130_fd_sc_hd__a21o_1 _18538_ (.A1(_13933_),
    .A2(_06978_),
    .B1(_13932_),
    .X(_06979_));
 sky130_fd_sc_hd__a21oi_2 _18539_ (.A1(_13942_),
    .A2(_06979_),
    .B1(_13941_),
    .Y(_06980_));
 sky130_fd_sc_hd__o31ai_4 _18540_ (.A1(net1048),
    .A2(_06977_),
    .A3(_06950_),
    .B1(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__xor2_2 _18541_ (.A(_06981_),
    .B(_13951_),
    .X(_12737_));
 sky130_fd_sc_hd__inv_1 _18542_ (.A(_12737_),
    .Y(_12553_));
 sky130_fd_sc_hd__clkinvlp_4 _18543_ (.A(_13957_),
    .Y(_06982_));
 sky130_fd_sc_hd__nor2_1 _18544_ (.A(_06969_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__nor3_1 _18545_ (.A(_06969_),
    .B(_06982_),
    .C(_06970_),
    .Y(_06984_));
 sky130_fd_sc_hd__a222oi_1 _18546_ (.A1(_13957_),
    .A2(_13946_),
    .B1(_06974_),
    .B2(_06983_),
    .C1(_06984_),
    .C2(_06956_),
    .Y(_06985_));
 sky130_fd_sc_hd__nand2b_1 _18547_ (.A_N(_13956_),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__a21oi_1 _18548_ (.A1(_13966_),
    .A2(_06986_),
    .B1(_13965_),
    .Y(_06987_));
 sky130_fd_sc_hd__xor2_2 _18549_ (.A(_13974_),
    .B(_06987_),
    .X(_12569_));
 sky130_fd_sc_hd__mux2_8 _18550_ (.A0(\hash.CA1.f[14] ),
    .A1(\hash.CA2.e_dash[14] ),
    .S(_06597_),
    .X(_13976_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1129 ();
 sky130_fd_sc_hd__a21o_4 _18552_ (.A1(_13961_),
    .A2(_13950_),
    .B1(_13960_),
    .X(_06989_));
 sky130_fd_sc_hd__inv_1 _18553_ (.A(_13916_),
    .Y(_06990_));
 sky130_fd_sc_hd__nand2_2 _18554_ (.A(_13951_),
    .B(_13961_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand3_1 _18555_ (.A(_13924_),
    .B(_13933_),
    .C(_13942_),
    .Y(_06992_));
 sky130_fd_sc_hd__nor3_1 _18556_ (.A(_06990_),
    .B(_06991_),
    .C(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__nor2b_1 _18557_ (.A(_06967_),
    .B_N(_13942_),
    .Y(_06994_));
 sky130_fd_sc_hd__nor2_1 _18558_ (.A(_13941_),
    .B(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__nand3_1 _18559_ (.A(_13951_),
    .B(_13961_),
    .C(_13915_),
    .Y(_06996_));
 sky130_fd_sc_hd__o22ai_1 _18560_ (.A1(_06991_),
    .A2(_06995_),
    .B1(_06992_),
    .B2(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__a21oi_2 _18561_ (.A1(_06993_),
    .A2(_06958_),
    .B1(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__nand2b_1 _18562_ (.A_N(_06989_),
    .B(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__a21oi_2 _18563_ (.A1(_13970_),
    .A2(_06999_),
    .B1(_13969_),
    .Y(_07000_));
 sky130_fd_sc_hd__xnor2_2 _18564_ (.A(_07000_),
    .B(_13978_),
    .Y(_12756_));
 sky130_fd_sc_hd__inv_1 _18565_ (.A(_12756_),
    .Y(_12568_));
 sky130_fd_sc_hd__a311o_1 _18566_ (.A1(_06940_),
    .A2(_06945_),
    .A3(_06971_),
    .B1(_06974_),
    .C1(_13946_),
    .X(_07001_));
 sky130_fd_sc_hd__inv_1 _18567_ (.A(_13946_),
    .Y(_07002_));
 sky130_fd_sc_hd__a21oi_2 _18568_ (.A1(_06969_),
    .A2(_07002_),
    .B1(_06982_),
    .Y(_07003_));
 sky130_fd_sc_hd__nor3_2 _18569_ (.A(_13956_),
    .B(_13965_),
    .C(_13973_),
    .Y(_07004_));
 sky130_fd_sc_hd__a21boi_4 _18570_ (.A1(_07001_),
    .A2(_07003_),
    .B1_N(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__or2_4 _18571_ (.A(_13966_),
    .B(_13965_),
    .X(_07006_));
 sky130_fd_sc_hd__a21oi_4 _18572_ (.A1(_13974_),
    .A2(_07006_),
    .B1(_13973_),
    .Y(_07007_));
 sky130_fd_sc_hd__nor2_4 _18573_ (.A(_07005_),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__xnor2_2 _18574_ (.A(_13983_),
    .B(_07008_),
    .Y(_12574_));
 sky130_fd_sc_hd__o21a_4 _18575_ (.A1(_06953_),
    .A2(_06977_),
    .B1(_06980_),
    .X(_07009_));
 sky130_fd_sc_hd__nand3_1 _18576_ (.A(_13951_),
    .B(_13961_),
    .C(_13970_),
    .Y(_07010_));
 sky130_fd_sc_hd__nand2_1 _18577_ (.A(_13970_),
    .B(_06989_),
    .Y(_07011_));
 sky130_fd_sc_hd__o21a_1 _18578_ (.A1(_07009_),
    .A2(_07010_),
    .B1(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__nand2b_1 _18579_ (.A_N(_13969_),
    .B(_07012_),
    .Y(_07013_));
 sky130_fd_sc_hd__a21oi_2 _18580_ (.A1(_13978_),
    .A2(_07013_),
    .B1(_13977_),
    .Y(_07014_));
 sky130_fd_sc_hd__xnor2_2 _18581_ (.A(_07014_),
    .B(_13987_),
    .Y(_12764_));
 sky130_fd_sc_hd__inv_1 _18582_ (.A(_12764_),
    .Y(_12573_));
 sky130_fd_sc_hd__nor3_4 _18583_ (.A(net351),
    .B(\hash.CA2.e_dash[16] ),
    .C(\hash.CA1.S1.X[16] ),
    .Y(_07015_));
 sky130_fd_sc_hd__a21oi_4 _18584_ (.A1(_06462_),
    .A2(\hash.CA1.S1.X[16] ),
    .B1(_07015_),
    .Y(_13995_));
 sky130_fd_sc_hd__inv_6 _18585_ (.A(_06568_),
    .Y(\hash.CA1.S1.X[10] ));
 sky130_fd_sc_hd__mux2_1 _18586_ (.A0(_06467_),
    .A1(\hash.CA2.e_dash[18] ),
    .S(_06634_),
    .X(_14012_));
 sky130_fd_sc_hd__and4_4 _18587_ (.A(_13983_),
    .B(_13993_),
    .C(_14002_),
    .D(_14010_),
    .X(_07016_));
 sky130_fd_sc_hd__nand3_1 _18588_ (.A(_14018_),
    .B(_14026_),
    .C(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__a211oi_2 _18589_ (.A1(_06985_),
    .A2(_07004_),
    .B1(_07007_),
    .C1(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__a21o_1 _18590_ (.A1(_13993_),
    .A2(_13982_),
    .B1(_13992_),
    .X(_07019_));
 sky130_fd_sc_hd__a21o_1 _18591_ (.A1(_14002_),
    .A2(_07019_),
    .B1(_14001_),
    .X(_07020_));
 sky130_fd_sc_hd__a21o_4 _18592_ (.A1(_14010_),
    .A2(_07020_),
    .B1(_14009_),
    .X(_07021_));
 sky130_fd_sc_hd__a21oi_1 _18593_ (.A1(_14018_),
    .A2(_07021_),
    .B1(_14017_),
    .Y(_07022_));
 sky130_fd_sc_hd__nor2b_4 _18594_ (.A(_07022_),
    .B_N(_14026_),
    .Y(_07023_));
 sky130_fd_sc_hd__a21oi_2 _18595_ (.A1(_06985_),
    .A2(_07004_),
    .B1(_07007_),
    .Y(_07024_));
 sky130_fd_sc_hd__and2_0 _18596_ (.A(_07024_),
    .B(_07016_),
    .X(_07025_));
 sky130_fd_sc_hd__o21ai_0 _18597_ (.A1(_07025_),
    .A2(_07021_),
    .B1(_14018_),
    .Y(_07026_));
 sky130_fd_sc_hd__nor3b_2 _18598_ (.A(_14026_),
    .B(_14017_),
    .C_N(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__nor3_4 _18599_ (.A(_07018_),
    .B(_07023_),
    .C(_07027_),
    .Y(_12599_));
 sky130_fd_sc_hd__inv_1 _18600_ (.A(_12599_),
    .Y(_12792_));
 sky130_fd_sc_hd__a21o_1 _18601_ (.A1(_14026_),
    .A2(_14017_),
    .B1(_14025_),
    .X(_07028_));
 sky130_fd_sc_hd__nand2_1 _18602_ (.A(_14018_),
    .B(_14026_),
    .Y(_07029_));
 sky130_fd_sc_hd__a21oi_2 _18603_ (.A1(_07008_),
    .A2(_07016_),
    .B1(_07021_),
    .Y(_07030_));
 sky130_fd_sc_hd__nor2_1 _18604_ (.A(_07029_),
    .B(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__nor2_1 _18605_ (.A(_07028_),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__xnor2_2 _18606_ (.A(_14034_),
    .B(_07032_),
    .Y(_12801_));
 sky130_fd_sc_hd__inv_1 _18607_ (.A(_12801_),
    .Y(_12604_));
 sky130_fd_sc_hd__nand2_4 _18608_ (.A(_13997_),
    .B(_14006_),
    .Y(_07033_));
 sky130_fd_sc_hd__nand2_1 _18609_ (.A(_13978_),
    .B(_13987_),
    .Y(_07034_));
 sky130_fd_sc_hd__nor2_1 _18610_ (.A(_07010_),
    .B(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__a21o_1 _18611_ (.A1(_13978_),
    .A2(_13969_),
    .B1(_13977_),
    .X(_07036_));
 sky130_fd_sc_hd__a21oi_1 _18612_ (.A1(_13987_),
    .A2(_07036_),
    .B1(_13986_),
    .Y(_07037_));
 sky130_fd_sc_hd__o21ai_0 _18613_ (.A1(_07011_),
    .A2(_07034_),
    .B1(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__a21oi_2 _18614_ (.A1(_06981_),
    .A2(_07035_),
    .B1(_07038_),
    .Y(_07039_));
 sky130_fd_sc_hd__nand2_4 _18615_ (.A(_14006_),
    .B(_13996_),
    .Y(_07040_));
 sky130_fd_sc_hd__o21ai_4 _18616_ (.A1(_07033_),
    .A2(_07039_),
    .B1(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__and3_4 _18617_ (.A(_14014_),
    .B(_14022_),
    .C(_14030_),
    .X(_07042_));
 sky130_fd_sc_hd__a21o_1 _18618_ (.A1(_14014_),
    .A2(_14005_),
    .B1(_14013_),
    .X(_07043_));
 sky130_fd_sc_hd__a21o_1 _18619_ (.A1(_14022_),
    .A2(_07043_),
    .B1(_14021_),
    .X(_07044_));
 sky130_fd_sc_hd__a21o_1 _18620_ (.A1(_14030_),
    .A2(_07044_),
    .B1(_14029_),
    .X(_07045_));
 sky130_fd_sc_hd__a21o_1 _18621_ (.A1(_07041_),
    .A2(_07042_),
    .B1(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__xor2_1 _18622_ (.A(_14038_),
    .B(_07046_),
    .X(_12807_));
 sky130_fd_sc_hd__clkinv_1 _18623_ (.A(_12807_),
    .Y(_12603_));
 sky130_fd_sc_hd__o31ai_1 _18624_ (.A1(_14025_),
    .A2(_07018_),
    .A3(_07023_),
    .B1(_14034_),
    .Y(_07047_));
 sky130_fd_sc_hd__nor2_1 _18625_ (.A(_14043_),
    .B(_14033_),
    .Y(_07048_));
 sky130_fd_sc_hd__o21a_1 _18626_ (.A1(_14034_),
    .A2(_14033_),
    .B1(_14043_),
    .X(_07049_));
 sky130_fd_sc_hd__o41a_1 _18627_ (.A1(_14025_),
    .A2(_14033_),
    .A3(_07018_),
    .A4(_07023_),
    .B1(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__a21o_4 _18628_ (.A1(_07047_),
    .A2(_07048_),
    .B1(_07050_),
    .X(_12609_));
 sky130_fd_sc_hd__nor3_1 _18629_ (.A(_13969_),
    .B(_13977_),
    .C(_06989_),
    .Y(_07051_));
 sky130_fd_sc_hd__or2_0 _18630_ (.A(_13970_),
    .B(_13969_),
    .X(_07052_));
 sky130_fd_sc_hd__a21oi_1 _18631_ (.A1(_13978_),
    .A2(_07052_),
    .B1(_13977_),
    .Y(_07053_));
 sky130_fd_sc_hd__a21oi_2 _18632_ (.A1(_06998_),
    .A2(_07051_),
    .B1(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__a21oi_4 _18633_ (.A1(_13987_),
    .A2(_07054_),
    .B1(_13986_),
    .Y(_07055_));
 sky130_fd_sc_hd__o21ai_4 _18634_ (.A1(_07033_),
    .A2(_07055_),
    .B1(_07040_),
    .Y(_07056_));
 sky130_fd_sc_hd__a21o_1 _18635_ (.A1(_14038_),
    .A2(_07045_),
    .B1(_14037_),
    .X(_07057_));
 sky130_fd_sc_hd__a31o_1 _18636_ (.A1(_14038_),
    .A2(_07042_),
    .A3(_07056_),
    .B1(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__xor2_1 _18637_ (.A(_14047_),
    .B(_07058_),
    .X(_12814_));
 sky130_fd_sc_hd__inv_1 _18638_ (.A(_12814_),
    .Y(_12608_));
 sky130_fd_sc_hd__and3_1 _18639_ (.A(_14018_),
    .B(_14026_),
    .C(_14034_),
    .X(_07059_));
 sky130_fd_sc_hd__nand3_1 _18640_ (.A(_14043_),
    .B(_07016_),
    .C(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_1 _18641_ (.A(_07021_),
    .B(_07059_),
    .Y(_07061_));
 sky130_fd_sc_hd__a21oi_1 _18642_ (.A1(_14034_),
    .A2(_07028_),
    .B1(_14033_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21bo_1 _18643_ (.A1(_07061_),
    .A2(_07062_),
    .B1_N(_14043_),
    .X(_07063_));
 sky130_fd_sc_hd__inv_1 _18644_ (.A(_14042_),
    .Y(_07064_));
 sky130_fd_sc_hd__o311ai_2 _18645_ (.A1(_07005_),
    .A2(_07007_),
    .A3(_07060_),
    .B1(_07063_),
    .C1(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__xor2_2 _18646_ (.A(_14053_),
    .B(_07065_),
    .X(_12817_));
 sky130_fd_sc_hd__inv_1 _18647_ (.A(_12817_),
    .Y(_12614_));
 sky130_fd_sc_hd__nand3_2 _18648_ (.A(_14038_),
    .B(_14047_),
    .C(_07042_),
    .Y(_07066_));
 sky130_fd_sc_hd__nor2b_1 _18649_ (.A(_07066_),
    .B_N(_07041_),
    .Y(_07067_));
 sky130_fd_sc_hd__a21oi_2 _18650_ (.A1(_14047_),
    .A2(_07057_),
    .B1(_14046_),
    .Y(_07068_));
 sky130_fd_sc_hd__nor2b_1 _18651_ (.A(_07067_),
    .B_N(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__xnor2_1 _18652_ (.A(_14057_),
    .B(_07069_),
    .Y(_12823_));
 sky130_fd_sc_hd__clkinv_1 _18653_ (.A(_12823_),
    .Y(_12613_));
 sky130_fd_sc_hd__o21ai_0 _18654_ (.A1(_14042_),
    .A2(_07050_),
    .B1(_14053_),
    .Y(_07070_));
 sky130_fd_sc_hd__nand2b_2 _18655_ (.A_N(_14052_),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__xnor2_2 _18656_ (.A(_14063_),
    .B(_07071_),
    .Y(_12619_));
 sky130_fd_sc_hd__mux2_1 _18657_ (.A0(_06487_),
    .A1(\hash.CA2.e_dash[24] ),
    .S(_06673_),
    .X(_14065_));
 sky130_fd_sc_hd__inv_1 _18658_ (.A(_07056_),
    .Y(_07072_));
 sky130_fd_sc_hd__o21ai_0 _18659_ (.A1(_07072_),
    .A2(_07066_),
    .B1(_07068_),
    .Y(_07073_));
 sky130_fd_sc_hd__a21oi_1 _18660_ (.A1(_14057_),
    .A2(_07073_),
    .B1(_14056_),
    .Y(_07074_));
 sky130_fd_sc_hd__xnor2_1 _18661_ (.A(_14067_),
    .B(_07074_),
    .Y(_12830_));
 sky130_fd_sc_hd__inv_1 _18662_ (.A(_12830_),
    .Y(_12618_));
 sky130_fd_sc_hd__a21o_1 _18663_ (.A1(_14053_),
    .A2(_07065_),
    .B1(_14052_),
    .X(_07075_));
 sky130_fd_sc_hd__a21o_4 _18664_ (.A1(_14063_),
    .A2(_07075_),
    .B1(_14062_),
    .X(_07076_));
 sky130_fd_sc_hd__xor2_2 _18665_ (.A(_14073_),
    .B(_07076_),
    .X(_12833_));
 sky130_fd_sc_hd__inv_1 _18666_ (.A(_12833_),
    .Y(_12624_));
 sky130_fd_sc_hd__nor3_2 _18667_ (.A(net354),
    .B(\hash.CA2.e_dash[25] ),
    .C(_06683_),
    .Y(_07077_));
 sky130_fd_sc_hd__a21oi_4 _18668_ (.A1(_06490_),
    .A2(_06683_),
    .B1(_07077_),
    .Y(_14075_));
 sky130_fd_sc_hd__clkinv_1 _18669_ (.A(_14077_),
    .Y(_07078_));
 sky130_fd_sc_hd__nand2_2 _18670_ (.A(_14067_),
    .B(_14057_),
    .Y(_07079_));
 sky130_fd_sc_hd__nor2_2 _18671_ (.A(_07066_),
    .B(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__nand2_1 _18672_ (.A(_14067_),
    .B(_14056_),
    .Y(_07081_));
 sky130_fd_sc_hd__o21ai_2 _18673_ (.A1(_07068_),
    .A2(_07079_),
    .B1(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__a211o_4 _18674_ (.A1(_07041_),
    .A2(_07080_),
    .B1(_07082_),
    .C1(_14066_),
    .X(_07083_));
 sky130_fd_sc_hd__xnor2_1 _18675_ (.A(_07078_),
    .B(_07083_),
    .Y(_12839_));
 sky130_fd_sc_hd__clkinv_1 _18676_ (.A(_12839_),
    .Y(_12623_));
 sky130_fd_sc_hd__nand2_2 _18677_ (.A(_14073_),
    .B(_07076_),
    .Y(_07084_));
 sky130_fd_sc_hd__nand2b_1 _18678_ (.A_N(_14072_),
    .B(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__a21o_1 _18679_ (.A1(_14083_),
    .A2(_07085_),
    .B1(_14082_),
    .X(_07086_));
 sky130_fd_sc_hd__xor2_2 _18680_ (.A(_14092_),
    .B(_07086_),
    .X(_12848_));
 sky130_fd_sc_hd__inv_1 _18681_ (.A(_12848_),
    .Y(_12634_));
 sky130_fd_sc_hd__nor3_1 _18682_ (.A(net354),
    .B(\hash.CA2.e_dash[27] ),
    .C(_06699_),
    .Y(_07087_));
 sky130_fd_sc_hd__a21oi_4 _18683_ (.A1(_06497_),
    .A2(_06699_),
    .B1(_07087_),
    .Y(_14094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1128 ();
 sky130_fd_sc_hd__a21o_1 _18685_ (.A1(_14077_),
    .A2(_07083_),
    .B1(_14076_),
    .X(_07089_));
 sky130_fd_sc_hd__a21oi_1 _18686_ (.A1(_14087_),
    .A2(_07089_),
    .B1(_14086_),
    .Y(_07090_));
 sky130_fd_sc_hd__xnor2_1 _18687_ (.A(_14096_),
    .B(_07090_),
    .Y(_12853_));
 sky130_fd_sc_hd__inv_1 _18688_ (.A(_12853_),
    .Y(_12633_));
 sky130_fd_sc_hd__o211ai_1 _18689_ (.A1(_14042_),
    .A2(_07050_),
    .B1(_14053_),
    .C1(_14063_),
    .Y(_07091_));
 sky130_fd_sc_hd__a21oi_1 _18690_ (.A1(_14063_),
    .A2(_14052_),
    .B1(_14062_),
    .Y(_07092_));
 sky130_fd_sc_hd__a21boi_2 _18691_ (.A1(_07091_),
    .A2(_07092_),
    .B1_N(_14073_),
    .Y(_07093_));
 sky130_fd_sc_hd__o21ai_2 _18692_ (.A1(_14083_),
    .A2(_14082_),
    .B1(_14092_),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2b_4 _18693_ (.A_N(_14091_),
    .B(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__o41ai_4 _18694_ (.A1(_14072_),
    .A2(_14082_),
    .A3(_14091_),
    .A4(_07093_),
    .B1(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__xnor2_1 _18695_ (.A(_14101_),
    .B(_07096_),
    .Y(_12856_));
 sky130_fd_sc_hd__inv_1 _18696_ (.A(_12856_),
    .Y(_12639_));
 sky130_fd_sc_hd__nor2_2 _18697_ (.A(\hash.CA2.e_dash[28] ),
    .B(_06707_),
    .Y(_07097_));
 sky130_fd_sc_hd__a31oi_4 _18698_ (.A1(_06002_),
    .A2(_06501_),
    .A3(_06707_),
    .B1(_07097_),
    .Y(_14103_));
 sky130_fd_sc_hd__a211oi_2 _18699_ (.A1(_07056_),
    .A2(_07080_),
    .B1(_07082_),
    .C1(_14066_),
    .Y(_07098_));
 sky130_fd_sc_hd__nand2_1 _18700_ (.A(_14077_),
    .B(_14087_),
    .Y(_07099_));
 sky130_fd_sc_hd__a21oi_1 _18701_ (.A1(_14087_),
    .A2(_14076_),
    .B1(_14086_),
    .Y(_07100_));
 sky130_fd_sc_hd__o21ai_0 _18702_ (.A1(_07098_),
    .A2(_07099_),
    .B1(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__a21o_1 _18703_ (.A1(_14096_),
    .A2(_07101_),
    .B1(_14095_),
    .X(_07102_));
 sky130_fd_sc_hd__xor2_1 _18704_ (.A(_14105_),
    .B(_07102_),
    .X(_12861_));
 sky130_fd_sc_hd__inv_1 _18705_ (.A(_12861_),
    .Y(_12638_));
 sky130_fd_sc_hd__nand2_1 _18706_ (.A(_14101_),
    .B(_14111_),
    .Y(_07103_));
 sky130_fd_sc_hd__inv_1 _18707_ (.A(_14101_),
    .Y(_07104_));
 sky130_fd_sc_hd__nor3b_1 _18708_ (.A(_14100_),
    .B(_14110_),
    .C_N(_14120_),
    .Y(_07105_));
 sky130_fd_sc_hd__o21ai_0 _18709_ (.A1(_07104_),
    .A2(_07096_),
    .B1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__o31ai_1 _18710_ (.A1(_14120_),
    .A2(_07096_),
    .A3(_07103_),
    .B1(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__a21oi_1 _18711_ (.A1(_14111_),
    .A2(_14100_),
    .B1(_14110_),
    .Y(_07108_));
 sky130_fd_sc_hd__nor2_1 _18712_ (.A(_14120_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__nor3b_1 _18713_ (.A(_14111_),
    .B(_14110_),
    .C_N(_14120_),
    .Y(_07110_));
 sky130_fd_sc_hd__nor3_2 _18714_ (.A(_07107_),
    .B(_07109_),
    .C(_07110_),
    .Y(_12649_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1127 ();
 sky130_fd_sc_hd__nand4_1 _18716_ (.A(_14096_),
    .B(_14105_),
    .C(_14115_),
    .D(_07101_),
    .Y(_07112_));
 sky130_fd_sc_hd__nand2_1 _18717_ (.A(_14115_),
    .B(_14104_),
    .Y(_07113_));
 sky130_fd_sc_hd__nand3_1 _18718_ (.A(_14105_),
    .B(_14115_),
    .C(_14095_),
    .Y(_07114_));
 sky130_fd_sc_hd__nand4b_1 _18719_ (.A_N(_14114_),
    .B(_07112_),
    .C(_07113_),
    .D(_07114_),
    .Y(_07115_));
 sky130_fd_sc_hd__xnor2_1 _18720_ (.A(_14124_),
    .B(_07115_),
    .Y(_12648_));
 sky130_fd_sc_hd__o21bai_1 _18721_ (.A1(_06990_),
    .A2(_06953_),
    .B1_N(_13915_),
    .Y(_07116_));
 sky130_fd_sc_hd__a21oi_2 _18722_ (.A1(_13924_),
    .A2(_07116_),
    .B1(_13923_),
    .Y(_07117_));
 sky130_fd_sc_hd__xnor2_2 _18723_ (.A(_13933_),
    .B(_07117_),
    .Y(_12720_));
 sky130_fd_sc_hd__o21ai_0 _18724_ (.A1(_06959_),
    .A2(_06992_),
    .B1(_06995_),
    .Y(_07118_));
 sky130_fd_sc_hd__a21oi_2 _18725_ (.A1(_13951_),
    .A2(_07118_),
    .B1(_13950_),
    .Y(_07119_));
 sky130_fd_sc_hd__xnor2_1 _18726_ (.A(_13961_),
    .B(_07119_),
    .Y(_12743_));
 sky130_fd_sc_hd__nor2_1 _18727_ (.A(_07009_),
    .B(_06991_),
    .Y(_07120_));
 sky130_fd_sc_hd__o31a_1 _18728_ (.A1(_13970_),
    .A2(_06989_),
    .A3(_07120_),
    .B1(_07012_),
    .X(_12749_));
 sky130_fd_sc_hd__xnor2_1 _18729_ (.A(_13997_),
    .B(_07055_),
    .Y(_12771_));
 sky130_fd_sc_hd__nor2_1 _18730_ (.A(_14006_),
    .B(_13996_),
    .Y(_07121_));
 sky130_fd_sc_hd__nand2b_1 _18731_ (.A_N(_07039_),
    .B(_13997_),
    .Y(_07122_));
 sky130_fd_sc_hd__a21oi_1 _18732_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07041_),
    .Y(_12777_));
 sky130_fd_sc_hd__nor2_2 _18733_ (.A(_14005_),
    .B(_07056_),
    .Y(_07123_));
 sky130_fd_sc_hd__xnor2_1 _18734_ (.A(_14014_),
    .B(_07123_),
    .Y(_12783_));
 sky130_fd_sc_hd__o21a_1 _18735_ (.A1(_14005_),
    .A2(_07041_),
    .B1(_14014_),
    .X(_07124_));
 sky130_fd_sc_hd__nor2_2 _18736_ (.A(_14013_),
    .B(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__xnor2_1 _18737_ (.A(_14022_),
    .B(_07125_),
    .Y(_12789_));
 sky130_fd_sc_hd__o21ai_0 _18738_ (.A1(_14005_),
    .A2(_07056_),
    .B1(_14014_),
    .Y(_07126_));
 sky130_fd_sc_hd__nand2b_1 _18739_ (.A_N(_14013_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21oi_2 _18740_ (.A1(_14022_),
    .A2(_07127_),
    .B1(_14021_),
    .Y(_07128_));
 sky130_fd_sc_hd__xnor2_1 _18741_ (.A(_14030_),
    .B(_07128_),
    .Y(_12798_));
 sky130_fd_sc_hd__o21bai_2 _18742_ (.A1(_07078_),
    .A2(_07098_),
    .B1_N(_14076_),
    .Y(_07129_));
 sky130_fd_sc_hd__xor2_1 _18743_ (.A(_14087_),
    .B(_07129_),
    .X(_12845_));
 sky130_fd_sc_hd__a2111o_1 _18744_ (.A1(_14077_),
    .A2(_07083_),
    .B1(_14095_),
    .C1(_14086_),
    .D1(_14076_),
    .X(_07130_));
 sky130_fd_sc_hd__nor3_1 _18745_ (.A(_14087_),
    .B(_14086_),
    .C(_14095_),
    .Y(_07131_));
 sky130_fd_sc_hd__nor2_1 _18746_ (.A(_14096_),
    .B(_14095_),
    .Y(_07132_));
 sky130_fd_sc_hd__nor2_1 _18747_ (.A(_07131_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__a31oi_4 _18748_ (.A1(_14105_),
    .A2(_07130_),
    .A3(_07133_),
    .B1(_14104_),
    .Y(_07134_));
 sky130_fd_sc_hd__xnor2_1 _18749_ (.A(_14115_),
    .B(_07134_),
    .Y(_12867_));
 sky130_fd_sc_hd__clkinvlp_4 _18750_ (.A(net1041),
    .Y(_00906_));
 sky130_fd_sc_hd__inv_1 _18751_ (.A(_12988_),
    .Y(_11600_));
 sky130_fd_sc_hd__inv_1 _18752_ (.A(_13111_),
    .Y(_11848_));
 sky130_fd_sc_hd__inv_2 _18753_ (.A(_13231_),
    .Y(_12083_));
 sky130_fd_sc_hd__inv_1 _18754_ (.A(_13240_),
    .Y(_12105_));
 sky130_fd_sc_hd__inv_1 _18755_ (.A(\hash.CA1.k_i2[1] ),
    .Y(_12366_));
 sky130_fd_sc_hd__inv_1 _18756_ (.A(\hash.CA1.k_i2[0] ),
    .Y(_12371_));
 sky130_fd_sc_hd__inv_1 _18757_ (.A(\hash.CA1.k_i2[3] ),
    .Y(_12381_));
 sky130_fd_sc_hd__inv_1 _18758_ (.A(\hash.CA1.k_i2[5] ),
    .Y(_12389_));
 sky130_fd_sc_hd__inv_1 _18759_ (.A(\hash.CA1.k_i2[7] ),
    .Y(_12397_));
 sky130_fd_sc_hd__clkinv_2 _18760_ (.A(\hash.CA1.k_i2[8] ),
    .Y(_12402_));
 sky130_fd_sc_hd__inv_1 _18761_ (.A(\hash.CA1.k_i2[11] ),
    .Y(_12413_));
 sky130_fd_sc_hd__inv_1 _18762_ (.A(\hash.CA1.k_i2[12] ),
    .Y(_12418_));
 sky130_fd_sc_hd__inv_1 _18763_ (.A(\hash.CA1.k_i2[14] ),
    .Y(_12426_));
 sky130_fd_sc_hd__inv_1 _18764_ (.A(\hash.CA1.k_i2[15] ),
    .Y(_12431_));
 sky130_fd_sc_hd__inv_1 _18765_ (.A(\hash.CA1.k_i2[16] ),
    .Y(_12436_));
 sky130_fd_sc_hd__inv_1 _18766_ (.A(\hash.CA1.k_i2[17] ),
    .Y(_12441_));
 sky130_fd_sc_hd__inv_1 _18767_ (.A(\hash.CA1.k_i2[23] ),
    .Y(_12461_));
 sky130_fd_sc_hd__inv_1 _18768_ (.A(\hash.CA1.k_i2[24] ),
    .Y(_12466_));
 sky130_fd_sc_hd__inv_1 _18769_ (.A(\hash.CA1.k_i2[25] ),
    .Y(_12471_));
 sky130_fd_sc_hd__inv_1 _18770_ (.A(\hash.CA1.k_i2[26] ),
    .Y(_12476_));
 sky130_fd_sc_hd__inv_1 _18771_ (.A(\hash.CA1.k_i2[27] ),
    .Y(_12481_));
 sky130_fd_sc_hd__clkinv_1 _18772_ (.A(\hash.CA1.k_i2[28] ),
    .Y(_12486_));
 sky130_fd_sc_hd__inv_1 _18773_ (.A(_12724_),
    .Y(_12736_));
 sky130_fd_sc_hd__inv_2 _18774_ (.A(_14204_),
    .Y(_12879_));
 sky130_fd_sc_hd__inv_1 _18775_ (.A(_14207_),
    .Y(_12884_));
 sky130_fd_sc_hd__inv_1 _18776_ (.A(_14208_),
    .Y(_12889_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1123 ();
 sky130_fd_sc_hd__mux4_2 _18781_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1119 ();
 sky130_fd_sc_hd__mux4_2 _18786_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1117 ();
 sky130_fd_sc_hd__mux4_2 _18789_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1114 ();
 sky130_fd_sc_hd__mux4_2 _18793_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1110 ();
 sky130_fd_sc_hd__mux4_2 _18798_ (.A0(_07139_),
    .A1(_07144_),
    .A2(_07147_),
    .A3(_07151_),
    .S0(net403),
    .S1(net401),
    .X(_07156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1108 ();
 sky130_fd_sc_hd__mux4_2 _18801_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1106 ();
 sky130_fd_sc_hd__mux4_2 _18804_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07162_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1104 ();
 sky130_fd_sc_hd__mux4_2 _18807_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1102 ();
 sky130_fd_sc_hd__mux4_2 _18810_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net409),
    .S1(net416),
    .X(_07168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1100 ();
 sky130_fd_sc_hd__mux4_2 _18813_ (.A0(_07159_),
    .A1(_07162_),
    .A2(_07165_),
    .A3(_07168_),
    .S0(net403),
    .S1(net401),
    .X(_07171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1099 ();
 sky130_fd_sc_hd__mux2i_4 _18815_ (.A0(_07156_),
    .A1(_07171_),
    .S(net400),
    .Y(_11580_));
 sky130_fd_sc_hd__mux4_2 _18816_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net408),
    .S1(net414),
    .X(_07173_));
 sky130_fd_sc_hd__mux4_2 _18817_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net408),
    .S1(net414),
    .X(_07174_));
 sky130_fd_sc_hd__mux4_2 _18818_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net408),
    .S1(net414),
    .X(_07175_));
 sky130_fd_sc_hd__mux4_2 _18819_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net408),
    .S1(net414),
    .X(_07176_));
 sky130_fd_sc_hd__mux4_2 _18820_ (.A0(_07173_),
    .A1(_07174_),
    .A2(_07175_),
    .A3(_07176_),
    .S0(net403),
    .S1(net401),
    .X(_07177_));
 sky130_fd_sc_hd__mux4_2 _18821_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net409),
    .S1(net416),
    .X(_07178_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1098 ();
 sky130_fd_sc_hd__mux4_2 _18823_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net409),
    .S1(net416),
    .X(_07180_));
 sky130_fd_sc_hd__mux4_2 _18824_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net409),
    .S1(net416),
    .X(_07181_));
 sky130_fd_sc_hd__mux4_2 _18825_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net409),
    .S1(net416),
    .X(_07182_));
 sky130_fd_sc_hd__mux4_2 _18826_ (.A0(_07178_),
    .A1(_07180_),
    .A2(_07181_),
    .A3(_07182_),
    .S0(net403),
    .S1(net401),
    .X(_07183_));
 sky130_fd_sc_hd__mux2i_4 _18827_ (.A0(_07177_),
    .A1(_07183_),
    .S(net400),
    .Y(_11585_));
 sky130_fd_sc_hd__mux4_2 _18828_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net409),
    .S1(net416),
    .X(_07184_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1097 ();
 sky130_fd_sc_hd__mux4_2 _18830_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net409),
    .S1(net416),
    .X(_07186_));
 sky130_fd_sc_hd__mux4_2 _18831_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net409),
    .S1(net416),
    .X(_07187_));
 sky130_fd_sc_hd__mux4_2 _18832_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net409),
    .S1(net416),
    .X(_07188_));
 sky130_fd_sc_hd__mux4_2 _18833_ (.A0(_07184_),
    .A1(_07186_),
    .A2(_07187_),
    .A3(_07188_),
    .S0(net403),
    .S1(net401),
    .X(_07189_));
 sky130_fd_sc_hd__mux4_2 _18834_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net407),
    .S1(net413),
    .X(_07190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1096 ();
 sky130_fd_sc_hd__mux4_2 _18836_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net407),
    .S1(net413),
    .X(_07192_));
 sky130_fd_sc_hd__mux4_2 _18837_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net407),
    .S1(net413),
    .X(_07193_));
 sky130_fd_sc_hd__mux4_2 _18838_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net407),
    .S1(net413),
    .X(_07194_));
 sky130_fd_sc_hd__mux4_2 _18839_ (.A0(_07190_),
    .A1(_07192_),
    .A2(_07193_),
    .A3(_07194_),
    .S0(net404),
    .S1(net401),
    .X(_07195_));
 sky130_fd_sc_hd__mux2i_4 _18840_ (.A0(_07189_),
    .A1(_07195_),
    .S(net399),
    .Y(_11593_));
 sky130_fd_sc_hd__mux4_2 _18841_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07196_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1095 ();
 sky130_fd_sc_hd__mux4_2 _18843_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07198_));
 sky130_fd_sc_hd__mux4_2 _18844_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07199_));
 sky130_fd_sc_hd__mux4_2 _18845_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07200_));
 sky130_fd_sc_hd__mux4_2 _18846_ (.A0(_07196_),
    .A1(_07198_),
    .A2(_07199_),
    .A3(_07200_),
    .S0(net403),
    .S1(net402),
    .X(_07201_));
 sky130_fd_sc_hd__mux4_2 _18847_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07202_));
 sky130_fd_sc_hd__mux4_2 _18848_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1094 ();
 sky130_fd_sc_hd__mux4_2 _18850_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07205_));
 sky130_fd_sc_hd__mux4_2 _18851_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net408),
    .S1(net414),
    .X(_07206_));
 sky130_fd_sc_hd__mux4_2 _18852_ (.A0(_07202_),
    .A1(_07203_),
    .A2(_07205_),
    .A3(_07206_),
    .S0(net403),
    .S1(net402),
    .X(_07207_));
 sky130_fd_sc_hd__mux2i_4 _18853_ (.A0(_07201_),
    .A1(_07207_),
    .S(net400),
    .Y(_11604_));
 sky130_fd_sc_hd__mux4_2 _18854_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net409),
    .S1(net416),
    .X(_07208_));
 sky130_fd_sc_hd__mux4_2 _18855_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net409),
    .S1(net416),
    .X(_07209_));
 sky130_fd_sc_hd__mux4_2 _18856_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net409),
    .S1(net416),
    .X(_07210_));
 sky130_fd_sc_hd__mux4_2 _18857_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net409),
    .S1(net416),
    .X(_07211_));
 sky130_fd_sc_hd__mux4_2 _18858_ (.A0(_07208_),
    .A1(_07209_),
    .A2(_07210_),
    .A3(_07211_),
    .S0(net403),
    .S1(net401),
    .X(_07212_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1093 ();
 sky130_fd_sc_hd__mux4_2 _18860_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net407),
    .S1(net413),
    .X(_07214_));
 sky130_fd_sc_hd__mux4_2 _18861_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net407),
    .S1(net416),
    .X(_07215_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1092 ();
 sky130_fd_sc_hd__mux4_2 _18863_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net407),
    .S1(net413),
    .X(_07217_));
 sky130_fd_sc_hd__mux4_2 _18864_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net407),
    .S1(net416),
    .X(_07218_));
 sky130_fd_sc_hd__mux4_2 _18865_ (.A0(_07214_),
    .A1(_07215_),
    .A2(_07217_),
    .A3(_07218_),
    .S0(net404),
    .S1(net401),
    .X(_07219_));
 sky130_fd_sc_hd__mux2i_4 _18866_ (.A0(_07212_),
    .A1(_07219_),
    .S(net399),
    .Y(_11612_));
 sky130_fd_sc_hd__mux4_2 _18867_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07220_));
 sky130_fd_sc_hd__mux4_2 _18868_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07221_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1091 ();
 sky130_fd_sc_hd__mux4_2 _18870_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07223_));
 sky130_fd_sc_hd__mux4_2 _18871_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07224_));
 sky130_fd_sc_hd__mux4_2 _18872_ (.A0(_07220_),
    .A1(_07221_),
    .A2(_07223_),
    .A3(_07224_),
    .S0(net403),
    .S1(net402),
    .X(_07225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1090 ();
 sky130_fd_sc_hd__mux4_2 _18874_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07227_));
 sky130_fd_sc_hd__mux4_2 _18875_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07228_));
 sky130_fd_sc_hd__mux4_2 _18876_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07229_));
 sky130_fd_sc_hd__mux4_2 _18877_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net408),
    .S1(net414),
    .X(_07230_));
 sky130_fd_sc_hd__mux4_2 _18878_ (.A0(_07227_),
    .A1(_07228_),
    .A2(_07229_),
    .A3(_07230_),
    .S0(net403),
    .S1(net402),
    .X(_07231_));
 sky130_fd_sc_hd__mux2i_4 _18879_ (.A0(_07225_),
    .A1(_07231_),
    .S(net400),
    .Y(_11620_));
 sky130_fd_sc_hd__mux4_2 _18880_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net412),
    .S1(net547),
    .X(_07232_));
 sky130_fd_sc_hd__mux4_2 _18881_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net412),
    .S1(net547),
    .X(_07233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1089 ();
 sky130_fd_sc_hd__mux4_2 _18883_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net412),
    .S1(net547),
    .X(_07235_));
 sky130_fd_sc_hd__mux4_2 _18884_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net412),
    .S1(net547),
    .X(_07236_));
 sky130_fd_sc_hd__mux4_2 _18885_ (.A0(_07232_),
    .A1(_07233_),
    .A2(_07235_),
    .A3(_07236_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07237_));
 sky130_fd_sc_hd__mux4_2 _18886_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(\count7_1[2] ),
    .S1(net417),
    .X(_07238_));
 sky130_fd_sc_hd__mux4_2 _18887_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(\count7_1[2] ),
    .S1(net417),
    .X(_07239_));
 sky130_fd_sc_hd__mux4_2 _18888_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net405),
    .S1(net417),
    .X(_07240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1088 ();
 sky130_fd_sc_hd__mux4_2 _18890_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(\count7_1[2] ),
    .S1(net417),
    .X(_07242_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1087 ();
 sky130_fd_sc_hd__mux4_2 _18892_ (.A0(_07238_),
    .A1(_07239_),
    .A2(_07240_),
    .A3(_07242_),
    .S0(net546),
    .S1(net545),
    .X(_07244_));
 sky130_fd_sc_hd__mux2i_2 _18893_ (.A0(_07237_),
    .A1(_07244_),
    .S(net400),
    .Y(_11628_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1086 ();
 sky130_fd_sc_hd__mux4_2 _18895_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net412),
    .S1(net547),
    .X(_07246_));
 sky130_fd_sc_hd__mux4_2 _18896_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net412),
    .S1(net547),
    .X(_07247_));
 sky130_fd_sc_hd__mux4_2 _18897_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net412),
    .S1(net547),
    .X(_07248_));
 sky130_fd_sc_hd__mux4_2 _18898_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net412),
    .S1(net547),
    .X(_07249_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1085 ();
 sky130_fd_sc_hd__mux4_2 _18900_ (.A0(_07246_),
    .A1(_07247_),
    .A2(_07248_),
    .A3(_07249_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07251_));
 sky130_fd_sc_hd__mux4_2 _18901_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(\count7_1[2] ),
    .S1(net417),
    .X(_07252_));
 sky130_fd_sc_hd__mux4_2 _18902_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(\count7_1[2] ),
    .S1(net417),
    .X(_07253_));
 sky130_fd_sc_hd__mux4_2 _18903_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(\count7_1[2] ),
    .S1(net417),
    .X(_07254_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1084 ();
 sky130_fd_sc_hd__mux4_2 _18905_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(\count7_1[2] ),
    .S1(net417),
    .X(_07256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1083 ();
 sky130_fd_sc_hd__mux4_2 _18907_ (.A0(_07252_),
    .A1(_07253_),
    .A2(_07254_),
    .A3(_07256_),
    .S0(net546),
    .S1(net401),
    .X(_07258_));
 sky130_fd_sc_hd__mux2i_4 _18908_ (.A0(_07251_),
    .A1(_07258_),
    .S(net400),
    .Y(_11636_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1082 ();
 sky130_fd_sc_hd__mux4_2 _18910_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net406),
    .S1(net413),
    .X(_07260_));
 sky130_fd_sc_hd__mux4_2 _18911_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net406),
    .S1(net413),
    .X(_07261_));
 sky130_fd_sc_hd__mux4_2 _18912_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net406),
    .S1(net413),
    .X(_07262_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1081 ();
 sky130_fd_sc_hd__mux4_2 _18914_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net406),
    .S1(net413),
    .X(_07264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1080 ();
 sky130_fd_sc_hd__mux4_2 _18916_ (.A0(_07260_),
    .A1(_07261_),
    .A2(_07262_),
    .A3(_07264_),
    .S0(net403),
    .S1(net401),
    .X(_07266_));
 sky130_fd_sc_hd__mux4_2 _18917_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net410),
    .S1(net415),
    .X(_07267_));
 sky130_fd_sc_hd__mux4_2 _18918_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net410),
    .S1(net415),
    .X(_07268_));
 sky130_fd_sc_hd__mux4_2 _18919_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net410),
    .S1(net415),
    .X(_07269_));
 sky130_fd_sc_hd__mux4_2 _18920_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net410),
    .S1(net415),
    .X(_07270_));
 sky130_fd_sc_hd__mux4_2 _18921_ (.A0(_07267_),
    .A1(_07268_),
    .A2(_07269_),
    .A3(_07270_),
    .S0(net404),
    .S1(net401),
    .X(_07271_));
 sky130_fd_sc_hd__mux2i_4 _18922_ (.A0(_07266_),
    .A1(_07271_),
    .S(net399),
    .Y(_11644_));
 sky130_fd_sc_hd__mux4_2 _18923_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07272_));
 sky130_fd_sc_hd__mux4_2 _18924_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07273_));
 sky130_fd_sc_hd__mux4_2 _18925_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07274_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1079 ();
 sky130_fd_sc_hd__mux4_2 _18927_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07276_));
 sky130_fd_sc_hd__mux4_2 _18928_ (.A0(_07272_),
    .A1(_07273_),
    .A2(_07274_),
    .A3(_07276_),
    .S0(net546),
    .S1(net545),
    .X(_07277_));
 sky130_fd_sc_hd__mux4_2 _18929_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07278_));
 sky130_fd_sc_hd__mux4_2 _18930_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07279_));
 sky130_fd_sc_hd__mux4_2 _18931_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07280_));
 sky130_fd_sc_hd__mux4_2 _18932_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net405),
    .S1(net417),
    .X(_07281_));
 sky130_fd_sc_hd__mux4_2 _18933_ (.A0(_07278_),
    .A1(_07279_),
    .A2(_07280_),
    .A3(_07281_),
    .S0(net546),
    .S1(net545),
    .X(_07282_));
 sky130_fd_sc_hd__mux2i_2 _18934_ (.A0(_07277_),
    .A1(_07282_),
    .S(net400),
    .Y(_11652_));
 sky130_fd_sc_hd__mux4_2 _18935_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net410),
    .S1(net415),
    .X(_07283_));
 sky130_fd_sc_hd__mux4_2 _18936_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net410),
    .S1(net415),
    .X(_07284_));
 sky130_fd_sc_hd__mux4_2 _18937_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net410),
    .S1(net415),
    .X(_07285_));
 sky130_fd_sc_hd__mux4_2 _18938_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net410),
    .S1(net415),
    .X(_07286_));
 sky130_fd_sc_hd__mux4_2 _18939_ (.A0(_07283_),
    .A1(_07284_),
    .A2(_07285_),
    .A3(_07286_),
    .S0(net404),
    .S1(net545),
    .X(_07287_));
 sky130_fd_sc_hd__mux4_2 _18940_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net405),
    .S1(net417),
    .X(_07288_));
 sky130_fd_sc_hd__mux4_2 _18941_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net405),
    .S1(net417),
    .X(_07289_));
 sky130_fd_sc_hd__mux4_2 _18942_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net405),
    .S1(net417),
    .X(_07290_));
 sky130_fd_sc_hd__mux4_2 _18943_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net405),
    .S1(net417),
    .X(_07291_));
 sky130_fd_sc_hd__mux4_2 _18944_ (.A0(_07288_),
    .A1(_07289_),
    .A2(_07290_),
    .A3(_07291_),
    .S0(net404),
    .S1(net545),
    .X(_07292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1078 ();
 sky130_fd_sc_hd__mux2i_4 _18946_ (.A0(_07287_),
    .A1(_07292_),
    .S(net399),
    .Y(_11660_));
 sky130_fd_sc_hd__mux4_2 _18947_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net407),
    .S1(net413),
    .X(_07294_));
 sky130_fd_sc_hd__mux4_2 _18948_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net406),
    .S1(net413),
    .X(_07295_));
 sky130_fd_sc_hd__mux4_2 _18949_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net407),
    .S1(net413),
    .X(_07296_));
 sky130_fd_sc_hd__mux4_2 _18950_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net407),
    .S1(net413),
    .X(_07297_));
 sky130_fd_sc_hd__mux4_2 _18951_ (.A0(_07294_),
    .A1(_07295_),
    .A2(_07296_),
    .A3(_07297_),
    .S0(net404),
    .S1(net545),
    .X(_07298_));
 sky130_fd_sc_hd__mux4_2 _18952_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net405),
    .S1(net417),
    .X(_07299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1077 ();
 sky130_fd_sc_hd__mux4_2 _18954_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net405),
    .S1(net417),
    .X(_07301_));
 sky130_fd_sc_hd__mux4_2 _18955_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net405),
    .S1(net417),
    .X(_07302_));
 sky130_fd_sc_hd__mux4_2 _18956_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net405),
    .S1(net417),
    .X(_07303_));
 sky130_fd_sc_hd__mux4_2 _18957_ (.A0(_07299_),
    .A1(_07301_),
    .A2(_07302_),
    .A3(_07303_),
    .S0(net546),
    .S1(net545),
    .X(_07304_));
 sky130_fd_sc_hd__mux2i_4 _18958_ (.A0(_07298_),
    .A1(_07304_),
    .S(net399),
    .Y(_11668_));
 sky130_fd_sc_hd__mux4_2 _18959_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net407),
    .S1(net413),
    .X(_07305_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1076 ();
 sky130_fd_sc_hd__mux4_2 _18961_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net407),
    .S1(net413),
    .X(_07307_));
 sky130_fd_sc_hd__mux4_2 _18962_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net407),
    .S1(net413),
    .X(_07308_));
 sky130_fd_sc_hd__mux4_2 _18963_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net407),
    .S1(net413),
    .X(_07309_));
 sky130_fd_sc_hd__mux4_2 _18964_ (.A0(_07305_),
    .A1(_07307_),
    .A2(_07308_),
    .A3(_07309_),
    .S0(net404),
    .S1(net401),
    .X(_07310_));
 sky130_fd_sc_hd__mux4_2 _18965_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net410),
    .S1(net415),
    .X(_07311_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1075 ();
 sky130_fd_sc_hd__mux4_2 _18967_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net410),
    .S1(net415),
    .X(_07313_));
 sky130_fd_sc_hd__mux4_2 _18968_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net410),
    .S1(net415),
    .X(_07314_));
 sky130_fd_sc_hd__mux4_2 _18969_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net410),
    .S1(net415),
    .X(_07315_));
 sky130_fd_sc_hd__mux4_2 _18970_ (.A0(_07311_),
    .A1(_07313_),
    .A2(_07314_),
    .A3(_07315_),
    .S0(net404),
    .S1(net401),
    .X(_07316_));
 sky130_fd_sc_hd__mux2i_4 _18971_ (.A0(_07310_),
    .A1(_07316_),
    .S(net399),
    .Y(_11676_));
 sky130_fd_sc_hd__mux4_2 _18972_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net410),
    .S1(net415),
    .X(_07317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1074 ();
 sky130_fd_sc_hd__mux4_2 _18974_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net410),
    .S1(net415),
    .X(_07319_));
 sky130_fd_sc_hd__mux4_2 _18975_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net410),
    .S1(net415),
    .X(_07320_));
 sky130_fd_sc_hd__mux4_2 _18976_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net410),
    .S1(net415),
    .X(_07321_));
 sky130_fd_sc_hd__mux4_2 _18977_ (.A0(_07317_),
    .A1(_07319_),
    .A2(_07320_),
    .A3(_07321_),
    .S0(net404),
    .S1(net545),
    .X(_07322_));
 sky130_fd_sc_hd__mux4_2 _18978_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net405),
    .S1(net417),
    .X(_07323_));
 sky130_fd_sc_hd__mux4_2 _18979_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net405),
    .S1(net417),
    .X(_07324_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1073 ();
 sky130_fd_sc_hd__mux4_2 _18981_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net405),
    .S1(net417),
    .X(_07326_));
 sky130_fd_sc_hd__mux4_2 _18982_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net405),
    .S1(net417),
    .X(_07327_));
 sky130_fd_sc_hd__mux4_2 _18983_ (.A0(_07323_),
    .A1(_07324_),
    .A2(_07326_),
    .A3(_07327_),
    .S0(net546),
    .S1(net545),
    .X(_07328_));
 sky130_fd_sc_hd__mux2i_4 _18984_ (.A0(_07322_),
    .A1(_07328_),
    .S(net399),
    .Y(_11684_));
 sky130_fd_sc_hd__mux4_2 _18985_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net406),
    .S1(net413),
    .X(_07329_));
 sky130_fd_sc_hd__mux4_2 _18986_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net406),
    .S1(net413),
    .X(_07330_));
 sky130_fd_sc_hd__mux4_2 _18987_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net406),
    .S1(net413),
    .X(_07331_));
 sky130_fd_sc_hd__mux4_2 _18988_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net406),
    .S1(net413),
    .X(_07332_));
 sky130_fd_sc_hd__mux4_2 _18989_ (.A0(_07329_),
    .A1(_07330_),
    .A2(_07331_),
    .A3(_07332_),
    .S0(net403),
    .S1(net401),
    .X(_07333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1072 ();
 sky130_fd_sc_hd__mux4_2 _18991_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net407),
    .S1(net413),
    .X(_07335_));
 sky130_fd_sc_hd__mux4_2 _18992_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net406),
    .S1(net413),
    .X(_07336_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1071 ();
 sky130_fd_sc_hd__mux4_2 _18994_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net406),
    .S1(net413),
    .X(_07338_));
 sky130_fd_sc_hd__mux4_2 _18995_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net407),
    .S1(net413),
    .X(_07339_));
 sky130_fd_sc_hd__mux4_2 _18996_ (.A0(_07335_),
    .A1(_07336_),
    .A2(_07338_),
    .A3(_07339_),
    .S0(net404),
    .S1(net401),
    .X(_07340_));
 sky130_fd_sc_hd__mux2i_4 _18997_ (.A0(_07333_),
    .A1(_07340_),
    .S(net399),
    .Y(_11692_));
 sky130_fd_sc_hd__mux4_2 _18998_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net411),
    .S1(net547),
    .X(_07341_));
 sky130_fd_sc_hd__mux4_2 _18999_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net412),
    .S1(net547),
    .X(_07342_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1070 ();
 sky130_fd_sc_hd__mux4_2 _19001_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net411),
    .S1(net547),
    .X(_07344_));
 sky130_fd_sc_hd__mux4_2 _19002_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net411),
    .S1(net547),
    .X(_07345_));
 sky130_fd_sc_hd__mux4_2 _19003_ (.A0(_07341_),
    .A1(_07342_),
    .A2(_07344_),
    .A3(_07345_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07346_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1069 ();
 sky130_fd_sc_hd__mux4_2 _19005_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net412),
    .S1(net415),
    .X(_07348_));
 sky130_fd_sc_hd__mux4_2 _19006_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net412),
    .S1(net416),
    .X(_07349_));
 sky130_fd_sc_hd__mux4_2 _19007_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net412),
    .S1(net416),
    .X(_07350_));
 sky130_fd_sc_hd__mux4_2 _19008_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net412),
    .S1(net416),
    .X(_07351_));
 sky130_fd_sc_hd__mux4_2 _19009_ (.A0(_07348_),
    .A1(_07349_),
    .A2(_07350_),
    .A3(_07351_),
    .S0(net546),
    .S1(net402),
    .X(_07352_));
 sky130_fd_sc_hd__mux2i_4 _19010_ (.A0(_07346_),
    .A1(_07352_),
    .S(net400),
    .Y(_11700_));
 sky130_fd_sc_hd__mux4_2 _19011_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net409),
    .S1(net416),
    .X(_07353_));
 sky130_fd_sc_hd__mux4_2 _19012_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net409),
    .S1(net416),
    .X(_07354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1068 ();
 sky130_fd_sc_hd__mux4_2 _19014_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net409),
    .S1(net416),
    .X(_07356_));
 sky130_fd_sc_hd__mux4_2 _19015_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net409),
    .S1(net416),
    .X(_07357_));
 sky130_fd_sc_hd__mux4_2 _19016_ (.A0(_07353_),
    .A1(_07354_),
    .A2(_07356_),
    .A3(_07357_),
    .S0(net403),
    .S1(net401),
    .X(_07358_));
 sky130_fd_sc_hd__mux4_2 _19017_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net410),
    .S1(net415),
    .X(_07359_));
 sky130_fd_sc_hd__mux4_2 _19018_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net410),
    .S1(net415),
    .X(_07360_));
 sky130_fd_sc_hd__mux4_2 _19019_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net410),
    .S1(net415),
    .X(_07361_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1067 ();
 sky130_fd_sc_hd__mux4_2 _19021_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net410),
    .S1(net415),
    .X(_07363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1066 ();
 sky130_fd_sc_hd__mux4_2 _19023_ (.A0(_07359_),
    .A1(_07360_),
    .A2(_07361_),
    .A3(_07363_),
    .S0(net404),
    .S1(net401),
    .X(_07365_));
 sky130_fd_sc_hd__mux2i_4 _19024_ (.A0(_07358_),
    .A1(_07365_),
    .S(net399),
    .Y(_11708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1065 ();
 sky130_fd_sc_hd__mux4_2 _19026_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net408),
    .S1(net414),
    .X(_07367_));
 sky130_fd_sc_hd__mux4_2 _19027_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net408),
    .S1(net414),
    .X(_07368_));
 sky130_fd_sc_hd__mux4_2 _19028_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net408),
    .S1(net414),
    .X(_07369_));
 sky130_fd_sc_hd__mux4_2 _19029_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net408),
    .S1(net414),
    .X(_07370_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1064 ();
 sky130_fd_sc_hd__mux4_2 _19031_ (.A0(_07367_),
    .A1(_07368_),
    .A2(_07369_),
    .A3(_07370_),
    .S0(net403),
    .S1(net402),
    .X(_07372_));
 sky130_fd_sc_hd__mux4_2 _19032_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net409),
    .S1(net416),
    .X(_07373_));
 sky130_fd_sc_hd__mux4_2 _19033_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net409),
    .S1(net416),
    .X(_07374_));
 sky130_fd_sc_hd__mux4_2 _19034_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net409),
    .S1(net416),
    .X(_07375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1063 ();
 sky130_fd_sc_hd__mux4_2 _19036_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net409),
    .S1(net416),
    .X(_07377_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1062 ();
 sky130_fd_sc_hd__mux4_2 _19038_ (.A0(_07373_),
    .A1(_07374_),
    .A2(_07375_),
    .A3(_07377_),
    .S0(net404),
    .S1(net401),
    .X(_07379_));
 sky130_fd_sc_hd__mux2i_4 _19039_ (.A0(_07372_),
    .A1(_07379_),
    .S(net400),
    .Y(_11716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1061 ();
 sky130_fd_sc_hd__mux4_2 _19041_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net410),
    .S1(net415),
    .X(_07381_));
 sky130_fd_sc_hd__mux4_2 _19042_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net410),
    .S1(net415),
    .X(_07382_));
 sky130_fd_sc_hd__mux4_2 _19043_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net410),
    .S1(net415),
    .X(_07383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1060 ();
 sky130_fd_sc_hd__mux4_2 _19045_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net410),
    .S1(net415),
    .X(_07385_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1059 ();
 sky130_fd_sc_hd__mux4_2 _19047_ (.A0(_07381_),
    .A1(_07382_),
    .A2(_07383_),
    .A3(_07385_),
    .S0(net404),
    .S1(net545),
    .X(_07387_));
 sky130_fd_sc_hd__mux4_2 _19048_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net407),
    .S1(net413),
    .X(_07388_));
 sky130_fd_sc_hd__mux4_2 _19049_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net407),
    .S1(net413),
    .X(_07389_));
 sky130_fd_sc_hd__mux4_2 _19050_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net407),
    .S1(net413),
    .X(_07390_));
 sky130_fd_sc_hd__mux4_2 _19051_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net407),
    .S1(net413),
    .X(_07391_));
 sky130_fd_sc_hd__mux4_2 _19052_ (.A0(_07388_),
    .A1(_07389_),
    .A2(_07390_),
    .A3(_07391_),
    .S0(net404),
    .S1(net401),
    .X(_07392_));
 sky130_fd_sc_hd__mux2i_4 _19053_ (.A0(_07387_),
    .A1(_07392_),
    .S(net399),
    .Y(_11724_));
 sky130_fd_sc_hd__mux4_2 _19054_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net406),
    .S1(net413),
    .X(_07393_));
 sky130_fd_sc_hd__mux4_2 _19055_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net406),
    .S1(net413),
    .X(_07394_));
 sky130_fd_sc_hd__mux4_2 _19056_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net406),
    .S1(net413),
    .X(_07395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1058 ();
 sky130_fd_sc_hd__mux4_2 _19058_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net406),
    .S1(net413),
    .X(_07397_));
 sky130_fd_sc_hd__mux4_2 _19059_ (.A0(_07393_),
    .A1(_07394_),
    .A2(_07395_),
    .A3(_07397_),
    .S0(net403),
    .S1(net401),
    .X(_07398_));
 sky130_fd_sc_hd__mux4_2 _19060_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net410),
    .S1(net415),
    .X(_07399_));
 sky130_fd_sc_hd__mux4_2 _19061_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net410),
    .S1(net415),
    .X(_07400_));
 sky130_fd_sc_hd__mux4_2 _19062_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net410),
    .S1(net415),
    .X(_07401_));
 sky130_fd_sc_hd__mux4_2 _19063_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net410),
    .S1(net415),
    .X(_07402_));
 sky130_fd_sc_hd__mux4_2 _19064_ (.A0(_07399_),
    .A1(_07400_),
    .A2(_07401_),
    .A3(_07402_),
    .S0(net404),
    .S1(net401),
    .X(_07403_));
 sky130_fd_sc_hd__mux2i_4 _19065_ (.A0(_07398_),
    .A1(_07403_),
    .S(net399),
    .Y(_11732_));
 sky130_fd_sc_hd__mux4_2 _19066_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07404_));
 sky130_fd_sc_hd__mux4_2 _19067_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07405_));
 sky130_fd_sc_hd__mux4_2 _19068_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07406_));
 sky130_fd_sc_hd__mux4_2 _19069_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07407_));
 sky130_fd_sc_hd__mux4_2 _19070_ (.A0(_07404_),
    .A1(_07405_),
    .A2(_07406_),
    .A3(_07407_),
    .S0(net546),
    .S1(net545),
    .X(_07408_));
 sky130_fd_sc_hd__mux4_2 _19071_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07409_));
 sky130_fd_sc_hd__mux4_2 _19072_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07410_));
 sky130_fd_sc_hd__mux4_2 _19073_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07411_));
 sky130_fd_sc_hd__mux4_2 _19074_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net405),
    .S1(net417),
    .X(_07412_));
 sky130_fd_sc_hd__mux4_2 _19075_ (.A0(_07409_),
    .A1(_07410_),
    .A2(_07411_),
    .A3(_07412_),
    .S0(net546),
    .S1(net545),
    .X(_07413_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1057 ();
 sky130_fd_sc_hd__mux2i_2 _19077_ (.A0(_07408_),
    .A1(_07413_),
    .S(net400),
    .Y(_11740_));
 sky130_fd_sc_hd__mux4_2 _19078_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07415_));
 sky130_fd_sc_hd__mux4_2 _19079_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07416_));
 sky130_fd_sc_hd__mux4_2 _19080_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07417_));
 sky130_fd_sc_hd__mux4_2 _19081_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07418_));
 sky130_fd_sc_hd__mux4_2 _19082_ (.A0(_07415_),
    .A1(_07416_),
    .A2(_07417_),
    .A3(_07418_),
    .S0(net404),
    .S1(net545),
    .X(_07419_));
 sky130_fd_sc_hd__mux4_2 _19083_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07420_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1056 ();
 sky130_fd_sc_hd__mux4_2 _19085_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07422_));
 sky130_fd_sc_hd__mux4_2 _19086_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07423_));
 sky130_fd_sc_hd__mux4_2 _19087_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net410),
    .S1(net415),
    .X(_07424_));
 sky130_fd_sc_hd__mux4_2 _19088_ (.A0(_07420_),
    .A1(_07422_),
    .A2(_07423_),
    .A3(_07424_),
    .S0(net404),
    .S1(net545),
    .X(_07425_));
 sky130_fd_sc_hd__mux2i_4 _19089_ (.A0(_07419_),
    .A1(_07425_),
    .S(net399),
    .Y(_11748_));
 sky130_fd_sc_hd__mux4_2 _19090_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net406),
    .S1(net413),
    .X(_07426_));
 sky130_fd_sc_hd__mux4_2 _19091_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net406),
    .S1(net413),
    .X(_07427_));
 sky130_fd_sc_hd__mux4_2 _19092_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net406),
    .S1(net413),
    .X(_07428_));
 sky130_fd_sc_hd__mux4_2 _19093_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net406),
    .S1(net413),
    .X(_07429_));
 sky130_fd_sc_hd__mux4_2 _19094_ (.A0(_07426_),
    .A1(_07427_),
    .A2(_07428_),
    .A3(_07429_),
    .S0(net404),
    .S1(net545),
    .X(_07430_));
 sky130_fd_sc_hd__mux4_2 _19095_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net407),
    .S1(net413),
    .X(_07431_));
 sky130_fd_sc_hd__mux4_2 _19096_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net407),
    .S1(net413),
    .X(_07432_));
 sky130_fd_sc_hd__mux4_2 _19097_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net407),
    .S1(net413),
    .X(_07433_));
 sky130_fd_sc_hd__mux4_2 _19098_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net407),
    .S1(net413),
    .X(_07434_));
 sky130_fd_sc_hd__mux4_2 _19099_ (.A0(_07431_),
    .A1(_07432_),
    .A2(_07433_),
    .A3(_07434_),
    .S0(net404),
    .S1(net401),
    .X(_07435_));
 sky130_fd_sc_hd__mux2i_4 _19100_ (.A0(_07430_),
    .A1(_07435_),
    .S(net399),
    .Y(_11756_));
 sky130_fd_sc_hd__mux4_2 _19101_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net411),
    .S1(net547),
    .X(_07436_));
 sky130_fd_sc_hd__mux4_2 _19102_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net411),
    .S1(net547),
    .X(_07437_));
 sky130_fd_sc_hd__mux4_2 _19103_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net411),
    .S1(net547),
    .X(_07438_));
 sky130_fd_sc_hd__mux4_2 _19104_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net411),
    .S1(net547),
    .X(_07439_));
 sky130_fd_sc_hd__mux4_2 _19105_ (.A0(_07436_),
    .A1(_07437_),
    .A2(_07438_),
    .A3(_07439_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07440_));
 sky130_fd_sc_hd__mux4_2 _19106_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net410),
    .S1(net415),
    .X(_07441_));
 sky130_fd_sc_hd__mux4_2 _19107_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net412),
    .S1(net415),
    .X(_07442_));
 sky130_fd_sc_hd__mux4_2 _19108_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net412),
    .S1(net415),
    .X(_07443_));
 sky130_fd_sc_hd__mux4_2 _19109_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net412),
    .S1(net415),
    .X(_07444_));
 sky130_fd_sc_hd__mux4_2 _19110_ (.A0(_07441_),
    .A1(_07442_),
    .A2(_07443_),
    .A3(_07444_),
    .S0(net404),
    .S1(net401),
    .X(_07445_));
 sky130_fd_sc_hd__mux2i_4 _19111_ (.A0(_07440_),
    .A1(_07445_),
    .S(net399),
    .Y(_11764_));
 sky130_fd_sc_hd__mux4_2 _19112_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net411),
    .S1(net547),
    .X(_07446_));
 sky130_fd_sc_hd__mux4_2 _19113_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net411),
    .S1(net547),
    .X(_07447_));
 sky130_fd_sc_hd__mux4_2 _19114_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net411),
    .S1(net547),
    .X(_07448_));
 sky130_fd_sc_hd__mux4_2 _19115_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net411),
    .S1(net547),
    .X(_07449_));
 sky130_fd_sc_hd__mux4_2 _19116_ (.A0(_07446_),
    .A1(_07447_),
    .A2(_07448_),
    .A3(_07449_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07450_));
 sky130_fd_sc_hd__mux4_2 _19117_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net409),
    .S1(net416),
    .X(_07451_));
 sky130_fd_sc_hd__mux4_2 _19118_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net409),
    .S1(net416),
    .X(_07452_));
 sky130_fd_sc_hd__mux4_2 _19119_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net408),
    .S1(net414),
    .X(_07453_));
 sky130_fd_sc_hd__mux4_2 _19120_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net409),
    .S1(net416),
    .X(_07454_));
 sky130_fd_sc_hd__mux4_2 _19121_ (.A0(_07451_),
    .A1(_07452_),
    .A2(_07453_),
    .A3(_07454_),
    .S0(net403),
    .S1(net402),
    .X(_07455_));
 sky130_fd_sc_hd__mux2i_4 _19122_ (.A0(_07450_),
    .A1(_07455_),
    .S(net400),
    .Y(_11772_));
 sky130_fd_sc_hd__mux4_2 _19123_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net406),
    .S1(net413),
    .X(_07456_));
 sky130_fd_sc_hd__mux4_2 _19124_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net406),
    .S1(net413),
    .X(_07457_));
 sky130_fd_sc_hd__mux4_2 _19125_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net406),
    .S1(net413),
    .X(_07458_));
 sky130_fd_sc_hd__mux4_2 _19126_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net406),
    .S1(net413),
    .X(_07459_));
 sky130_fd_sc_hd__mux4_2 _19127_ (.A0(_07456_),
    .A1(_07457_),
    .A2(_07458_),
    .A3(_07459_),
    .S0(net403),
    .S1(net401),
    .X(_07460_));
 sky130_fd_sc_hd__mux4_2 _19128_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net407),
    .S1(net413),
    .X(_07461_));
 sky130_fd_sc_hd__mux4_2 _19129_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net407),
    .S1(net413),
    .X(_07462_));
 sky130_fd_sc_hd__mux4_2 _19130_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net407),
    .S1(net413),
    .X(_07463_));
 sky130_fd_sc_hd__mux4_2 _19131_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net407),
    .S1(net413),
    .X(_07464_));
 sky130_fd_sc_hd__mux4_2 _19132_ (.A0(_07461_),
    .A1(_07462_),
    .A2(_07463_),
    .A3(_07464_),
    .S0(net404),
    .S1(net401),
    .X(_07465_));
 sky130_fd_sc_hd__mux2i_4 _19133_ (.A0(_07460_),
    .A1(_07465_),
    .S(net399),
    .Y(_11780_));
 sky130_fd_sc_hd__mux4_2 _19134_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net411),
    .S1(net547),
    .X(_07466_));
 sky130_fd_sc_hd__mux4_2 _19135_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net411),
    .S1(net547),
    .X(_07467_));
 sky130_fd_sc_hd__mux4_2 _19136_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net411),
    .S1(net547),
    .X(_07468_));
 sky130_fd_sc_hd__mux4_2 _19137_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net411),
    .S1(net547),
    .X(_07469_));
 sky130_fd_sc_hd__mux4_2 _19138_ (.A0(_07466_),
    .A1(_07467_),
    .A2(_07468_),
    .A3(_07469_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07470_));
 sky130_fd_sc_hd__mux4_2 _19139_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net412),
    .S1(net415),
    .X(_07471_));
 sky130_fd_sc_hd__mux4_2 _19140_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net412),
    .S1(net415),
    .X(_07472_));
 sky130_fd_sc_hd__mux4_2 _19141_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net412),
    .S1(net415),
    .X(_07473_));
 sky130_fd_sc_hd__mux4_2 _19142_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net412),
    .S1(net415),
    .X(_07474_));
 sky130_fd_sc_hd__mux4_2 _19143_ (.A0(_07471_),
    .A1(_07472_),
    .A2(_07473_),
    .A3(_07474_),
    .S0(net404),
    .S1(net401),
    .X(_07475_));
 sky130_fd_sc_hd__mux2i_4 _19144_ (.A0(_07470_),
    .A1(_07475_),
    .S(net400),
    .Y(_11788_));
 sky130_fd_sc_hd__mux4_2 _19145_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net408),
    .S1(net414),
    .X(_07476_));
 sky130_fd_sc_hd__mux4_2 _19146_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net408),
    .S1(net414),
    .X(_07477_));
 sky130_fd_sc_hd__mux4_2 _19147_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net408),
    .S1(net414),
    .X(_07478_));
 sky130_fd_sc_hd__mux4_2 _19148_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net408),
    .S1(net414),
    .X(_07479_));
 sky130_fd_sc_hd__mux4_2 _19149_ (.A0(_07476_),
    .A1(_07477_),
    .A2(_07478_),
    .A3(_07479_),
    .S0(net403),
    .S1(net401),
    .X(_07480_));
 sky130_fd_sc_hd__mux4_2 _19150_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net412),
    .S1(net415),
    .X(_07481_));
 sky130_fd_sc_hd__mux4_2 _19151_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net412),
    .S1(net415),
    .X(_07482_));
 sky130_fd_sc_hd__mux4_2 _19152_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net412),
    .S1(net415),
    .X(_07483_));
 sky130_fd_sc_hd__mux4_2 _19153_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net412),
    .S1(net415),
    .X(_07484_));
 sky130_fd_sc_hd__mux4_2 _19154_ (.A0(_07481_),
    .A1(_07482_),
    .A2(_07483_),
    .A3(_07484_),
    .S0(net404),
    .S1(net401),
    .X(_07485_));
 sky130_fd_sc_hd__mux2i_4 _19155_ (.A0(_07480_),
    .A1(_07485_),
    .S(net399),
    .Y(_11796_));
 sky130_fd_sc_hd__mux4_2 _19156_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net411),
    .S1(net547),
    .X(_07486_));
 sky130_fd_sc_hd__mux4_2 _19157_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net411),
    .S1(net547),
    .X(_07487_));
 sky130_fd_sc_hd__mux4_2 _19158_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net411),
    .S1(net547),
    .X(_07488_));
 sky130_fd_sc_hd__mux4_2 _19159_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net411),
    .S1(net547),
    .X(_07489_));
 sky130_fd_sc_hd__mux4_2 _19160_ (.A0(_07486_),
    .A1(_07487_),
    .A2(_07488_),
    .A3(_07489_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07490_));
 sky130_fd_sc_hd__mux4_2 _19161_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net409),
    .S1(net416),
    .X(_07491_));
 sky130_fd_sc_hd__mux4_2 _19162_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net409),
    .S1(net416),
    .X(_07492_));
 sky130_fd_sc_hd__mux4_2 _19163_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net409),
    .S1(net416),
    .X(_07493_));
 sky130_fd_sc_hd__mux4_2 _19164_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net409),
    .S1(net416),
    .X(_07494_));
 sky130_fd_sc_hd__mux4_2 _19165_ (.A0(_07491_),
    .A1(_07492_),
    .A2(_07493_),
    .A3(_07494_),
    .S0(net403),
    .S1(net402),
    .X(_07495_));
 sky130_fd_sc_hd__mux2i_4 _19166_ (.A0(_07490_),
    .A1(_07495_),
    .S(net400),
    .Y(_11804_));
 sky130_fd_sc_hd__mux4_2 _19167_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net411),
    .S1(net547),
    .X(_07496_));
 sky130_fd_sc_hd__mux4_2 _19168_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net411),
    .S1(net547),
    .X(_07497_));
 sky130_fd_sc_hd__mux4_2 _19169_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net411),
    .S1(net547),
    .X(_07498_));
 sky130_fd_sc_hd__mux4_2 _19170_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net411),
    .S1(net547),
    .X(_07499_));
 sky130_fd_sc_hd__mux4_2 _19171_ (.A0(_07496_),
    .A1(_07497_),
    .A2(_07498_),
    .A3(_07499_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07500_));
 sky130_fd_sc_hd__mux4_2 _19172_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net412),
    .S1(net416),
    .X(_07501_));
 sky130_fd_sc_hd__mux4_2 _19173_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net412),
    .S1(net416),
    .X(_07502_));
 sky130_fd_sc_hd__mux4_2 _19174_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net412),
    .S1(net416),
    .X(_07503_));
 sky130_fd_sc_hd__mux4_2 _19175_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net412),
    .S1(net416),
    .X(_07504_));
 sky130_fd_sc_hd__mux4_2 _19176_ (.A0(_07501_),
    .A1(_07502_),
    .A2(_07503_),
    .A3(_07504_),
    .S0(net403),
    .S1(net402),
    .X(_07505_));
 sky130_fd_sc_hd__mux2i_4 _19177_ (.A0(_07500_),
    .A1(_07505_),
    .S(net400),
    .Y(_11812_));
 sky130_fd_sc_hd__mux4_2 _19178_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net412),
    .S1(\count7_1[1] ),
    .X(_07506_));
 sky130_fd_sc_hd__mux4_2 _19179_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net412),
    .S1(\count7_1[1] ),
    .X(_07507_));
 sky130_fd_sc_hd__mux4_2 _19180_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net412),
    .S1(\count7_1[1] ),
    .X(_07508_));
 sky130_fd_sc_hd__mux4_2 _19181_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net412),
    .S1(\count7_1[1] ),
    .X(_07509_));
 sky130_fd_sc_hd__mux4_2 _19182_ (.A0(_07506_),
    .A1(_07507_),
    .A2(_07508_),
    .A3(_07509_),
    .S0(\count7_1[3] ),
    .S1(net402),
    .X(_07510_));
 sky130_fd_sc_hd__mux4_2 _19183_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net405),
    .S1(net417),
    .X(_07511_));
 sky130_fd_sc_hd__mux4_2 _19184_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net405),
    .S1(net417),
    .X(_07512_));
 sky130_fd_sc_hd__mux4_2 _19185_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net405),
    .S1(net417),
    .X(_07513_));
 sky130_fd_sc_hd__mux4_2 _19186_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net405),
    .S1(net417),
    .X(_07514_));
 sky130_fd_sc_hd__mux4_2 _19187_ (.A0(_07511_),
    .A1(_07512_),
    .A2(_07513_),
    .A3(_07514_),
    .S0(net546),
    .S1(net545),
    .X(_07515_));
 sky130_fd_sc_hd__mux2i_2 _19188_ (.A0(_07510_),
    .A1(_07515_),
    .S(net400),
    .Y(_11820_));
 sky130_fd_sc_hd__inv_1 _19189_ (.A(\hash.CA1.w_i2[1] ),
    .Y(_12367_));
 sky130_fd_sc_hd__inv_1 _19190_ (.A(\hash.CA1.w_i2[0] ),
    .Y(_12372_));
 sky130_fd_sc_hd__inv_2 _19191_ (.A(\hash.CA1.w_i2[3] ),
    .Y(_12382_));
 sky130_fd_sc_hd__clkinv_1 _19192_ (.A(\hash.CA1.w_i2[5] ),
    .Y(_12390_));
 sky130_fd_sc_hd__inv_2 _19193_ (.A(\hash.CA1.w_i2[7] ),
    .Y(_12398_));
 sky130_fd_sc_hd__clkinv_4 _19194_ (.A(\hash.CA1.w_i2[8] ),
    .Y(_12403_));
 sky130_fd_sc_hd__inv_2 _19195_ (.A(\hash.CA1.w_i2[11] ),
    .Y(_12414_));
 sky130_fd_sc_hd__clkinvlp_2 _19196_ (.A(\hash.CA1.w_i2[12] ),
    .Y(_12419_));
 sky130_fd_sc_hd__inv_1 _19197_ (.A(\hash.CA1.w_i2[14] ),
    .Y(_12427_));
 sky130_fd_sc_hd__clkinv_4 _19198_ (.A(\hash.CA1.w_i2[15] ),
    .Y(_12432_));
 sky130_fd_sc_hd__inv_2 _19199_ (.A(\hash.CA1.w_i2[16] ),
    .Y(_12437_));
 sky130_fd_sc_hd__clkinvlp_2 _19200_ (.A(\hash.CA1.w_i2[17] ),
    .Y(_12442_));
 sky130_fd_sc_hd__inv_1 _19201_ (.A(\hash.CA1.w_i2[23] ),
    .Y(_12462_));
 sky130_fd_sc_hd__inv_1 _19202_ (.A(\hash.CA1.w_i2[24] ),
    .Y(_12467_));
 sky130_fd_sc_hd__inv_2 _19203_ (.A(\hash.CA1.w_i2[25] ),
    .Y(_12472_));
 sky130_fd_sc_hd__clkinvlp_4 _19204_ (.A(\hash.CA1.w_i2[26] ),
    .Y(_12477_));
 sky130_fd_sc_hd__inv_1 _19205_ (.A(\hash.CA1.w_i2[27] ),
    .Y(_12482_));
 sky130_fd_sc_hd__inv_1 _19206_ (.A(\hash.CA1.w_i2[28] ),
    .Y(_12487_));
 sky130_fd_sc_hd__inv_1 _19207_ (.A(_12725_),
    .Y(_12727_));
 sky130_fd_sc_hd__clkinv_1 _19208_ (.A(_06771_),
    .Y(_12793_));
 sky130_fd_sc_hd__inv_1 _19209_ (.A(_12898_),
    .Y(_12894_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1052 ();
 sky130_fd_sc_hd__mux4_2 _19214_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07520_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1048 ();
 sky130_fd_sc_hd__mux4_2 _19219_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1046 ();
 sky130_fd_sc_hd__mux4_2 _19222_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1043 ();
 sky130_fd_sc_hd__mux4_2 _19226_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1039 ();
 sky130_fd_sc_hd__mux4_2 _19231_ (.A0(_07520_),
    .A1(_07525_),
    .A2(_07528_),
    .A3(_07532_),
    .S0(net482),
    .S1(net480),
    .X(_07537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1037 ();
 sky130_fd_sc_hd__mux4_2 _19234_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07540_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1035 ();
 sky130_fd_sc_hd__mux4_2 _19237_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07543_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1033 ();
 sky130_fd_sc_hd__mux4_2 _19240_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1031 ();
 sky130_fd_sc_hd__mux4_2 _19243_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net486),
    .S1(net492),
    .X(_07549_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1029 ();
 sky130_fd_sc_hd__mux4_2 _19246_ (.A0(_07540_),
    .A1(_07543_),
    .A2(_07546_),
    .A3(_07549_),
    .S0(net483),
    .S1(net481),
    .X(_07552_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1028 ();
 sky130_fd_sc_hd__mux2i_4 _19248_ (.A0(_07537_),
    .A1(_07552_),
    .S(net478),
    .Y(_11581_));
 sky130_fd_sc_hd__mux4_2 _19249_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net487),
    .S1(net494),
    .X(_07554_));
 sky130_fd_sc_hd__mux4_2 _19250_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net487),
    .S1(net494),
    .X(_07555_));
 sky130_fd_sc_hd__mux4_2 _19251_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net487),
    .S1(net494),
    .X(_07556_));
 sky130_fd_sc_hd__mux4_2 _19252_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net487),
    .S1(net494),
    .X(_07557_));
 sky130_fd_sc_hd__mux4_2 _19253_ (.A0(_07554_),
    .A1(_07555_),
    .A2(_07556_),
    .A3(_07557_),
    .S0(net482),
    .S1(net480),
    .X(_07558_));
 sky130_fd_sc_hd__mux4_2 _19254_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net488),
    .S1(net493),
    .X(_07559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1027 ();
 sky130_fd_sc_hd__mux4_2 _19256_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net488),
    .S1(net493),
    .X(_07561_));
 sky130_fd_sc_hd__mux4_2 _19257_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net488),
    .S1(net493),
    .X(_07562_));
 sky130_fd_sc_hd__mux4_2 _19258_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net488),
    .S1(net493),
    .X(_07563_));
 sky130_fd_sc_hd__mux4_2 _19259_ (.A0(_07559_),
    .A1(_07561_),
    .A2(_07562_),
    .A3(_07563_),
    .S0(net483),
    .S1(net481),
    .X(_07564_));
 sky130_fd_sc_hd__mux2i_4 _19260_ (.A0(_07558_),
    .A1(_07564_),
    .S(net478),
    .Y(_11586_));
 sky130_fd_sc_hd__mux4_2 _19261_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net555),
    .S1(net496),
    .X(_07565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1026 ();
 sky130_fd_sc_hd__mux4_2 _19263_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net555),
    .S1(net496),
    .X(_07567_));
 sky130_fd_sc_hd__mux4_2 _19264_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net555),
    .S1(net496),
    .X(_07568_));
 sky130_fd_sc_hd__mux4_2 _19265_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net555),
    .S1(net496),
    .X(_07569_));
 sky130_fd_sc_hd__mux4_2 _19266_ (.A0(_07565_),
    .A1(_07567_),
    .A2(_07568_),
    .A3(_07569_),
    .S0(net484),
    .S1(net554),
    .X(_07570_));
 sky130_fd_sc_hd__mux4_2 _19267_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net555),
    .S1(net495),
    .X(_07571_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1025 ();
 sky130_fd_sc_hd__mux4_2 _19269_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net555),
    .S1(net495),
    .X(_07573_));
 sky130_fd_sc_hd__mux4_2 _19270_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net555),
    .S1(net495),
    .X(_07574_));
 sky130_fd_sc_hd__mux4_2 _19271_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net555),
    .S1(net495),
    .X(_07575_));
 sky130_fd_sc_hd__mux4_2 _19272_ (.A0(_07571_),
    .A1(_07573_),
    .A2(_07574_),
    .A3(_07575_),
    .S0(net484),
    .S1(net554),
    .X(_07576_));
 sky130_fd_sc_hd__mux2i_4 _19273_ (.A0(_07570_),
    .A1(_07576_),
    .S(net479),
    .Y(_11594_));
 sky130_fd_sc_hd__mux4_2 _19274_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net490),
    .S1(net496),
    .X(_07577_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1024 ();
 sky130_fd_sc_hd__mux4_2 _19276_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net490),
    .S1(net496),
    .X(_07579_));
 sky130_fd_sc_hd__mux4_2 _19277_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net490),
    .S1(net496),
    .X(_07580_));
 sky130_fd_sc_hd__mux4_2 _19278_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net490),
    .S1(net496),
    .X(_07581_));
 sky130_fd_sc_hd__mux4_2 _19279_ (.A0(_07577_),
    .A1(_07579_),
    .A2(_07580_),
    .A3(_07581_),
    .S0(net484),
    .S1(\count16_1[4] ),
    .X(_07582_));
 sky130_fd_sc_hd__mux4_2 _19280_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net491),
    .S1(net556),
    .X(_07583_));
 sky130_fd_sc_hd__mux4_2 _19281_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net491),
    .S1(net556),
    .X(_07584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1023 ();
 sky130_fd_sc_hd__mux4_2 _19283_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net491),
    .S1(net556),
    .X(_07586_));
 sky130_fd_sc_hd__mux4_2 _19284_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net491),
    .S1(net556),
    .X(_07587_));
 sky130_fd_sc_hd__mux4_2 _19285_ (.A0(_07583_),
    .A1(_07584_),
    .A2(_07586_),
    .A3(_07587_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07588_));
 sky130_fd_sc_hd__mux2i_2 _19286_ (.A0(_07582_),
    .A1(_07588_),
    .S(\count16_1[5] ),
    .Y(_11605_));
 sky130_fd_sc_hd__mux4_2 _19287_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net490),
    .S1(net496),
    .X(_07589_));
 sky130_fd_sc_hd__mux4_2 _19288_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net490),
    .S1(net496),
    .X(_07590_));
 sky130_fd_sc_hd__mux4_2 _19289_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net490),
    .S1(net496),
    .X(_07591_));
 sky130_fd_sc_hd__mux4_2 _19290_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net490),
    .S1(net496),
    .X(_07592_));
 sky130_fd_sc_hd__mux4_2 _19291_ (.A0(_07589_),
    .A1(_07590_),
    .A2(_07591_),
    .A3(_07592_),
    .S0(net484),
    .S1(net554),
    .X(_07593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1022 ();
 sky130_fd_sc_hd__mux4_2 _19293_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net490),
    .S1(net495),
    .X(_07595_));
 sky130_fd_sc_hd__mux4_2 _19294_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net490),
    .S1(net495),
    .X(_07596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1021 ();
 sky130_fd_sc_hd__mux4_2 _19296_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net490),
    .S1(net495),
    .X(_07598_));
 sky130_fd_sc_hd__mux4_2 _19297_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net490),
    .S1(net495),
    .X(_07599_));
 sky130_fd_sc_hd__mux4_2 _19298_ (.A0(_07595_),
    .A1(_07596_),
    .A2(_07598_),
    .A3(_07599_),
    .S0(net484),
    .S1(net554),
    .X(_07600_));
 sky130_fd_sc_hd__mux2i_4 _19299_ (.A0(_07593_),
    .A1(_07600_),
    .S(net479),
    .Y(_11613_));
 sky130_fd_sc_hd__mux4_2 _19300_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net490),
    .S1(net496),
    .X(_07601_));
 sky130_fd_sc_hd__mux4_2 _19301_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net490),
    .S1(net496),
    .X(_07602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1020 ();
 sky130_fd_sc_hd__mux4_2 _19303_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net490),
    .S1(net496),
    .X(_07604_));
 sky130_fd_sc_hd__mux4_2 _19304_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net490),
    .S1(net496),
    .X(_07605_));
 sky130_fd_sc_hd__mux4_2 _19305_ (.A0(_07601_),
    .A1(_07602_),
    .A2(_07604_),
    .A3(_07605_),
    .S0(net484),
    .S1(net554),
    .X(_07606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1019 ();
 sky130_fd_sc_hd__mux4_2 _19307_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net555),
    .S1(net495),
    .X(_07608_));
 sky130_fd_sc_hd__mux4_2 _19308_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net555),
    .S1(net495),
    .X(_07609_));
 sky130_fd_sc_hd__mux4_2 _19309_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net555),
    .S1(net495),
    .X(_07610_));
 sky130_fd_sc_hd__mux4_2 _19310_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net555),
    .S1(net495),
    .X(_07611_));
 sky130_fd_sc_hd__mux4_2 _19311_ (.A0(_07608_),
    .A1(_07609_),
    .A2(_07610_),
    .A3(_07611_),
    .S0(net484),
    .S1(net554),
    .X(_07612_));
 sky130_fd_sc_hd__mux2i_4 _19312_ (.A0(_07606_),
    .A1(_07612_),
    .S(net479),
    .Y(_11621_));
 sky130_fd_sc_hd__mux4_2 _19313_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net490),
    .S1(net496),
    .X(_07613_));
 sky130_fd_sc_hd__mux4_2 _19314_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net490),
    .S1(net496),
    .X(_07614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1018 ();
 sky130_fd_sc_hd__mux4_2 _19316_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net490),
    .S1(net496),
    .X(_07616_));
 sky130_fd_sc_hd__mux4_2 _19317_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net490),
    .S1(net496),
    .X(_07617_));
 sky130_fd_sc_hd__mux4_2 _19318_ (.A0(_07613_),
    .A1(_07614_),
    .A2(_07616_),
    .A3(_07617_),
    .S0(net484),
    .S1(net554),
    .X(_07618_));
 sky130_fd_sc_hd__mux4_2 _19319_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(\count16_1[2] ),
    .S1(net556),
    .X(_07619_));
 sky130_fd_sc_hd__mux4_2 _19320_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(\count16_1[2] ),
    .S1(net556),
    .X(_07620_));
 sky130_fd_sc_hd__mux4_2 _19321_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(\count16_1[2] ),
    .S1(net556),
    .X(_07621_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1017 ();
 sky130_fd_sc_hd__mux4_2 _19323_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count16_1[2] ),
    .S1(net556),
    .X(_07623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1016 ();
 sky130_fd_sc_hd__mux4_2 _19325_ (.A0(_07619_),
    .A1(_07620_),
    .A2(_07621_),
    .A3(_07623_),
    .S0(net484),
    .S1(\count16_1[4] ),
    .X(_07625_));
 sky130_fd_sc_hd__mux2i_2 _19326_ (.A0(_07618_),
    .A1(_07625_),
    .S(\count16_1[5] ),
    .Y(_11629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1015 ();
 sky130_fd_sc_hd__mux4_2 _19328_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net491),
    .S1(net495),
    .X(_07627_));
 sky130_fd_sc_hd__mux4_2 _19329_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net491),
    .S1(net495),
    .X(_07628_));
 sky130_fd_sc_hd__mux4_2 _19330_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net491),
    .S1(net495),
    .X(_07629_));
 sky130_fd_sc_hd__mux4_2 _19331_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net491),
    .S1(net495),
    .X(_07630_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1014 ();
 sky130_fd_sc_hd__mux4_2 _19333_ (.A0(_07627_),
    .A1(_07628_),
    .A2(_07629_),
    .A3(_07630_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07632_));
 sky130_fd_sc_hd__mux4_2 _19334_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net489),
    .S1(net493),
    .X(_07633_));
 sky130_fd_sc_hd__mux4_2 _19335_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net489),
    .S1(net493),
    .X(_07634_));
 sky130_fd_sc_hd__mux4_2 _19336_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net489),
    .S1(net556),
    .X(_07635_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1013 ();
 sky130_fd_sc_hd__mux4_2 _19338_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net489),
    .S1(net556),
    .X(_07637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1012 ();
 sky130_fd_sc_hd__mux4_2 _19340_ (.A0(_07633_),
    .A1(_07634_),
    .A2(_07635_),
    .A3(_07637_),
    .S0(net483),
    .S1(net481),
    .X(_07639_));
 sky130_fd_sc_hd__mux2i_2 _19341_ (.A0(_07632_),
    .A1(_07639_),
    .S(net479),
    .Y(_11637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1011 ();
 sky130_fd_sc_hd__mux4_2 _19343_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net487),
    .S1(net492),
    .X(_07641_));
 sky130_fd_sc_hd__mux4_2 _19344_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net487),
    .S1(net492),
    .X(_07642_));
 sky130_fd_sc_hd__mux4_2 _19345_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net487),
    .S1(net492),
    .X(_07643_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1010 ();
 sky130_fd_sc_hd__mux4_2 _19347_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net487),
    .S1(net492),
    .X(_07645_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1009 ();
 sky130_fd_sc_hd__mux4_2 _19349_ (.A0(_07641_),
    .A1(_07642_),
    .A2(_07643_),
    .A3(_07645_),
    .S0(net482),
    .S1(net480),
    .X(_07647_));
 sky130_fd_sc_hd__mux4_2 _19350_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net486),
    .S1(net492),
    .X(_07648_));
 sky130_fd_sc_hd__mux4_2 _19351_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net486),
    .S1(net492),
    .X(_07649_));
 sky130_fd_sc_hd__mux4_2 _19352_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net486),
    .S1(net492),
    .X(_07650_));
 sky130_fd_sc_hd__mux4_2 _19353_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net486),
    .S1(net492),
    .X(_07651_));
 sky130_fd_sc_hd__mux4_2 _19354_ (.A0(_07648_),
    .A1(_07649_),
    .A2(_07650_),
    .A3(_07651_),
    .S0(net482),
    .S1(net480),
    .X(_07652_));
 sky130_fd_sc_hd__mux2i_4 _19355_ (.A0(_07647_),
    .A1(_07652_),
    .S(net478),
    .Y(_11645_));
 sky130_fd_sc_hd__mux4_2 _19356_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07653_));
 sky130_fd_sc_hd__mux4_2 _19357_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07654_));
 sky130_fd_sc_hd__mux4_2 _19358_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07655_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1008 ();
 sky130_fd_sc_hd__mux4_2 _19360_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07657_));
 sky130_fd_sc_hd__mux4_2 _19361_ (.A0(_07653_),
    .A1(_07654_),
    .A2(_07655_),
    .A3(_07657_),
    .S0(net482),
    .S1(net480),
    .X(_07658_));
 sky130_fd_sc_hd__mux4_2 _19362_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07659_));
 sky130_fd_sc_hd__mux4_2 _19363_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07660_));
 sky130_fd_sc_hd__mux4_2 _19364_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07661_));
 sky130_fd_sc_hd__mux4_2 _19365_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net486),
    .S1(net492),
    .X(_07662_));
 sky130_fd_sc_hd__mux4_2 _19366_ (.A0(_07659_),
    .A1(_07660_),
    .A2(_07661_),
    .A3(_07662_),
    .S0(net483),
    .S1(net481),
    .X(_07663_));
 sky130_fd_sc_hd__mux2i_4 _19367_ (.A0(_07658_),
    .A1(_07663_),
    .S(net478),
    .Y(_11653_));
 sky130_fd_sc_hd__mux4_2 _19368_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net486),
    .S1(net492),
    .X(_07664_));
 sky130_fd_sc_hd__mux4_2 _19369_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net486),
    .S1(net492),
    .X(_07665_));
 sky130_fd_sc_hd__mux4_2 _19370_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net486),
    .S1(net492),
    .X(_07666_));
 sky130_fd_sc_hd__mux4_2 _19371_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net486),
    .S1(net492),
    .X(_07667_));
 sky130_fd_sc_hd__mux4_2 _19372_ (.A0(_07664_),
    .A1(_07665_),
    .A2(_07666_),
    .A3(_07667_),
    .S0(net483),
    .S1(net481),
    .X(_07668_));
 sky130_fd_sc_hd__mux4_2 _19373_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net488),
    .S1(net493),
    .X(_07669_));
 sky130_fd_sc_hd__mux4_2 _19374_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net488),
    .S1(net493),
    .X(_07670_));
 sky130_fd_sc_hd__mux4_2 _19375_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net488),
    .S1(net493),
    .X(_07671_));
 sky130_fd_sc_hd__mux4_2 _19376_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net488),
    .S1(net493),
    .X(_07672_));
 sky130_fd_sc_hd__mux4_2 _19377_ (.A0(_07669_),
    .A1(_07670_),
    .A2(_07671_),
    .A3(_07672_),
    .S0(net483),
    .S1(net481),
    .X(_07673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1007 ();
 sky130_fd_sc_hd__mux2i_4 _19379_ (.A0(_07668_),
    .A1(_07673_),
    .S(net478),
    .Y(_11661_));
 sky130_fd_sc_hd__mux4_2 _19380_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net485),
    .S1(net494),
    .X(_07675_));
 sky130_fd_sc_hd__mux4_2 _19381_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net485),
    .S1(net494),
    .X(_07676_));
 sky130_fd_sc_hd__mux4_2 _19382_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net485),
    .S1(net494),
    .X(_07677_));
 sky130_fd_sc_hd__mux4_2 _19383_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net485),
    .S1(net494),
    .X(_07678_));
 sky130_fd_sc_hd__mux4_2 _19384_ (.A0(_07675_),
    .A1(_07676_),
    .A2(_07677_),
    .A3(_07678_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07679_));
 sky130_fd_sc_hd__mux4_2 _19385_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net488),
    .S1(net493),
    .X(_07680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1006 ();
 sky130_fd_sc_hd__mux4_2 _19387_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net488),
    .S1(net493),
    .X(_07682_));
 sky130_fd_sc_hd__mux4_2 _19388_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net488),
    .S1(net493),
    .X(_07683_));
 sky130_fd_sc_hd__mux4_2 _19389_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net488),
    .S1(net493),
    .X(_07684_));
 sky130_fd_sc_hd__mux4_2 _19390_ (.A0(_07680_),
    .A1(_07682_),
    .A2(_07683_),
    .A3(_07684_),
    .S0(net483),
    .S1(net481),
    .X(_07685_));
 sky130_fd_sc_hd__mux2i_2 _19391_ (.A0(_07679_),
    .A1(_07685_),
    .S(net479),
    .Y(_11669_));
 sky130_fd_sc_hd__mux4_2 _19392_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net485),
    .S1(net495),
    .X(_07686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1005 ();
 sky130_fd_sc_hd__mux4_2 _19394_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net485),
    .S1(net495),
    .X(_07688_));
 sky130_fd_sc_hd__mux4_2 _19395_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net485),
    .S1(net495),
    .X(_07689_));
 sky130_fd_sc_hd__mux4_2 _19396_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net485),
    .S1(net495),
    .X(_07690_));
 sky130_fd_sc_hd__mux4_2 _19397_ (.A0(_07686_),
    .A1(_07688_),
    .A2(_07689_),
    .A3(_07690_),
    .S0(net484),
    .S1(net554),
    .X(_07691_));
 sky130_fd_sc_hd__mux4_2 _19398_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net491),
    .S1(net556),
    .X(_07692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1004 ();
 sky130_fd_sc_hd__mux4_2 _19400_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net491),
    .S1(net556),
    .X(_07694_));
 sky130_fd_sc_hd__mux4_2 _19401_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net491),
    .S1(net556),
    .X(_07695_));
 sky130_fd_sc_hd__mux4_2 _19402_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net491),
    .S1(net556),
    .X(_07696_));
 sky130_fd_sc_hd__mux4_2 _19403_ (.A0(_07692_),
    .A1(_07694_),
    .A2(_07695_),
    .A3(_07696_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07697_));
 sky130_fd_sc_hd__mux2i_4 _19404_ (.A0(_07691_),
    .A1(_07697_),
    .S(net479),
    .Y(_11677_));
 sky130_fd_sc_hd__mux4_2 _19405_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net485),
    .S1(net495),
    .X(_07698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1003 ();
 sky130_fd_sc_hd__mux4_2 _19407_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net485),
    .S1(net495),
    .X(_07700_));
 sky130_fd_sc_hd__mux4_2 _19408_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net485),
    .S1(net495),
    .X(_07701_));
 sky130_fd_sc_hd__mux4_2 _19409_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net485),
    .S1(net495),
    .X(_07702_));
 sky130_fd_sc_hd__mux4_2 _19410_ (.A0(_07698_),
    .A1(_07700_),
    .A2(_07701_),
    .A3(_07702_),
    .S0(net484),
    .S1(net554),
    .X(_07703_));
 sky130_fd_sc_hd__mux4_2 _19411_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net491),
    .S1(net556),
    .X(_07704_));
 sky130_fd_sc_hd__mux4_2 _19412_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net491),
    .S1(net556),
    .X(_07705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1002 ();
 sky130_fd_sc_hd__mux4_2 _19414_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net491),
    .S1(net556),
    .X(_07707_));
 sky130_fd_sc_hd__mux4_2 _19415_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net491),
    .S1(net556),
    .X(_07708_));
 sky130_fd_sc_hd__mux4_2 _19416_ (.A0(_07704_),
    .A1(_07705_),
    .A2(_07707_),
    .A3(_07708_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07709_));
 sky130_fd_sc_hd__mux2i_4 _19417_ (.A0(_07703_),
    .A1(_07709_),
    .S(net479),
    .Y(_11685_));
 sky130_fd_sc_hd__mux4_2 _19418_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net485),
    .S1(net495),
    .X(_07710_));
 sky130_fd_sc_hd__mux4_2 _19419_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net485),
    .S1(net495),
    .X(_07711_));
 sky130_fd_sc_hd__mux4_2 _19420_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net485),
    .S1(net495),
    .X(_07712_));
 sky130_fd_sc_hd__mux4_2 _19421_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net485),
    .S1(net495),
    .X(_07713_));
 sky130_fd_sc_hd__mux4_2 _19422_ (.A0(_07710_),
    .A1(_07711_),
    .A2(_07712_),
    .A3(_07713_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1001 ();
 sky130_fd_sc_hd__mux4_2 _19424_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net489),
    .S1(net493),
    .X(_07716_));
 sky130_fd_sc_hd__mux4_2 _19425_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net489),
    .S1(net493),
    .X(_07717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1000 ();
 sky130_fd_sc_hd__mux4_2 _19427_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net489),
    .S1(net493),
    .X(_07719_));
 sky130_fd_sc_hd__mux4_2 _19428_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net489),
    .S1(net493),
    .X(_07720_));
 sky130_fd_sc_hd__mux4_2 _19429_ (.A0(_07716_),
    .A1(_07717_),
    .A2(_07719_),
    .A3(_07720_),
    .S0(net483),
    .S1(net481),
    .X(_07721_));
 sky130_fd_sc_hd__mux2i_4 _19430_ (.A0(_07714_),
    .A1(_07721_),
    .S(net478),
    .Y(_11693_));
 sky130_fd_sc_hd__mux4_2 _19431_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net555),
    .S1(net496),
    .X(_07722_));
 sky130_fd_sc_hd__mux4_2 _19432_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net555),
    .S1(net496),
    .X(_07723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_999 ();
 sky130_fd_sc_hd__mux4_2 _19434_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net555),
    .S1(net495),
    .X(_07725_));
 sky130_fd_sc_hd__mux4_2 _19435_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net555),
    .S1(net495),
    .X(_07726_));
 sky130_fd_sc_hd__mux4_2 _19436_ (.A0(_07722_),
    .A1(_07723_),
    .A2(_07725_),
    .A3(_07726_),
    .S0(net484),
    .S1(net554),
    .X(_07727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_998 ();
 sky130_fd_sc_hd__mux4_2 _19438_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net555),
    .S1(net495),
    .X(_07729_));
 sky130_fd_sc_hd__mux4_2 _19439_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net555),
    .S1(net495),
    .X(_07730_));
 sky130_fd_sc_hd__mux4_2 _19440_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net555),
    .S1(net495),
    .X(_07731_));
 sky130_fd_sc_hd__mux4_2 _19441_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net555),
    .S1(net495),
    .X(_07732_));
 sky130_fd_sc_hd__mux4_2 _19442_ (.A0(_07729_),
    .A1(_07730_),
    .A2(_07731_),
    .A3(_07732_),
    .S0(net484),
    .S1(net554),
    .X(_07733_));
 sky130_fd_sc_hd__mux2i_4 _19443_ (.A0(_07727_),
    .A1(_07733_),
    .S(net479),
    .Y(_11701_));
 sky130_fd_sc_hd__mux4_2 _19444_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net555),
    .S1(net496),
    .X(_07734_));
 sky130_fd_sc_hd__mux4_2 _19445_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net490),
    .S1(net496),
    .X(_07735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_997 ();
 sky130_fd_sc_hd__mux4_2 _19447_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net490),
    .S1(net496),
    .X(_07737_));
 sky130_fd_sc_hd__mux4_2 _19448_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net490),
    .S1(net496),
    .X(_07738_));
 sky130_fd_sc_hd__mux4_2 _19449_ (.A0(_07734_),
    .A1(_07735_),
    .A2(_07737_),
    .A3(_07738_),
    .S0(net484),
    .S1(net554),
    .X(_07739_));
 sky130_fd_sc_hd__mux4_2 _19450_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net491),
    .S1(net556),
    .X(_07740_));
 sky130_fd_sc_hd__mux4_2 _19451_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net491),
    .S1(net556),
    .X(_07741_));
 sky130_fd_sc_hd__mux4_2 _19452_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net491),
    .S1(net556),
    .X(_07742_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_996 ();
 sky130_fd_sc_hd__mux4_2 _19454_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net491),
    .S1(net556),
    .X(_07744_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_995 ();
 sky130_fd_sc_hd__mux4_2 _19456_ (.A0(_07740_),
    .A1(_07741_),
    .A2(_07742_),
    .A3(_07744_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07746_));
 sky130_fd_sc_hd__mux2i_2 _19457_ (.A0(_07739_),
    .A1(_07746_),
    .S(\count16_1[5] ),
    .Y(_11709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_994 ();
 sky130_fd_sc_hd__mux4_2 _19459_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07748_));
 sky130_fd_sc_hd__mux4_2 _19460_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07749_));
 sky130_fd_sc_hd__mux4_2 _19461_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07750_));
 sky130_fd_sc_hd__mux4_2 _19462_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07751_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_993 ();
 sky130_fd_sc_hd__mux4_2 _19464_ (.A0(_07748_),
    .A1(_07749_),
    .A2(_07750_),
    .A3(_07751_),
    .S0(net482),
    .S1(net480),
    .X(_07753_));
 sky130_fd_sc_hd__mux4_2 _19465_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07754_));
 sky130_fd_sc_hd__mux4_2 _19466_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07755_));
 sky130_fd_sc_hd__mux4_2 _19467_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07756_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_992 ();
 sky130_fd_sc_hd__mux4_2 _19469_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net489),
    .S1(net494),
    .X(_07758_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_991 ();
 sky130_fd_sc_hd__mux4_2 _19471_ (.A0(_07754_),
    .A1(_07755_),
    .A2(_07756_),
    .A3(_07758_),
    .S0(net482),
    .S1(net480),
    .X(_07760_));
 sky130_fd_sc_hd__mux2i_4 _19472_ (.A0(_07753_),
    .A1(_07760_),
    .S(net479),
    .Y(_11717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_990 ();
 sky130_fd_sc_hd__mux4_2 _19474_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07762_));
 sky130_fd_sc_hd__mux4_2 _19475_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07763_));
 sky130_fd_sc_hd__mux4_2 _19476_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07764_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_989 ();
 sky130_fd_sc_hd__mux4_2 _19478_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_988 ();
 sky130_fd_sc_hd__mux4_2 _19480_ (.A0(_07762_),
    .A1(_07763_),
    .A2(_07764_),
    .A3(_07766_),
    .S0(net483),
    .S1(net481),
    .X(_07768_));
 sky130_fd_sc_hd__mux4_2 _19481_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07769_));
 sky130_fd_sc_hd__mux4_2 _19482_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07770_));
 sky130_fd_sc_hd__mux4_2 _19483_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07771_));
 sky130_fd_sc_hd__mux4_2 _19484_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net488),
    .S1(net493),
    .X(_07772_));
 sky130_fd_sc_hd__mux4_2 _19485_ (.A0(_07769_),
    .A1(_07770_),
    .A2(_07771_),
    .A3(_07772_),
    .S0(net483),
    .S1(net481),
    .X(_07773_));
 sky130_fd_sc_hd__mux2i_2 _19486_ (.A0(_07768_),
    .A1(_07773_),
    .S(net479),
    .Y(_11725_));
 sky130_fd_sc_hd__mux4_2 _19487_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net487),
    .S1(net494),
    .X(_07774_));
 sky130_fd_sc_hd__mux4_2 _19488_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net487),
    .S1(net494),
    .X(_07775_));
 sky130_fd_sc_hd__mux4_2 _19489_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net487),
    .S1(net494),
    .X(_07776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_987 ();
 sky130_fd_sc_hd__mux4_2 _19491_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net487),
    .S1(net494),
    .X(_07778_));
 sky130_fd_sc_hd__mux4_2 _19492_ (.A0(_07774_),
    .A1(_07775_),
    .A2(_07776_),
    .A3(_07778_),
    .S0(net482),
    .S1(net480),
    .X(_07779_));
 sky130_fd_sc_hd__mux4_2 _19493_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net486),
    .S1(net492),
    .X(_07780_));
 sky130_fd_sc_hd__mux4_2 _19494_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net487),
    .S1(net492),
    .X(_07781_));
 sky130_fd_sc_hd__mux4_2 _19495_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net487),
    .S1(net492),
    .X(_07782_));
 sky130_fd_sc_hd__mux4_2 _19496_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net487),
    .S1(net492),
    .X(_07783_));
 sky130_fd_sc_hd__mux4_2 _19497_ (.A0(_07780_),
    .A1(_07781_),
    .A2(_07782_),
    .A3(_07783_),
    .S0(net483),
    .S1(net481),
    .X(_07784_));
 sky130_fd_sc_hd__mux2i_4 _19498_ (.A0(_07779_),
    .A1(_07784_),
    .S(net478),
    .Y(_11733_));
 sky130_fd_sc_hd__mux4_2 _19499_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net486),
    .S1(net492),
    .X(_07785_));
 sky130_fd_sc_hd__mux4_2 _19500_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net486),
    .S1(net492),
    .X(_07786_));
 sky130_fd_sc_hd__mux4_2 _19501_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net486),
    .S1(net492),
    .X(_07787_));
 sky130_fd_sc_hd__mux4_2 _19502_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net486),
    .S1(net492),
    .X(_07788_));
 sky130_fd_sc_hd__mux4_2 _19503_ (.A0(_07785_),
    .A1(_07786_),
    .A2(_07787_),
    .A3(_07788_),
    .S0(net483),
    .S1(net481),
    .X(_07789_));
 sky130_fd_sc_hd__mux4_2 _19504_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net488),
    .S1(net493),
    .X(_07790_));
 sky130_fd_sc_hd__mux4_2 _19505_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net488),
    .S1(net493),
    .X(_07791_));
 sky130_fd_sc_hd__mux4_2 _19506_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net488),
    .S1(net493),
    .X(_07792_));
 sky130_fd_sc_hd__mux4_2 _19507_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net488),
    .S1(net493),
    .X(_07793_));
 sky130_fd_sc_hd__mux4_2 _19508_ (.A0(_07790_),
    .A1(_07791_),
    .A2(_07792_),
    .A3(_07793_),
    .S0(net483),
    .S1(net481),
    .X(_07794_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_986 ();
 sky130_fd_sc_hd__mux2i_2 _19510_ (.A0(_07789_),
    .A1(_07794_),
    .S(net479),
    .Y(_11741_));
 sky130_fd_sc_hd__mux4_2 _19511_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net485),
    .S1(net494),
    .X(_07796_));
 sky130_fd_sc_hd__mux4_2 _19512_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net485),
    .S1(net494),
    .X(_07797_));
 sky130_fd_sc_hd__mux4_2 _19513_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net485),
    .S1(net494),
    .X(_07798_));
 sky130_fd_sc_hd__mux4_2 _19514_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net485),
    .S1(net494),
    .X(_07799_));
 sky130_fd_sc_hd__mux4_2 _19515_ (.A0(_07796_),
    .A1(_07797_),
    .A2(_07798_),
    .A3(_07799_),
    .S0(net482),
    .S1(net480),
    .X(_07800_));
 sky130_fd_sc_hd__mux4_2 _19516_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net489),
    .S1(net492),
    .X(_07801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_985 ();
 sky130_fd_sc_hd__mux4_2 _19518_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net489),
    .S1(net493),
    .X(_07803_));
 sky130_fd_sc_hd__mux4_2 _19519_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net489),
    .S1(net493),
    .X(_07804_));
 sky130_fd_sc_hd__mux4_2 _19520_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net489),
    .S1(net493),
    .X(_07805_));
 sky130_fd_sc_hd__mux4_2 _19521_ (.A0(_07801_),
    .A1(_07803_),
    .A2(_07804_),
    .A3(_07805_),
    .S0(net483),
    .S1(net481),
    .X(_07806_));
 sky130_fd_sc_hd__mux2i_4 _19522_ (.A0(_07800_),
    .A1(_07806_),
    .S(net478),
    .Y(_11749_));
 sky130_fd_sc_hd__mux4_2 _19523_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net486),
    .S1(net492),
    .X(_07807_));
 sky130_fd_sc_hd__mux4_2 _19524_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net486),
    .S1(net492),
    .X(_07808_));
 sky130_fd_sc_hd__mux4_2 _19525_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net486),
    .S1(net492),
    .X(_07809_));
 sky130_fd_sc_hd__mux4_2 _19526_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net486),
    .S1(net492),
    .X(_07810_));
 sky130_fd_sc_hd__mux4_2 _19527_ (.A0(_07807_),
    .A1(_07808_),
    .A2(_07809_),
    .A3(_07810_),
    .S0(net482),
    .S1(net480),
    .X(_07811_));
 sky130_fd_sc_hd__mux4_2 _19528_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net488),
    .S1(net493),
    .X(_07812_));
 sky130_fd_sc_hd__mux4_2 _19529_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net488),
    .S1(net493),
    .X(_07813_));
 sky130_fd_sc_hd__mux4_2 _19530_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net488),
    .S1(net493),
    .X(_07814_));
 sky130_fd_sc_hd__mux4_2 _19531_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net488),
    .S1(net493),
    .X(_07815_));
 sky130_fd_sc_hd__mux4_2 _19532_ (.A0(_07812_),
    .A1(_07813_),
    .A2(_07814_),
    .A3(_07815_),
    .S0(net483),
    .S1(net481),
    .X(_07816_));
 sky130_fd_sc_hd__mux2i_4 _19533_ (.A0(_07811_),
    .A1(_07816_),
    .S(net478),
    .Y(_11757_));
 sky130_fd_sc_hd__mux4_2 _19534_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net485),
    .S1(net495),
    .X(_07817_));
 sky130_fd_sc_hd__mux4_2 _19535_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net485),
    .S1(net495),
    .X(_07818_));
 sky130_fd_sc_hd__mux4_2 _19536_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net485),
    .S1(net495),
    .X(_07819_));
 sky130_fd_sc_hd__mux4_2 _19537_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net485),
    .S1(net495),
    .X(_07820_));
 sky130_fd_sc_hd__mux4_2 _19538_ (.A0(_07817_),
    .A1(_07818_),
    .A2(_07819_),
    .A3(_07820_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07821_));
 sky130_fd_sc_hd__mux4_2 _19539_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net491),
    .S1(net495),
    .X(_07822_));
 sky130_fd_sc_hd__mux4_2 _19540_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net491),
    .S1(net495),
    .X(_07823_));
 sky130_fd_sc_hd__mux4_2 _19541_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net491),
    .S1(net495),
    .X(_07824_));
 sky130_fd_sc_hd__mux4_2 _19542_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net491),
    .S1(net495),
    .X(_07825_));
 sky130_fd_sc_hd__mux4_2 _19543_ (.A0(_07822_),
    .A1(_07823_),
    .A2(_07824_),
    .A3(_07825_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07826_));
 sky130_fd_sc_hd__mux2i_4 _19544_ (.A0(_07821_),
    .A1(_07826_),
    .S(net479),
    .Y(_11765_));
 sky130_fd_sc_hd__mux4_2 _19545_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net487),
    .S1(net494),
    .X(_07827_));
 sky130_fd_sc_hd__mux4_2 _19546_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net487),
    .S1(net494),
    .X(_07828_));
 sky130_fd_sc_hd__mux4_2 _19547_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net487),
    .S1(net494),
    .X(_07829_));
 sky130_fd_sc_hd__mux4_2 _19548_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net487),
    .S1(net494),
    .X(_07830_));
 sky130_fd_sc_hd__mux4_2 _19549_ (.A0(_07827_),
    .A1(_07828_),
    .A2(_07829_),
    .A3(_07830_),
    .S0(net482),
    .S1(net480),
    .X(_07831_));
 sky130_fd_sc_hd__mux4_2 _19550_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net487),
    .S1(net492),
    .X(_07832_));
 sky130_fd_sc_hd__mux4_2 _19551_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net487),
    .S1(net492),
    .X(_07833_));
 sky130_fd_sc_hd__mux4_2 _19552_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net487),
    .S1(net492),
    .X(_07834_));
 sky130_fd_sc_hd__mux4_2 _19553_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net487),
    .S1(net492),
    .X(_07835_));
 sky130_fd_sc_hd__mux4_2 _19554_ (.A0(_07832_),
    .A1(_07833_),
    .A2(_07834_),
    .A3(_07835_),
    .S0(net482),
    .S1(net480),
    .X(_07836_));
 sky130_fd_sc_hd__mux2i_4 _19555_ (.A0(_07831_),
    .A1(_07836_),
    .S(net478),
    .Y(_11773_));
 sky130_fd_sc_hd__mux4_2 _19556_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07837_));
 sky130_fd_sc_hd__mux4_2 _19557_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07838_));
 sky130_fd_sc_hd__mux4_2 _19558_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07839_));
 sky130_fd_sc_hd__mux4_2 _19559_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07840_));
 sky130_fd_sc_hd__mux4_2 _19560_ (.A0(_07837_),
    .A1(_07838_),
    .A2(_07839_),
    .A3(_07840_),
    .S0(net482),
    .S1(net480),
    .X(_07841_));
 sky130_fd_sc_hd__mux4_2 _19561_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07842_));
 sky130_fd_sc_hd__mux4_2 _19562_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07843_));
 sky130_fd_sc_hd__mux4_2 _19563_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07844_));
 sky130_fd_sc_hd__mux4_2 _19564_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net489),
    .S1(net494),
    .X(_07845_));
 sky130_fd_sc_hd__mux4_2 _19565_ (.A0(_07842_),
    .A1(_07843_),
    .A2(_07844_),
    .A3(_07845_),
    .S0(net482),
    .S1(net480),
    .X(_07846_));
 sky130_fd_sc_hd__mux2i_4 _19566_ (.A0(_07841_),
    .A1(_07846_),
    .S(net478),
    .Y(_11781_));
 sky130_fd_sc_hd__mux4_2 _19567_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net487),
    .S1(net494),
    .X(_07847_));
 sky130_fd_sc_hd__mux4_2 _19568_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net487),
    .S1(net494),
    .X(_07848_));
 sky130_fd_sc_hd__mux4_2 _19569_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net487),
    .S1(net494),
    .X(_07849_));
 sky130_fd_sc_hd__mux4_2 _19570_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net487),
    .S1(net494),
    .X(_07850_));
 sky130_fd_sc_hd__mux4_2 _19571_ (.A0(_07847_),
    .A1(_07848_),
    .A2(_07849_),
    .A3(_07850_),
    .S0(net482),
    .S1(net480),
    .X(_07851_));
 sky130_fd_sc_hd__mux4_2 _19572_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net487),
    .S1(net492),
    .X(_07852_));
 sky130_fd_sc_hd__mux4_2 _19573_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net487),
    .S1(net492),
    .X(_07853_));
 sky130_fd_sc_hd__mux4_2 _19574_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net487),
    .S1(net492),
    .X(_07854_));
 sky130_fd_sc_hd__mux4_2 _19575_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net487),
    .S1(net492),
    .X(_07855_));
 sky130_fd_sc_hd__mux4_2 _19576_ (.A0(_07852_),
    .A1(_07853_),
    .A2(_07854_),
    .A3(_07855_),
    .S0(net482),
    .S1(net480),
    .X(_07856_));
 sky130_fd_sc_hd__mux2i_4 _19577_ (.A0(_07851_),
    .A1(_07856_),
    .S(net478),
    .Y(_11789_));
 sky130_fd_sc_hd__mux4_2 _19578_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07857_));
 sky130_fd_sc_hd__mux4_2 _19579_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07858_));
 sky130_fd_sc_hd__mux4_2 _19580_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07859_));
 sky130_fd_sc_hd__mux4_2 _19581_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07860_));
 sky130_fd_sc_hd__mux4_2 _19582_ (.A0(_07857_),
    .A1(_07858_),
    .A2(_07859_),
    .A3(_07860_),
    .S0(net484),
    .S1(net554),
    .X(_07861_));
 sky130_fd_sc_hd__mux4_2 _19583_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07862_));
 sky130_fd_sc_hd__mux4_2 _19584_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07863_));
 sky130_fd_sc_hd__mux4_2 _19585_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07864_));
 sky130_fd_sc_hd__mux4_2 _19586_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net485),
    .S1(net495),
    .X(_07865_));
 sky130_fd_sc_hd__mux4_2 _19587_ (.A0(_07862_),
    .A1(_07863_),
    .A2(_07864_),
    .A3(_07865_),
    .S0(net484),
    .S1(net554),
    .X(_07866_));
 sky130_fd_sc_hd__mux2i_4 _19588_ (.A0(_07861_),
    .A1(_07866_),
    .S(net479),
    .Y(_11797_));
 sky130_fd_sc_hd__mux4_2 _19589_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net485),
    .S1(net494),
    .X(_07867_));
 sky130_fd_sc_hd__mux4_2 _19590_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net485),
    .S1(net494),
    .X(_07868_));
 sky130_fd_sc_hd__mux4_2 _19591_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net485),
    .S1(net494),
    .X(_07869_));
 sky130_fd_sc_hd__mux4_2 _19592_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net485),
    .S1(net494),
    .X(_07870_));
 sky130_fd_sc_hd__mux4_2 _19593_ (.A0(_07867_),
    .A1(_07868_),
    .A2(_07869_),
    .A3(_07870_),
    .S0(\count16_1[3] ),
    .S1(net481),
    .X(_07871_));
 sky130_fd_sc_hd__mux4_2 _19594_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net488),
    .S1(net493),
    .X(_07872_));
 sky130_fd_sc_hd__mux4_2 _19595_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net489),
    .S1(net493),
    .X(_07873_));
 sky130_fd_sc_hd__mux4_2 _19596_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net489),
    .S1(net493),
    .X(_07874_));
 sky130_fd_sc_hd__mux4_2 _19597_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net489),
    .S1(net493),
    .X(_07875_));
 sky130_fd_sc_hd__mux4_2 _19598_ (.A0(_07872_),
    .A1(_07873_),
    .A2(_07874_),
    .A3(_07875_),
    .S0(net483),
    .S1(net481),
    .X(_07876_));
 sky130_fd_sc_hd__mux2i_4 _19599_ (.A0(_07871_),
    .A1(_07876_),
    .S(net478),
    .Y(_11805_));
 sky130_fd_sc_hd__mux4_2 _19600_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07877_));
 sky130_fd_sc_hd__mux4_2 _19601_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07878_));
 sky130_fd_sc_hd__mux4_2 _19602_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07879_));
 sky130_fd_sc_hd__mux4_2 _19603_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07880_));
 sky130_fd_sc_hd__mux4_2 _19604_ (.A0(_07877_),
    .A1(_07878_),
    .A2(_07879_),
    .A3(_07880_),
    .S0(net484),
    .S1(net554),
    .X(_07881_));
 sky130_fd_sc_hd__mux4_2 _19605_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07882_));
 sky130_fd_sc_hd__mux4_2 _19606_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07883_));
 sky130_fd_sc_hd__mux4_2 _19607_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07884_));
 sky130_fd_sc_hd__mux4_2 _19608_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net490),
    .S1(net496),
    .X(_07885_));
 sky130_fd_sc_hd__mux4_2 _19609_ (.A0(_07882_),
    .A1(_07883_),
    .A2(_07884_),
    .A3(_07885_),
    .S0(net484),
    .S1(net554),
    .X(_07886_));
 sky130_fd_sc_hd__mux2i_4 _19610_ (.A0(_07881_),
    .A1(_07886_),
    .S(net479),
    .Y(_11813_));
 sky130_fd_sc_hd__mux4_2 _19611_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07887_));
 sky130_fd_sc_hd__mux4_2 _19612_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07888_));
 sky130_fd_sc_hd__mux4_2 _19613_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07889_));
 sky130_fd_sc_hd__mux4_2 _19614_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07890_));
 sky130_fd_sc_hd__mux4_2 _19615_ (.A0(_07887_),
    .A1(_07888_),
    .A2(_07889_),
    .A3(_07890_),
    .S0(net484),
    .S1(net554),
    .X(_07891_));
 sky130_fd_sc_hd__mux4_2 _19616_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07892_));
 sky130_fd_sc_hd__mux4_2 _19617_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07893_));
 sky130_fd_sc_hd__mux4_2 _19618_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07894_));
 sky130_fd_sc_hd__mux4_2 _19619_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net490),
    .S1(net496),
    .X(_07895_));
 sky130_fd_sc_hd__mux4_2 _19620_ (.A0(_07892_),
    .A1(_07893_),
    .A2(_07894_),
    .A3(_07895_),
    .S0(net484),
    .S1(net554),
    .X(_07896_));
 sky130_fd_sc_hd__mux2i_4 _19621_ (.A0(_07891_),
    .A1(_07896_),
    .S(net479),
    .Y(_11821_));
 sky130_fd_sc_hd__inv_1 _19622_ (.A(_12504_),
    .Y(_12662_));
 sky130_fd_sc_hd__inv_1 _19623_ (.A(_12883_),
    .Y(\hash.CA1.p1[1] ));
 sky130_fd_sc_hd__inv_1 _19624_ (.A(_12886_),
    .Y(\hash.CA1.p2[2] ));
 sky130_fd_sc_hd__inv_1 _19625_ (.A(_12893_),
    .Y(\hash.CA1.p3[2] ));
 sky130_fd_sc_hd__inv_1 _19626_ (.A(_12897_),
    .Y(\hash.CA1.p5[1] ));
 sky130_fd_sc_hd__inv_1 _19627_ (.A(_12104_),
    .Y(_12107_));
 sky130_fd_sc_hd__inv_1 _19628_ (.A(_12512_),
    .Y(_12891_));
 sky130_fd_sc_hd__inv_1 _19629_ (.A(_12659_),
    .Y(_12661_));
 sky130_fd_sc_hd__inv_1 _19630_ (.A(_12686_),
    .Y(_12687_));
 sky130_fd_sc_hd__inv_1 _19631_ (.A(_12874_),
    .Y(_12876_));
 sky130_fd_sc_hd__inv_1 _19632_ (.A(_12094_),
    .Y(_12106_));
 sky130_fd_sc_hd__inv_1 _19633_ (.A(_12506_),
    .Y(_12890_));
 sky130_fd_sc_hd__inv_1 _19634_ (.A(_12655_),
    .Y(_12660_));
 sky130_fd_sc_hd__inv_1 _19635_ (.A(_12658_),
    .Y(_12670_));
 sky130_fd_sc_hd__inv_1 _19636_ (.A(_12685_),
    .Y(_12696_));
 sky130_fd_sc_hd__inv_1 _19637_ (.A(_12865_),
    .Y(_12875_));
 sky130_fd_sc_hd__clkinvlp_4 _19638_ (.A(\count_hash2[1] ),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_4 _19639_ (.A(\count_hash1[1] ),
    .Y(_00654_));
 sky130_fd_sc_hd__xor2_1 _19640_ (.A(_11335_),
    .B(_02699_),
    .X(_07897_));
 sky130_fd_sc_hd__xnor2_1 _19641_ (.A(_11090_),
    .B(_07897_),
    .Y(_12983_));
 sky130_fd_sc_hd__inv_1 _19642_ (.A(_11590_),
    .Y(_12990_));
 sky130_fd_sc_hd__inv_1 _19643_ (.A(_11598_),
    .Y(_12994_));
 sky130_fd_sc_hd__inv_1 _19644_ (.A(_11609_),
    .Y(_12998_));
 sky130_fd_sc_hd__inv_1 _19645_ (.A(_11617_),
    .Y(_13002_));
 sky130_fd_sc_hd__inv_1 _19646_ (.A(_11625_),
    .Y(_13006_));
 sky130_fd_sc_hd__clkinvlp_4 _19647_ (.A(_11633_),
    .Y(_13010_));
 sky130_fd_sc_hd__clkinv_1 _19648_ (.A(_11641_),
    .Y(_13014_));
 sky130_fd_sc_hd__inv_2 _19649_ (.A(_11649_),
    .Y(_13018_));
 sky130_fd_sc_hd__clkinv_1 _19650_ (.A(_11657_),
    .Y(_13022_));
 sky130_fd_sc_hd__clkinv_2 _19651_ (.A(_11665_),
    .Y(_13026_));
 sky130_fd_sc_hd__inv_1 _19652_ (.A(_11673_),
    .Y(_13030_));
 sky130_fd_sc_hd__inv_1 _19653_ (.A(_11681_),
    .Y(_13034_));
 sky130_fd_sc_hd__inv_1 _19654_ (.A(_11689_),
    .Y(_13038_));
 sky130_fd_sc_hd__inv_1 _19655_ (.A(_11697_),
    .Y(_13042_));
 sky130_fd_sc_hd__inv_1 _19656_ (.A(_11705_),
    .Y(_13046_));
 sky130_fd_sc_hd__inv_1 _19657_ (.A(_11713_),
    .Y(_13050_));
 sky130_fd_sc_hd__inv_1 _19658_ (.A(_11721_),
    .Y(_13054_));
 sky130_fd_sc_hd__inv_1 _19659_ (.A(_11729_),
    .Y(_13058_));
 sky130_fd_sc_hd__clkinv_1 _19660_ (.A(_11737_),
    .Y(_13062_));
 sky130_fd_sc_hd__inv_1 _19661_ (.A(_11745_),
    .Y(_13066_));
 sky130_fd_sc_hd__clkinv_1 _19662_ (.A(_11753_),
    .Y(_13070_));
 sky130_fd_sc_hd__inv_1 _19663_ (.A(_11761_),
    .Y(_13074_));
 sky130_fd_sc_hd__inv_1 _19664_ (.A(_11769_),
    .Y(_13078_));
 sky130_fd_sc_hd__inv_2 _19665_ (.A(_11777_),
    .Y(_13082_));
 sky130_fd_sc_hd__clkinv_1 _19666_ (.A(_11785_),
    .Y(_13086_));
 sky130_fd_sc_hd__clkinv_1 _19667_ (.A(_11793_),
    .Y(_13090_));
 sky130_fd_sc_hd__clkinv_1 _19668_ (.A(_11801_),
    .Y(_13094_));
 sky130_fd_sc_hd__clkinv_1 _19669_ (.A(_11809_),
    .Y(_13098_));
 sky130_fd_sc_hd__clkinv_1 _19670_ (.A(_11817_),
    .Y(_13102_));
 sky130_fd_sc_hd__mux4_2 _19671_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net465),
    .S1(net475),
    .X(_07898_));
 sky130_fd_sc_hd__mux4_2 _19672_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net465),
    .S1(net475),
    .X(_07899_));
 sky130_fd_sc_hd__mux4_2 _19673_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net465),
    .S1(net475),
    .X(_07900_));
 sky130_fd_sc_hd__mux4_2 _19674_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net465),
    .S1(net475),
    .X(_07901_));
 sky130_fd_sc_hd__mux4_2 _19675_ (.A0(_07898_),
    .A1(_07899_),
    .A2(_07900_),
    .A3(_07901_),
    .S0(net462),
    .S1(net460),
    .X(_07902_));
 sky130_fd_sc_hd__mux4_2 _19676_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net465),
    .S1(net476),
    .X(_07903_));
 sky130_fd_sc_hd__mux4_2 _19677_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net465),
    .S1(net476),
    .X(_07904_));
 sky130_fd_sc_hd__mux4_2 _19678_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net465),
    .S1(net476),
    .X(_07905_));
 sky130_fd_sc_hd__mux4_2 _19679_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net465),
    .S1(net476),
    .X(_07906_));
 sky130_fd_sc_hd__mux4_2 _19680_ (.A0(_07903_),
    .A1(_07904_),
    .A2(_07905_),
    .A3(_07906_),
    .S0(net462),
    .S1(net460),
    .X(_07907_));
 sky130_fd_sc_hd__mux2_8 _19681_ (.A0(_07902_),
    .A1(_07907_),
    .S(net458),
    .X(_13106_));
 sky130_fd_sc_hd__inv_1 _19682_ (.A(_11838_),
    .Y(_13113_));
 sky130_fd_sc_hd__inv_1 _19683_ (.A(_11846_),
    .Y(_13117_));
 sky130_fd_sc_hd__inv_1 _19684_ (.A(_11857_),
    .Y(_13121_));
 sky130_fd_sc_hd__inv_1 _19685_ (.A(_11865_),
    .Y(_13125_));
 sky130_fd_sc_hd__inv_1 _19686_ (.A(_11873_),
    .Y(_13129_));
 sky130_fd_sc_hd__clkinv_1 _19687_ (.A(_11881_),
    .Y(_13133_));
 sky130_fd_sc_hd__inv_2 _19688_ (.A(_11889_),
    .Y(_13137_));
 sky130_fd_sc_hd__clkinv_1 _19689_ (.A(_11897_),
    .Y(_13141_));
 sky130_fd_sc_hd__clkinv_1 _19690_ (.A(_11905_),
    .Y(_13145_));
 sky130_fd_sc_hd__clkinv_1 _19691_ (.A(_11913_),
    .Y(_13149_));
 sky130_fd_sc_hd__clkinv_1 _19692_ (.A(_11921_),
    .Y(_13153_));
 sky130_fd_sc_hd__inv_1 _19693_ (.A(_11929_),
    .Y(_13157_));
 sky130_fd_sc_hd__inv_1 _19694_ (.A(_11937_),
    .Y(_13161_));
 sky130_fd_sc_hd__inv_1 _19695_ (.A(_11945_),
    .Y(_13165_));
 sky130_fd_sc_hd__inv_1 _19696_ (.A(_11953_),
    .Y(_13169_));
 sky130_fd_sc_hd__clkinv_1 _19697_ (.A(_11961_),
    .Y(_13173_));
 sky130_fd_sc_hd__clkinv_1 _19698_ (.A(_11969_),
    .Y(_13177_));
 sky130_fd_sc_hd__clkinv_1 _19699_ (.A(_11977_),
    .Y(_13181_));
 sky130_fd_sc_hd__inv_1 _19700_ (.A(_11985_),
    .Y(_13185_));
 sky130_fd_sc_hd__inv_1 _19701_ (.A(_11993_),
    .Y(_13189_));
 sky130_fd_sc_hd__clkinv_1 _19702_ (.A(_12001_),
    .Y(_13193_));
 sky130_fd_sc_hd__clkinv_1 _19703_ (.A(_12009_),
    .Y(_13197_));
 sky130_fd_sc_hd__inv_1 _19704_ (.A(_12017_),
    .Y(_13201_));
 sky130_fd_sc_hd__inv_1 _19705_ (.A(_12025_),
    .Y(_13205_));
 sky130_fd_sc_hd__clkinv_1 _19706_ (.A(_12033_),
    .Y(_13209_));
 sky130_fd_sc_hd__clkinv_1 _19707_ (.A(_12041_),
    .Y(_13213_));
 sky130_fd_sc_hd__inv_1 _19708_ (.A(_12049_),
    .Y(_13217_));
 sky130_fd_sc_hd__inv_1 _19709_ (.A(_12057_),
    .Y(_13221_));
 sky130_fd_sc_hd__inv_1 _19710_ (.A(_12065_),
    .Y(_13225_));
 sky130_fd_sc_hd__mux2_1 _19711_ (.A0(\hash.CA2.f_dash[0] ),
    .A1(\hash.CA2.e_dash[0] ),
    .S(\hash.CA2.S1.X[0] ),
    .X(_13229_));
 sky130_fd_sc_hd__inv_1 _19712_ (.A(_12078_),
    .Y(_12092_));
 sky130_fd_sc_hd__mux2_4 _19713_ (.A0(\hash.CA2.f_dash[2] ),
    .A1(\hash.CA2.e_dash[2] ),
    .S(\hash.CA2.S1.X[2] ),
    .X(_13242_));
 sky130_fd_sc_hd__inv_1 _19714_ (.A(_12090_),
    .Y(_12101_));
 sky130_fd_sc_hd__mux2_1 _19715_ (.A0(\hash.CA2.f_dash[3] ),
    .A1(\hash.CA2.e_dash[3] ),
    .S(\hash.CA2.S1.X[3] ),
    .X(_13249_));
 sky130_fd_sc_hd__inv_1 _19716_ (.A(_12099_),
    .Y(_12115_));
 sky130_fd_sc_hd__mux2_1 _19717_ (.A0(\hash.CA2.f_dash[4] ),
    .A1(\hash.CA2.e_dash[4] ),
    .S(\hash.CA2.S1.X[4] ),
    .X(_13256_));
 sky130_fd_sc_hd__inv_1 _19718_ (.A(_12113_),
    .Y(_12124_));
 sky130_fd_sc_hd__mux2_8 _19719_ (.A0(\hash.CA2.f_dash[5] ),
    .A1(\hash.CA2.e_dash[5] ),
    .S(\hash.CA2.S1.X[5] ),
    .X(_13263_));
 sky130_fd_sc_hd__inv_1 _19720_ (.A(_12122_),
    .Y(_12133_));
 sky130_fd_sc_hd__mux2_1 _19721_ (.A0(\hash.CA2.f_dash[6] ),
    .A1(\hash.CA2.e_dash[6] ),
    .S(\hash.CA2.S1.X[6] ),
    .X(_13270_));
 sky130_fd_sc_hd__inv_1 _19722_ (.A(_12131_),
    .Y(_12142_));
 sky130_fd_sc_hd__mux2_1 _19723_ (.A0(\hash.CA2.f_dash[7] ),
    .A1(\hash.CA2.e_dash[7] ),
    .S(net1058),
    .X(_13277_));
 sky130_fd_sc_hd__inv_1 _19724_ (.A(_12140_),
    .Y(_12151_));
 sky130_fd_sc_hd__mux2_1 _19725_ (.A0(\hash.CA2.f_dash[8] ),
    .A1(\hash.CA2.e_dash[8] ),
    .S(\hash.CA2.S1.X[8] ),
    .X(_13284_));
 sky130_fd_sc_hd__inv_1 _19726_ (.A(_12149_),
    .Y(_12160_));
 sky130_fd_sc_hd__mux2_4 _19727_ (.A0(\hash.CA2.f_dash[9] ),
    .A1(\hash.CA2.e_dash[9] ),
    .S(\hash.CA2.S1.X[9] ),
    .X(_13291_));
 sky130_fd_sc_hd__inv_1 _19728_ (.A(_12158_),
    .Y(_12169_));
 sky130_fd_sc_hd__mux2_8 _19729_ (.A0(\hash.CA2.f_dash[10] ),
    .A1(\hash.CA2.e_dash[10] ),
    .S(\hash.CA2.S1.X[10] ),
    .X(_13298_));
 sky130_fd_sc_hd__inv_1 _19730_ (.A(_12167_),
    .Y(_12178_));
 sky130_fd_sc_hd__mux2_4 _19731_ (.A0(\hash.CA2.f_dash[11] ),
    .A1(\hash.CA2.e_dash[11] ),
    .S(\hash.CA2.S1.X[11] ),
    .X(_13305_));
 sky130_fd_sc_hd__inv_1 _19732_ (.A(_12176_),
    .Y(_12187_));
 sky130_fd_sc_hd__mux2_4 _19733_ (.A0(\hash.CA2.f_dash[12] ),
    .A1(\hash.CA2.e_dash[12] ),
    .S(\hash.CA2.S1.X[12] ),
    .X(_13312_));
 sky130_fd_sc_hd__inv_1 _19734_ (.A(_12185_),
    .Y(_12196_));
 sky130_fd_sc_hd__nand2_1 _19735_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA2.e_dash[13] ),
    .Y(_07908_));
 sky130_fd_sc_hd__o21ai_2 _19736_ (.A1(\hash.CA2.S1.X[13] ),
    .A2(_06314_),
    .B1(_07908_),
    .Y(_13319_));
 sky130_fd_sc_hd__inv_1 _19737_ (.A(_12194_),
    .Y(_12205_));
 sky130_fd_sc_hd__mux2_8 _19738_ (.A0(\hash.CA2.f_dash[14] ),
    .A1(\hash.CA2.e_dash[14] ),
    .S(\hash.CA2.S1.X[14] ),
    .X(_13326_));
 sky130_fd_sc_hd__inv_1 _19739_ (.A(_12203_),
    .Y(_12214_));
 sky130_fd_sc_hd__mux2_4 _19740_ (.A0(\hash.CA2.f_dash[15] ),
    .A1(\hash.CA2.e_dash[15] ),
    .S(\hash.CA2.S1.X[15] ),
    .X(_13333_));
 sky130_fd_sc_hd__inv_1 _19741_ (.A(_12212_),
    .Y(_12223_));
 sky130_fd_sc_hd__mux2_1 _19742_ (.A0(\hash.CA2.f_dash[16] ),
    .A1(\hash.CA2.e_dash[16] ),
    .S(\hash.CA2.S1.X[16] ),
    .X(_13340_));
 sky130_fd_sc_hd__inv_1 _19743_ (.A(_12221_),
    .Y(_12232_));
 sky130_fd_sc_hd__mux2_1 _19744_ (.A0(\hash.CA2.f_dash[17] ),
    .A1(\hash.CA2.e_dash[17] ),
    .S(\hash.CA2.S1.X[17] ),
    .X(_13347_));
 sky130_fd_sc_hd__inv_1 _19745_ (.A(_12230_),
    .Y(_12241_));
 sky130_fd_sc_hd__mux2_8 _19746_ (.A0(\hash.CA2.f_dash[18] ),
    .A1(\hash.CA2.e_dash[18] ),
    .S(\hash.CA2.S1.X[18] ),
    .X(_13354_));
 sky130_fd_sc_hd__inv_1 _19747_ (.A(_12239_),
    .Y(_12250_));
 sky130_fd_sc_hd__mux2_8 _19748_ (.A0(\hash.CA2.f_dash[19] ),
    .A1(\hash.CA2.e_dash[19] ),
    .S(\hash.CA2.S1.X[19] ),
    .X(_13361_));
 sky130_fd_sc_hd__inv_1 _19749_ (.A(_12248_),
    .Y(_12259_));
 sky130_fd_sc_hd__mux2_4 _19750_ (.A0(\hash.CA2.f_dash[20] ),
    .A1(\hash.CA2.e_dash[20] ),
    .S(\hash.CA2.S1.X[20] ),
    .X(_13368_));
 sky130_fd_sc_hd__inv_1 _19751_ (.A(_12257_),
    .Y(_12268_));
 sky130_fd_sc_hd__mux2_1 _19752_ (.A0(\hash.CA2.f_dash[21] ),
    .A1(\hash.CA2.e_dash[21] ),
    .S(\hash.CA2.S1.X[21] ),
    .X(_13375_));
 sky130_fd_sc_hd__inv_1 _19753_ (.A(_12266_),
    .Y(_12277_));
 sky130_fd_sc_hd__mux2_1 _19754_ (.A0(\hash.CA2.f_dash[22] ),
    .A1(\hash.CA2.e_dash[22] ),
    .S(\hash.CA2.S1.X[22] ),
    .X(_13382_));
 sky130_fd_sc_hd__inv_1 _19755_ (.A(_12275_),
    .Y(_12286_));
 sky130_fd_sc_hd__mux2_8 _19756_ (.A0(\hash.CA2.f_dash[23] ),
    .A1(\hash.CA2.e_dash[23] ),
    .S(\hash.CA2.S1.X[23] ),
    .X(_13389_));
 sky130_fd_sc_hd__inv_1 _19757_ (.A(_12284_),
    .Y(_12295_));
 sky130_fd_sc_hd__mux2_8 _19758_ (.A0(\hash.CA2.f_dash[24] ),
    .A1(\hash.CA2.e_dash[24] ),
    .S(\hash.CA2.S1.X[24] ),
    .X(_13396_));
 sky130_fd_sc_hd__inv_1 _19759_ (.A(_12293_),
    .Y(_12304_));
 sky130_fd_sc_hd__mux2_1 _19760_ (.A0(\hash.CA2.f_dash[25] ),
    .A1(\hash.CA2.e_dash[25] ),
    .S(\hash.CA2.S1.X[25] ),
    .X(_13403_));
 sky130_fd_sc_hd__inv_1 _19761_ (.A(_12302_),
    .Y(_12313_));
 sky130_fd_sc_hd__mux2_8 _19762_ (.A0(\hash.CA2.f_dash[26] ),
    .A1(\hash.CA2.e_dash[26] ),
    .S(net1064),
    .X(_13410_));
 sky130_fd_sc_hd__inv_1 _19763_ (.A(_12311_),
    .Y(_12322_));
 sky130_fd_sc_hd__mux2_8 _19764_ (.A0(\hash.CA2.f_dash[27] ),
    .A1(\hash.CA2.e_dash[27] ),
    .S(\hash.CA2.S1.X[27] ),
    .X(_13417_));
 sky130_fd_sc_hd__inv_1 _19765_ (.A(_12320_),
    .Y(_12331_));
 sky130_fd_sc_hd__mux2_8 _19766_ (.A0(\hash.CA2.f_dash[28] ),
    .A1(\hash.CA2.e_dash[28] ),
    .S(\hash.CA2.S1.X[28] ),
    .X(_13424_));
 sky130_fd_sc_hd__inv_1 _19767_ (.A(_12329_),
    .Y(_12340_));
 sky130_fd_sc_hd__mux2_4 _19768_ (.A0(\hash.CA2.f_dash[29] ),
    .A1(\hash.CA2.e_dash[29] ),
    .S(\hash.CA2.S1.X[29] ),
    .X(_13431_));
 sky130_fd_sc_hd__inv_1 _19769_ (.A(_12338_),
    .Y(_12349_));
 sky130_fd_sc_hd__mux2_8 _19770_ (.A0(\hash.CA2.f_dash[30] ),
    .A1(\hash.CA2.e_dash[30] ),
    .S(\hash.CA2.S1.X[30] ),
    .X(_13438_));
 sky130_fd_sc_hd__inv_1 _19771_ (.A(_12347_),
    .Y(_12358_));
 sky130_fd_sc_hd__inv_4 _19772_ (.A(\count_1[1] ),
    .Y(_00650_));
 sky130_fd_sc_hd__inv_4 _19773_ (.A(\count_2[1] ),
    .Y(_00652_));
 sky130_fd_sc_hd__a21oi_1 _19774_ (.A1(\hash.CA2.a_dash[2] ),
    .A2(_05998_),
    .B1(_04421_),
    .Y(_07909_));
 sky130_fd_sc_hd__nor2_1 _19775_ (.A(\hash.CA2.a_dash[2] ),
    .B(_05998_),
    .Y(_07910_));
 sky130_fd_sc_hd__o21ai_0 _19776_ (.A1(_07909_),
    .A2(_07910_),
    .B1(_06002_),
    .Y(_13551_));
 sky130_fd_sc_hd__o21ai_0 _19777_ (.A1(\hash.CA1.S0.X[3] ),
    .A2(\hash.CA1.b[3] ),
    .B1(\hash.CA2.a_dash[3] ),
    .Y(_07911_));
 sky130_fd_sc_hd__nand2_1 _19778_ (.A(_04470_),
    .B(\hash.CA1.S0.X[3] ),
    .Y(_07912_));
 sky130_fd_sc_hd__nand2_1 _19779_ (.A(_07911_),
    .B(_07912_),
    .Y(_13555_));
 sky130_fd_sc_hd__nor2_1 _19780_ (.A(_06010_),
    .B(\hash.CA1.b[4] ),
    .Y(_07913_));
 sky130_fd_sc_hd__a21oi_1 _19781_ (.A1(_04487_),
    .A2(_06010_),
    .B1(\hash.CA2.a_dash[4] ),
    .Y(_07914_));
 sky130_fd_sc_hd__nor2_1 _19782_ (.A(_07913_),
    .B(_07914_),
    .Y(_13559_));
 sky130_fd_sc_hd__nor2_1 _19783_ (.A(net349),
    .B(_04501_),
    .Y(_07915_));
 sky130_fd_sc_hd__nor2_1 _19784_ (.A(_06016_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__o22a_1 _19785_ (.A1(\hash.CA1.S0.X[5] ),
    .A2(\hash.CA1.b[5] ),
    .B1(_07916_),
    .B2(\hash.CA2.a_dash[5] ),
    .X(_13563_));
 sky130_fd_sc_hd__nor2_1 _19786_ (.A(net349),
    .B(_04522_),
    .Y(_07917_));
 sky130_fd_sc_hd__o21ai_0 _19787_ (.A1(\hash.CA1.S0.X[6] ),
    .A2(\hash.CA1.b[6] ),
    .B1(\hash.CA2.a_dash[6] ),
    .Y(_07918_));
 sky130_fd_sc_hd__o21ai_0 _19788_ (.A1(_06024_),
    .A2(_07917_),
    .B1(_07918_),
    .Y(_13567_));
 sky130_fd_sc_hd__nand2_1 _19789_ (.A(_06030_),
    .B(_06031_),
    .Y(_07919_));
 sky130_fd_sc_hd__a21oi_1 _19790_ (.A1(\hash.CA1.S0.X[7] ),
    .A2(\hash.CA1.b[7] ),
    .B1(\hash.CA2.a_dash[7] ),
    .Y(_07920_));
 sky130_fd_sc_hd__a211oi_1 _19791_ (.A1(_04543_),
    .A2(_07919_),
    .B1(_07920_),
    .C1(net349),
    .Y(_13571_));
 sky130_fd_sc_hd__maj3_1 _19792_ (.A(\hash.CA2.a_dash[8] ),
    .B(_06043_),
    .C(_06279_),
    .X(_13575_));
 sky130_fd_sc_hd__maj3_1 _19793_ (.A(\hash.CA2.a_dash[9] ),
    .B(\hash.CA1.S0.X[9] ),
    .C(_06280_),
    .X(_13579_));
 sky130_fd_sc_hd__maj3_1 _19794_ (.A(\hash.CA2.a_dash[10] ),
    .B(\hash.CA1.S0.X[10] ),
    .C(\hash.CA1.b[10] ),
    .X(_13583_));
 sky130_fd_sc_hd__o211ai_1 _19795_ (.A1(_04614_),
    .A2(_06065_),
    .B1(_06002_),
    .C1(\hash.CA2.a_dash[11] ),
    .Y(_07921_));
 sky130_fd_sc_hd__o21ai_2 _19796_ (.A1(_06066_),
    .A2(_06282_),
    .B1(_07921_),
    .Y(_13587_));
 sky130_fd_sc_hd__maj3_1 _19797_ (.A(\hash.CA2.a_dash[12] ),
    .B(\hash.CA1.S0.X[12] ),
    .C(_06283_),
    .X(_13591_));
 sky130_fd_sc_hd__a21oi_1 _19798_ (.A1(\hash.CA2.a_dash[13] ),
    .A2(_04437_),
    .B1(_06079_),
    .Y(_07922_));
 sky130_fd_sc_hd__o21ai_4 _19799_ (.A1(_04638_),
    .A2(_07922_),
    .B1(_06002_),
    .Y(_13595_));
 sky130_fd_sc_hd__a21boi_0 _19800_ (.A1(\hash.CA2.a_dash[14] ),
    .A2(_04636_),
    .B1_N(_06091_),
    .Y(_07923_));
 sky130_fd_sc_hd__o21ai_2 _19801_ (.A1(_04646_),
    .A2(_07923_),
    .B1(_06002_),
    .Y(_13599_));
 sky130_fd_sc_hd__maj3_1 _19802_ (.A(\hash.CA2.a_dash[15] ),
    .B(\hash.CA1.S0.X[15] ),
    .C(\hash.CA1.b[15] ),
    .X(_13603_));
 sky130_fd_sc_hd__maj3_1 _19803_ (.A(\hash.CA2.a_dash[16] ),
    .B(\hash.CA1.S0.X[16] ),
    .C(\hash.CA1.b[16] ),
    .X(_13607_));
 sky130_fd_sc_hd__nor2_1 _19804_ (.A(\hash.CA2.a_dash[17] ),
    .B(_04520_),
    .Y(_07924_));
 sky130_fd_sc_hd__a21oi_1 _19805_ (.A1(\hash.CA2.a_dash[17] ),
    .A2(_04520_),
    .B1(\hash.CA1.S0.X[17] ),
    .Y(_07925_));
 sky130_fd_sc_hd__o21ai_1 _19806_ (.A1(_07924_),
    .A2(_07925_),
    .B1(_06002_),
    .Y(_13611_));
 sky130_fd_sc_hd__a21oi_1 _19807_ (.A1(\hash.CA2.a_dash[18] ),
    .A2(_04541_),
    .B1(_06121_),
    .Y(_07926_));
 sky130_fd_sc_hd__o21ai_2 _19808_ (.A1(_04672_),
    .A2(_07926_),
    .B1(_06002_),
    .Y(_13615_));
 sky130_fd_sc_hd__a211oi_1 _19809_ (.A1(_04559_),
    .A2(_06132_),
    .B1(net350),
    .C1(\hash.CA2.a_dash[19] ),
    .Y(_07927_));
 sky130_fd_sc_hd__nor2_1 _19810_ (.A(\hash.CA1.S0.X[19] ),
    .B(_06284_),
    .Y(_07928_));
 sky130_fd_sc_hd__nor2_2 _19811_ (.A(_07927_),
    .B(_07928_),
    .Y(_13619_));
 sky130_fd_sc_hd__nand2_1 _19812_ (.A(_04577_),
    .B(_06148_),
    .Y(_07929_));
 sky130_fd_sc_hd__o21ai_2 _19813_ (.A1(_06148_),
    .A2(\hash.CA1.b[20] ),
    .B1(\hash.CA2.a_dash[20] ),
    .Y(_07930_));
 sky130_fd_sc_hd__nand2_4 _19814_ (.A(_07929_),
    .B(_07930_),
    .Y(_13623_));
 sky130_fd_sc_hd__a21oi_1 _19815_ (.A1(\hash.CA2.a_dash[21] ),
    .A2(_04596_),
    .B1(_06155_),
    .Y(_07931_));
 sky130_fd_sc_hd__o21ai_2 _19816_ (.A1(_04697_),
    .A2(_07931_),
    .B1(_06002_),
    .Y(_13627_));
 sky130_fd_sc_hd__nand2_1 _19817_ (.A(_04704_),
    .B(_06164_),
    .Y(_07932_));
 sky130_fd_sc_hd__o21ai_2 _19818_ (.A1(\hash.CA2.a_dash[22] ),
    .A2(_04420_),
    .B1(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__nand2_1 _19819_ (.A(_06002_),
    .B(_07933_),
    .Y(_13631_));
 sky130_fd_sc_hd__o21ai_0 _19820_ (.A1(\hash.CA1.S0.X[23] ),
    .A2(_06285_),
    .B1(\hash.CA2.a_dash[23] ),
    .Y(_07934_));
 sky130_fd_sc_hd__o21ai_2 _19821_ (.A1(_06172_),
    .A2(_06895_),
    .B1(_07934_),
    .Y(_13635_));
 sky130_fd_sc_hd__o31a_1 _19822_ (.A1(_13402_),
    .A2(_13394_),
    .A3(_06177_),
    .B1(_06178_),
    .X(_07935_));
 sky130_fd_sc_hd__o21ai_0 _19823_ (.A1(\hash.CA2.a_dash[24] ),
    .A2(_04726_),
    .B1(_07935_),
    .Y(_07936_));
 sky130_fd_sc_hd__a21oi_2 _19824_ (.A1(_04727_),
    .A2(_07936_),
    .B1(net351),
    .Y(_13639_));
 sky130_fd_sc_hd__maj3_4 _19825_ (.A(\hash.CA2.a_dash[25] ),
    .B(\hash.CA1.S0.X[25] ),
    .C(\hash.CA1.b[25] ),
    .X(_13643_));
 sky130_fd_sc_hd__maj3_4 _19826_ (.A(\hash.CA2.a_dash[26] ),
    .B(_06201_),
    .C(\hash.CA1.b[26] ),
    .X(_13647_));
 sky130_fd_sc_hd__maj3_1 _19827_ (.A(\hash.CA2.a_dash[27] ),
    .B(_04537_),
    .C(_06210_),
    .X(_07937_));
 sky130_fd_sc_hd__or2_4 _19828_ (.A(net350),
    .B(_07937_),
    .X(_13651_));
 sky130_fd_sc_hd__o21ai_0 _19829_ (.A1(_06215_),
    .A2(_06217_),
    .B1(_04756_),
    .Y(_07938_));
 sky130_fd_sc_hd__o21ai_1 _19830_ (.A1(\hash.CA2.a_dash[28] ),
    .A2(_04554_),
    .B1(_07938_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_2 _19831_ (.A(_06002_),
    .B(_07939_),
    .Y(_13655_));
 sky130_fd_sc_hd__a21oi_1 _19832_ (.A1(\hash.CA2.a_dash[29] ),
    .A2(_04754_),
    .B1(\hash.CA1.S0.X[29] ),
    .Y(_07940_));
 sky130_fd_sc_hd__o21ai_4 _19833_ (.A1(_04762_),
    .A2(_07940_),
    .B1(_06002_),
    .Y(_13659_));
 sky130_fd_sc_hd__a31oi_1 _19834_ (.A1(_04770_),
    .A2(_06232_),
    .A3(_06233_),
    .B1(_04771_),
    .Y(_07941_));
 sky130_fd_sc_hd__nor2_2 _19835_ (.A(net351),
    .B(_07941_),
    .Y(_13663_));
 sky130_fd_sc_hd__inv_1 _19836_ (.A(_12373_),
    .Y(_13667_));
 sky130_fd_sc_hd__clkinv_1 _19837_ (.A(_12369_),
    .Y(_12379_));
 sky130_fd_sc_hd__xor2_1 _19838_ (.A(_13678_),
    .B(_12380_),
    .X(\hash.CA1.p4[3] ));
 sky130_fd_sc_hd__inv_1 _19839_ (.A(_12384_),
    .Y(_13682_));
 sky130_fd_sc_hd__a21o_1 _19840_ (.A1(_12378_),
    .A2(_13672_),
    .B1(_13671_),
    .X(_07942_));
 sky130_fd_sc_hd__a21oi_1 _19841_ (.A1(_13678_),
    .A2(_07942_),
    .B1(_13677_),
    .Y(_07943_));
 sky130_fd_sc_hd__xnor2_1 _19842_ (.A(_13684_),
    .B(_07943_),
    .Y(\hash.CA1.p4[4] ));
 sky130_fd_sc_hd__a21o_1 _19843_ (.A1(_13678_),
    .A2(_12380_),
    .B1(_13677_),
    .X(_07944_));
 sky130_fd_sc_hd__a21oi_2 _19844_ (.A1(_13684_),
    .A2(_07944_),
    .B1(_13683_),
    .Y(_07945_));
 sky130_fd_sc_hd__xnor2_1 _19845_ (.A(_13690_),
    .B(_07945_),
    .Y(\hash.CA1.p4[5] ));
 sky130_fd_sc_hd__inv_1 _19846_ (.A(_12392_),
    .Y(_13694_));
 sky130_fd_sc_hd__inv_1 _19847_ (.A(_13684_),
    .Y(_07946_));
 sky130_fd_sc_hd__o21bai_1 _19848_ (.A1(_07946_),
    .A2(_07943_),
    .B1_N(_13683_),
    .Y(_07947_));
 sky130_fd_sc_hd__a21o_4 _19849_ (.A1(_13690_),
    .A2(_07947_),
    .B1(_13689_),
    .X(_07948_));
 sky130_fd_sc_hd__xor2_2 _19850_ (.A(_13696_),
    .B(_07948_),
    .X(\hash.CA1.p4[6] ));
 sky130_fd_sc_hd__inv_1 _19851_ (.A(_13690_),
    .Y(_07949_));
 sky130_fd_sc_hd__o21bai_2 _19852_ (.A1(_07949_),
    .A2(_07945_),
    .B1_N(_13689_),
    .Y(_07950_));
 sky130_fd_sc_hd__a21oi_2 _19853_ (.A1(_13696_),
    .A2(_07950_),
    .B1(_13695_),
    .Y(_07951_));
 sky130_fd_sc_hd__xnor2_1 _19854_ (.A(_13702_),
    .B(_07951_),
    .Y(\hash.CA1.p4[7] ));
 sky130_fd_sc_hd__clkinv_2 _19855_ (.A(_12400_),
    .Y(_13706_));
 sky130_fd_sc_hd__a21oi_2 _19856_ (.A1(_13696_),
    .A2(_07948_),
    .B1(_13695_),
    .Y(_07952_));
 sky130_fd_sc_hd__inv_1 _19857_ (.A(_07952_),
    .Y(_07953_));
 sky130_fd_sc_hd__a21oi_1 _19858_ (.A1(_13702_),
    .A2(_07953_),
    .B1(_13701_),
    .Y(_07954_));
 sky130_fd_sc_hd__xnor2_1 _19859_ (.A(_13709_),
    .B(_07954_),
    .Y(\hash.CA1.p4[8] ));
 sky130_fd_sc_hd__clkinv_1 _19860_ (.A(_12405_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand2_4 _19861_ (.A(_13702_),
    .B(_13709_),
    .Y(_07955_));
 sky130_fd_sc_hd__a21oi_2 _19862_ (.A1(_13709_),
    .A2(_13701_),
    .B1(_13708_),
    .Y(_07956_));
 sky130_fd_sc_hd__o21ai_0 _19863_ (.A1(_07951_),
    .A2(_07955_),
    .B1(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__xor2_1 _19864_ (.A(_13715_),
    .B(_07957_),
    .X(\hash.CA1.p4[9] ));
 sky130_fd_sc_hd__nand2b_1 _19865_ (.A_N(_13714_),
    .B(_07956_),
    .Y(_07958_));
 sky130_fd_sc_hd__o21bai_4 _19866_ (.A1(_07952_),
    .A2(_07955_),
    .B1_N(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__o21a_4 _19867_ (.A1(_13715_),
    .A2(_13714_),
    .B1(_13720_),
    .X(_07960_));
 sky130_fd_sc_hd__o21ai_0 _19868_ (.A1(_07952_),
    .A2(_07955_),
    .B1(_07956_),
    .Y(_07961_));
 sky130_fd_sc_hd__a211oi_1 _19869_ (.A1(_13715_),
    .A2(_07961_),
    .B1(_13714_),
    .C1(_13720_),
    .Y(_07962_));
 sky130_fd_sc_hd__a21oi_4 _19870_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_07962_),
    .Y(\hash.CA1.p4[10] ));
 sky130_fd_sc_hd__a211oi_1 _19871_ (.A1(_13696_),
    .A2(_07950_),
    .B1(_07958_),
    .C1(_13695_),
    .Y(_07963_));
 sky130_fd_sc_hd__a21boi_0 _19872_ (.A1(_07956_),
    .A2(_07955_),
    .B1_N(_13715_),
    .Y(_07964_));
 sky130_fd_sc_hd__o21ai_1 _19873_ (.A1(_13714_),
    .A2(_07964_),
    .B1(_13720_),
    .Y(_07965_));
 sky130_fd_sc_hd__nor2_1 _19874_ (.A(_07963_),
    .B(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__nor2_2 _19875_ (.A(_13719_),
    .B(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__xnor2_2 _19876_ (.A(_13726_),
    .B(_07967_),
    .Y(\hash.CA1.p4[11] ));
 sky130_fd_sc_hd__clkinv_1 _19877_ (.A(_12416_),
    .Y(_13730_));
 sky130_fd_sc_hd__inv_1 _19878_ (.A(_13726_),
    .Y(_07968_));
 sky130_fd_sc_hd__a21oi_1 _19879_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_13719_),
    .Y(_07969_));
 sky130_fd_sc_hd__o21bai_1 _19880_ (.A1(_07968_),
    .A2(_07969_),
    .B1_N(_13725_),
    .Y(_07970_));
 sky130_fd_sc_hd__xor2_2 _19881_ (.A(_13733_),
    .B(_07970_),
    .X(\hash.CA1.p4[12] ));
 sky130_fd_sc_hd__inv_1 _19882_ (.A(_12421_),
    .Y(_13737_));
 sky130_fd_sc_hd__o21bai_1 _19883_ (.A1(_07968_),
    .A2(_07967_),
    .B1_N(_13725_),
    .Y(_07971_));
 sky130_fd_sc_hd__a21oi_1 _19884_ (.A1(_13733_),
    .A2(_07971_),
    .B1(_13732_),
    .Y(_07972_));
 sky130_fd_sc_hd__xnor2_2 _19885_ (.A(_13739_),
    .B(_07972_),
    .Y(\hash.CA1.p4[13] ));
 sky130_fd_sc_hd__a2111oi_2 _19886_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_13719_),
    .C1(_13725_),
    .D1(_13732_),
    .Y(_07973_));
 sky130_fd_sc_hd__o21a_1 _19887_ (.A1(_13726_),
    .A2(_13725_),
    .B1(_13733_),
    .X(_07974_));
 sky130_fd_sc_hd__nor2_1 _19888_ (.A(_13732_),
    .B(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__nor2_1 _19889_ (.A(_07973_),
    .B(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__a21oi_1 _19890_ (.A1(_13739_),
    .A2(_07976_),
    .B1(_13738_),
    .Y(_07977_));
 sky130_fd_sc_hd__xnor2_2 _19891_ (.A(_13745_),
    .B(_07977_),
    .Y(\hash.CA1.p4[14] ));
 sky130_fd_sc_hd__inv_1 _19892_ (.A(_12429_),
    .Y(_13749_));
 sky130_fd_sc_hd__nand3_1 _19893_ (.A(_13726_),
    .B(_13733_),
    .C(_13739_),
    .Y(_07978_));
 sky130_fd_sc_hd__a21o_1 _19894_ (.A1(_13733_),
    .A2(_13725_),
    .B1(_13732_),
    .X(_07979_));
 sky130_fd_sc_hd__a21oi_1 _19895_ (.A1(_13739_),
    .A2(_07979_),
    .B1(_13738_),
    .Y(_07980_));
 sky130_fd_sc_hd__o21ai_0 _19896_ (.A1(_07967_),
    .A2(_07978_),
    .B1(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__a21oi_1 _19897_ (.A1(_13745_),
    .A2(_07981_),
    .B1(_13744_),
    .Y(_07982_));
 sky130_fd_sc_hd__xnor2_2 _19898_ (.A(_13752_),
    .B(_07982_),
    .Y(\hash.CA1.p4[15] ));
 sky130_fd_sc_hd__inv_1 _19899_ (.A(_12434_),
    .Y(_13756_));
 sky130_fd_sc_hd__and2_4 _19900_ (.A(_13745_),
    .B(_13752_),
    .X(_07983_));
 sky130_fd_sc_hd__o211ai_1 _19901_ (.A1(_13732_),
    .A2(_07974_),
    .B1(_07983_),
    .C1(_13739_),
    .Y(_07984_));
 sky130_fd_sc_hd__a22oi_1 _19902_ (.A1(_13752_),
    .A2(_13744_),
    .B1(_07983_),
    .B2(_13738_),
    .Y(_07985_));
 sky130_fd_sc_hd__nor2b_1 _19903_ (.A(_13751_),
    .B_N(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__o21ai_2 _19904_ (.A1(_07973_),
    .A2(_07984_),
    .B1(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__xor2_2 _19905_ (.A(_13759_),
    .B(_07987_),
    .X(\hash.CA1.p4[16] ));
 sky130_fd_sc_hd__inv_1 _19906_ (.A(_12439_),
    .Y(_13763_));
 sky130_fd_sc_hd__nor3_1 _19907_ (.A(_07963_),
    .B(_07965_),
    .C(_07978_),
    .Y(_07988_));
 sky130_fd_sc_hd__inv_1 _19908_ (.A(_13719_),
    .Y(_07989_));
 sky130_fd_sc_hd__o21ai_0 _19909_ (.A1(_07989_),
    .A2(_07978_),
    .B1(_07980_),
    .Y(_07990_));
 sky130_fd_sc_hd__o211ai_1 _19910_ (.A1(_07988_),
    .A2(_07990_),
    .B1(_07983_),
    .C1(_13759_),
    .Y(_07991_));
 sky130_fd_sc_hd__and3_1 _19911_ (.A(_13752_),
    .B(_13759_),
    .C(_13744_),
    .X(_07992_));
 sky130_fd_sc_hd__a21oi_2 _19912_ (.A1(_13759_),
    .A2(_13751_),
    .B1(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__nand3b_1 _19913_ (.A_N(_13758_),
    .B(_07991_),
    .C(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__xor2_2 _19914_ (.A(_13766_),
    .B(_07994_),
    .X(\hash.CA1.p4[17] ));
 sky130_fd_sc_hd__clkinv_1 _19915_ (.A(_12444_),
    .Y(_13770_));
 sky130_fd_sc_hd__nor3_1 _19916_ (.A(_13751_),
    .B(_13758_),
    .C(_13765_),
    .Y(_07995_));
 sky130_fd_sc_hd__o211ai_1 _19917_ (.A1(_07973_),
    .A2(_07984_),
    .B1(_07985_),
    .C1(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__or2_0 _19918_ (.A(_13766_),
    .B(_13765_),
    .X(_07997_));
 sky130_fd_sc_hd__o31a_1 _19919_ (.A1(_13759_),
    .A2(_13758_),
    .A3(_13765_),
    .B1(_07997_),
    .X(_07998_));
 sky130_fd_sc_hd__nand2_4 _19920_ (.A(_07996_),
    .B(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__xnor2_2 _19921_ (.A(_13772_),
    .B(_07999_),
    .Y(\hash.CA1.p4[18] ));
 sky130_fd_sc_hd__nor3_1 _19922_ (.A(_13758_),
    .B(_13765_),
    .C(_13771_),
    .Y(_08000_));
 sky130_fd_sc_hd__a21oi_1 _19923_ (.A1(_13772_),
    .A2(_07997_),
    .B1(_13771_),
    .Y(_08001_));
 sky130_fd_sc_hd__a31oi_4 _19924_ (.A1(_07991_),
    .A2(_07993_),
    .A3(_08000_),
    .B1(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__xor2_2 _19925_ (.A(_13777_),
    .B(_08002_),
    .X(\hash.CA1.p4[19] ));
 sky130_fd_sc_hd__nand3_2 _19926_ (.A(_13772_),
    .B(_13777_),
    .C(_13782_),
    .Y(_08003_));
 sky130_fd_sc_hd__and3_1 _19927_ (.A(_13777_),
    .B(_13782_),
    .C(_13771_),
    .X(_08004_));
 sky130_fd_sc_hd__a21oi_2 _19928_ (.A1(_13782_),
    .A2(_13776_),
    .B1(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__o21ai_4 _19929_ (.A1(_07999_),
    .A2(_08003_),
    .B1(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__a31o_1 _19930_ (.A1(_13772_),
    .A2(_07996_),
    .A3(_07998_),
    .B1(_13771_),
    .X(_08007_));
 sky130_fd_sc_hd__a211oi_2 _19931_ (.A1(_13777_),
    .A2(_08007_),
    .B1(_13776_),
    .C1(_13782_),
    .Y(_08008_));
 sky130_fd_sc_hd__nor2_4 _19932_ (.A(_08006_),
    .B(_08008_),
    .Y(\hash.CA1.p4[20] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_984 ();
 sky130_fd_sc_hd__a21o_1 _19934_ (.A1(_13777_),
    .A2(_08002_),
    .B1(_13776_),
    .X(_08010_));
 sky130_fd_sc_hd__a21oi_1 _19935_ (.A1(_13782_),
    .A2(_08010_),
    .B1(_13781_),
    .Y(_08011_));
 sky130_fd_sc_hd__xnor2_2 _19936_ (.A(_13787_),
    .B(_08011_),
    .Y(\hash.CA1.p4[21] ));
 sky130_fd_sc_hd__inv_1 _19937_ (.A(_13781_),
    .Y(_08012_));
 sky130_fd_sc_hd__o211ai_1 _19938_ (.A1(_07999_),
    .A2(_08003_),
    .B1(_08005_),
    .C1(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__a21oi_2 _19939_ (.A1(_13787_),
    .A2(_08013_),
    .B1(_13786_),
    .Y(_08014_));
 sky130_fd_sc_hd__xnor2_2 _19940_ (.A(_13792_),
    .B(_08014_),
    .Y(\hash.CA1.p4[22] ));
 sky130_fd_sc_hd__and3_1 _19941_ (.A(_13777_),
    .B(_13782_),
    .C(_13787_),
    .X(_08015_));
 sky130_fd_sc_hd__nand2_1 _19942_ (.A(_13787_),
    .B(_13781_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand3_1 _19943_ (.A(_13782_),
    .B(_13787_),
    .C(_13776_),
    .Y(_08017_));
 sky130_fd_sc_hd__nand2_1 _19944_ (.A(_08016_),
    .B(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__a211o_1 _19945_ (.A1(_08002_),
    .A2(_08015_),
    .B1(_08018_),
    .C1(_13786_),
    .X(_08019_));
 sky130_fd_sc_hd__a21o_4 _19946_ (.A1(_13792_),
    .A2(_08019_),
    .B1(_13791_),
    .X(_08020_));
 sky130_fd_sc_hd__xor2_2 _19947_ (.A(_13798_),
    .B(_08020_),
    .X(\hash.CA1.p4[23] ));
 sky130_fd_sc_hd__inv_1 _19948_ (.A(_12464_),
    .Y(_13802_));
 sky130_fd_sc_hd__a21o_4 _19949_ (.A1(_13798_),
    .A2(_13791_),
    .B1(_13797_),
    .X(_08021_));
 sky130_fd_sc_hd__nand2_2 _19950_ (.A(_13792_),
    .B(_13798_),
    .Y(_08022_));
 sky130_fd_sc_hd__nor2_1 _19951_ (.A(_13787_),
    .B(_13786_),
    .Y(_08023_));
 sky130_fd_sc_hd__o21bai_1 _19952_ (.A1(_08022_),
    .A2(_08023_),
    .B1_N(_08021_),
    .Y(_08024_));
 sky130_fd_sc_hd__o41ai_2 _19953_ (.A1(_13781_),
    .A2(_13786_),
    .A3(_08006_),
    .A4(_08021_),
    .B1(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__xnor2_2 _19954_ (.A(_13805_),
    .B(_08025_),
    .Y(\hash.CA1.p4[24] ));
 sky130_fd_sc_hd__inv_1 _19955_ (.A(_12469_),
    .Y(_13809_));
 sky130_fd_sc_hd__clkinvlp_4 _19956_ (.A(_13812_),
    .Y(_08026_));
 sky130_fd_sc_hd__a21oi_1 _19957_ (.A1(_13805_),
    .A2(_13797_),
    .B1(_13804_),
    .Y(_08027_));
 sky130_fd_sc_hd__nand3_1 _19958_ (.A(_13798_),
    .B(_13805_),
    .C(_08020_),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_1 _19959_ (.A(_08027_),
    .B(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__xnor2_2 _19960_ (.A(_08026_),
    .B(_08029_),
    .Y(\hash.CA1.p4[25] ));
 sky130_fd_sc_hd__inv_1 _19961_ (.A(_12474_),
    .Y(_13816_));
 sky130_fd_sc_hd__nor2_1 _19962_ (.A(_08014_),
    .B(_08022_),
    .Y(_08030_));
 sky130_fd_sc_hd__a21oi_1 _19963_ (.A1(_13805_),
    .A2(_08021_),
    .B1(_13804_),
    .Y(_08031_));
 sky130_fd_sc_hd__o21bai_2 _19964_ (.A1(_08026_),
    .A2(_08031_),
    .B1_N(_13811_),
    .Y(_08032_));
 sky130_fd_sc_hd__a31oi_1 _19965_ (.A1(_13805_),
    .A2(_13812_),
    .A3(_08030_),
    .B1(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__xnor2_2 _19966_ (.A(_13819_),
    .B(_08033_),
    .Y(\hash.CA1.p4[26] ));
 sky130_fd_sc_hd__clkinv_1 _19967_ (.A(_12479_),
    .Y(_13823_));
 sky130_fd_sc_hd__inv_4 _19968_ (.A(_13826_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand2_2 _19969_ (.A(_13798_),
    .B(_08020_),
    .Y(_08035_));
 sky130_fd_sc_hd__nand3_2 _19970_ (.A(_13805_),
    .B(_13812_),
    .C(_13819_),
    .Y(_08036_));
 sky130_fd_sc_hd__o21bai_1 _19971_ (.A1(_08026_),
    .A2(_08027_),
    .B1_N(_13811_),
    .Y(_08037_));
 sky130_fd_sc_hd__a21oi_2 _19972_ (.A1(_13819_),
    .A2(_08037_),
    .B1(_13818_),
    .Y(_08038_));
 sky130_fd_sc_hd__o21ai_4 _19973_ (.A1(_08035_),
    .A2(_08036_),
    .B1(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__xnor2_4 _19974_ (.A(_08034_),
    .B(_08039_),
    .Y(\hash.CA1.p4[27] ));
 sky130_fd_sc_hd__clkinv_1 _19975_ (.A(_12484_),
    .Y(_13830_));
 sky130_fd_sc_hd__a21o_1 _19976_ (.A1(_13812_),
    .A2(_13804_),
    .B1(_13811_),
    .X(_08040_));
 sky130_fd_sc_hd__a21oi_1 _19977_ (.A1(_13819_),
    .A2(_08040_),
    .B1(_13818_),
    .Y(_08041_));
 sky130_fd_sc_hd__o21ai_0 _19978_ (.A1(_08025_),
    .A2(_08036_),
    .B1(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__a21oi_2 _19979_ (.A1(_13826_),
    .A2(_08042_),
    .B1(_13825_),
    .Y(_08043_));
 sky130_fd_sc_hd__xnor2_4 _19980_ (.A(_13833_),
    .B(_08043_),
    .Y(\hash.CA1.p4[28] ));
 sky130_fd_sc_hd__clkinv_1 _19981_ (.A(_12489_),
    .Y(_13837_));
 sky130_fd_sc_hd__a21o_1 _19982_ (.A1(_13826_),
    .A2(_08039_),
    .B1(_13825_),
    .X(_08044_));
 sky130_fd_sc_hd__a21oi_2 _19983_ (.A1(_13833_),
    .A2(_08044_),
    .B1(_13832_),
    .Y(_08045_));
 sky130_fd_sc_hd__xnor2_4 _19984_ (.A(_13839_),
    .B(_08045_),
    .Y(\hash.CA1.p4[29] ));
 sky130_fd_sc_hd__a21oi_1 _19985_ (.A1(_13819_),
    .A2(_08032_),
    .B1(_13818_),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_1 _19986_ (.A(_08034_),
    .B(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__o21a_1 _19987_ (.A1(_13825_),
    .A2(_08047_),
    .B1(_13833_),
    .X(_08048_));
 sky130_fd_sc_hd__o21ai_2 _19988_ (.A1(_13832_),
    .A2(_08048_),
    .B1(_13839_),
    .Y(_08049_));
 sky130_fd_sc_hd__nand2_1 _19989_ (.A(_13833_),
    .B(_13839_),
    .Y(_08050_));
 sky130_fd_sc_hd__or3_4 _19990_ (.A(_08034_),
    .B(_08036_),
    .C(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__nor2_1 _19991_ (.A(_08022_),
    .B(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__nand2b_1 _19992_ (.A_N(_13786_),
    .B(_08016_),
    .Y(_08053_));
 sky130_fd_sc_hd__a21oi_1 _19993_ (.A1(_08052_),
    .A2(_08053_),
    .B1(_13838_),
    .Y(_08054_));
 sky130_fd_sc_hd__nand3_1 _19994_ (.A(_13787_),
    .B(_08006_),
    .C(_08052_),
    .Y(_08055_));
 sky130_fd_sc_hd__nand3_2 _19995_ (.A(_08049_),
    .B(_08054_),
    .C(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__xor2_4 _19996_ (.A(_13844_),
    .B(_08056_),
    .X(\hash.CA1.p4[30] ));
 sky130_fd_sc_hd__xnor2_1 _19997_ (.A(\hash.CA1.S1.X[6] ),
    .B(_06575_),
    .Y(_08057_));
 sky130_fd_sc_hd__xnor2_2 _19998_ (.A(_08057_),
    .B(_06683_),
    .Y(_13861_));
 sky130_fd_sc_hd__xor2_1 _19999_ (.A(\hash.CA1.S1.X[7] ),
    .B(_06581_),
    .X(_08058_));
 sky130_fd_sc_hd__xnor2_2 _20000_ (.A(_06689_),
    .B(_08058_),
    .Y(_12501_));
 sky130_fd_sc_hd__xnor2_1 _20001_ (.A(_06552_),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_08059_));
 sky130_fd_sc_hd__xnor2_1 _20002_ (.A(_06699_),
    .B(_08059_),
    .Y(_13869_));
 sky130_fd_sc_hd__xnor2_1 _20003_ (.A(_06559_),
    .B(_06597_),
    .Y(_08060_));
 sky130_fd_sc_hd__xnor2_2 _20004_ (.A(_06707_),
    .B(_08060_),
    .Y(_13877_));
 sky130_fd_sc_hd__xnor2_1 _20005_ (.A(\hash.CA1.S1.X[10] ),
    .B(_06610_),
    .Y(_08061_));
 sky130_fd_sc_hd__xnor2_1 _20006_ (.A(\hash.CA1.S1.X[29] ),
    .B(_08061_),
    .Y(_13886_));
 sky130_fd_sc_hd__inv_1 _20007_ (.A(_12516_),
    .Y(_13890_));
 sky130_fd_sc_hd__nand3b_1 _20008_ (.A_N(_13884_),
    .B(_06942_),
    .C(_06943_),
    .Y(_08062_));
 sky130_fd_sc_hd__xor2_2 _20009_ (.A(_13895_),
    .B(_08062_),
    .X(_12524_));
 sky130_fd_sc_hd__xnor2_1 _20010_ (.A(_06575_),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_08063_));
 sky130_fd_sc_hd__xnor2_2 _20011_ (.A(\hash.CA1.S1.X[30] ),
    .B(_08063_),
    .Y(_13896_));
 sky130_fd_sc_hd__inv_1 _20012_ (.A(_12521_),
    .Y(_13900_));
 sky130_fd_sc_hd__xnor2_1 _20013_ (.A(_06581_),
    .B(_06624_),
    .Y(_08064_));
 sky130_fd_sc_hd__xnor2_2 _20014_ (.A(_08064_),
    .B(\hash.CA1.S1.X[31] ),
    .Y(_13905_));
 sky130_fd_sc_hd__nor2_1 _20015_ (.A(\hash.CA1.S1.X[0] ),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_08065_));
 sky130_fd_sc_hd__a21oi_1 _20016_ (.A1(_13445_),
    .A2(\hash.CA1.S1.X[13] ),
    .B1(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__xnor2_1 _20017_ (.A(_06634_),
    .B(_08066_),
    .Y(_13913_));
 sky130_fd_sc_hd__nor2_1 _20018_ (.A(\hash.CA1.S1.X[1] ),
    .B(_06642_),
    .Y(_08067_));
 sky130_fd_sc_hd__a21oi_1 _20019_ (.A1(_12365_),
    .A2(_06642_),
    .B1(_08067_),
    .Y(_08068_));
 sky130_fd_sc_hd__xnor2_1 _20020_ (.A(\hash.CA1.S1.X[14] ),
    .B(_08068_),
    .Y(_13921_));
 sky130_fd_sc_hd__xnor2_1 _20021_ (.A(\hash.CA1.S1.X[2] ),
    .B(_06610_),
    .Y(_08069_));
 sky130_fd_sc_hd__xnor2_1 _20022_ (.A(\hash.CA1.S1.X[20] ),
    .B(_08069_),
    .Y(_13930_));
 sky130_fd_sc_hd__xnor2_1 _20023_ (.A(_13933_),
    .B(_07117_),
    .Y(_12543_));
 sky130_fd_sc_hd__clkinv_1 _20024_ (.A(_12541_),
    .Y(_13934_));
 sky130_fd_sc_hd__xnor2_1 _20025_ (.A(\hash.CA1.S1.X[3] ),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_08070_));
 sky130_fd_sc_hd__xnor2_1 _20026_ (.A(\hash.CA1.S1.X[21] ),
    .B(_08070_),
    .Y(_13939_));
 sky130_fd_sc_hd__xnor2_1 _20027_ (.A(_06524_),
    .B(_06624_),
    .Y(_08071_));
 sky130_fd_sc_hd__xnor2_1 _20028_ (.A(\hash.CA1.S1.X[22] ),
    .B(_08071_),
    .Y(_13948_));
 sky130_fd_sc_hd__clkinv_1 _20029_ (.A(_12551_),
    .Y(_13952_));
 sky130_fd_sc_hd__a21oi_1 _20030_ (.A1(_06956_),
    .A2(_06971_),
    .B1(_06974_),
    .Y(_08072_));
 sky130_fd_sc_hd__o21ai_1 _20031_ (.A1(_06969_),
    .A2(_08072_),
    .B1(_07002_),
    .Y(_08073_));
 sky130_fd_sc_hd__xnor2_2 _20032_ (.A(_06982_),
    .B(_08073_),
    .Y(_12559_));
 sky130_fd_sc_hd__xnor2_1 _20033_ (.A(_06531_),
    .B(_06634_),
    .Y(_08074_));
 sky130_fd_sc_hd__xnor2_1 _20034_ (.A(\hash.CA1.S1.X[23] ),
    .B(_08074_),
    .Y(_13958_));
 sky130_fd_sc_hd__xnor2_1 _20035_ (.A(_13961_),
    .B(_07119_),
    .Y(_12558_));
 sky130_fd_sc_hd__clkinv_1 _20036_ (.A(_12556_),
    .Y(_13962_));
 sky130_fd_sc_hd__a21oi_1 _20037_ (.A1(_07001_),
    .A2(_07003_),
    .B1(_13956_),
    .Y(_08075_));
 sky130_fd_sc_hd__xnor2_2 _20038_ (.A(_13966_),
    .B(_08075_),
    .Y(_12564_));
 sky130_fd_sc_hd__xnor2_1 _20039_ (.A(\hash.CA1.S1.X[6] ),
    .B(_06642_),
    .Y(_08076_));
 sky130_fd_sc_hd__xnor2_1 _20040_ (.A(_06673_),
    .B(_08076_),
    .Y(_13967_));
 sky130_fd_sc_hd__o31a_1 _20041_ (.A1(_13970_),
    .A2(_06989_),
    .A3(_07120_),
    .B1(_07012_),
    .X(_12563_));
 sky130_fd_sc_hd__xnor2_1 _20042_ (.A(\hash.CA1.S1.X[7] ),
    .B(\hash.CA1.S1.X[20] ),
    .Y(_08077_));
 sky130_fd_sc_hd__xnor2_1 _20043_ (.A(_06683_),
    .B(_08077_),
    .Y(_13975_));
 sky130_fd_sc_hd__xnor2_1 _20044_ (.A(_06552_),
    .B(\hash.CA1.S1.X[21] ),
    .Y(_08078_));
 sky130_fd_sc_hd__xnor2_1 _20045_ (.A(_06689_),
    .B(_08078_),
    .Y(_13984_));
 sky130_fd_sc_hd__clkinv_1 _20046_ (.A(_12571_),
    .Y(_13988_));
 sky130_fd_sc_hd__a21oi_1 _20047_ (.A1(_13983_),
    .A2(_07024_),
    .B1(_13982_),
    .Y(_08079_));
 sky130_fd_sc_hd__xnor2_2 _20048_ (.A(_13993_),
    .B(_08079_),
    .Y(_12579_));
 sky130_fd_sc_hd__xnor2_1 _20049_ (.A(\hash.CA1.S1.X[9] ),
    .B(\hash.CA1.S1.X[22] ),
    .Y(_08080_));
 sky130_fd_sc_hd__xnor2_1 _20050_ (.A(_06699_),
    .B(_08080_),
    .Y(_13994_));
 sky130_fd_sc_hd__xnor2_1 _20051_ (.A(_13997_),
    .B(_07055_),
    .Y(_12578_));
 sky130_fd_sc_hd__clkinv_1 _20052_ (.A(_12576_),
    .Y(_13998_));
 sky130_fd_sc_hd__a31oi_1 _20053_ (.A1(_13983_),
    .A2(_13993_),
    .A3(_07008_),
    .B1(_07019_),
    .Y(_08081_));
 sky130_fd_sc_hd__xnor2_2 _20054_ (.A(_14002_),
    .B(_08081_),
    .Y(_12584_));
 sky130_fd_sc_hd__xnor2_1 _20055_ (.A(\hash.CA1.S1.X[10] ),
    .B(\hash.CA1.S1.X[23] ),
    .Y(_08082_));
 sky130_fd_sc_hd__xnor2_1 _20056_ (.A(_06707_),
    .B(_08082_),
    .Y(_14003_));
 sky130_fd_sc_hd__a21oi_1 _20057_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07041_),
    .Y(_12583_));
 sky130_fd_sc_hd__a31o_1 _20058_ (.A1(_13983_),
    .A2(_13993_),
    .A3(_07024_),
    .B1(_07019_),
    .X(_08083_));
 sky130_fd_sc_hd__a21oi_2 _20059_ (.A1(_14002_),
    .A2(_08083_),
    .B1(_14001_),
    .Y(_08084_));
 sky130_fd_sc_hd__xnor2_2 _20060_ (.A(_14010_),
    .B(_08084_),
    .Y(_12589_));
 sky130_fd_sc_hd__xnor3_1 _20061_ (.A(_06575_),
    .B(_06673_),
    .C(\hash.CA1.S1.X[29] ),
    .X(_14011_));
 sky130_fd_sc_hd__xnor2_1 _20062_ (.A(_14014_),
    .B(_07123_),
    .Y(_12588_));
 sky130_fd_sc_hd__xnor2_2 _20063_ (.A(_14018_),
    .B(_07030_),
    .Y(_12594_));
 sky130_fd_sc_hd__xnor2_1 _20064_ (.A(\hash.CA1.S1.X[12] ),
    .B(_06683_),
    .Y(_08085_));
 sky130_fd_sc_hd__xnor2_1 _20065_ (.A(net1046),
    .B(_08085_),
    .Y(_14019_));
 sky130_fd_sc_hd__xnor2_1 _20066_ (.A(_14022_),
    .B(_07125_),
    .Y(_12593_));
 sky130_fd_sc_hd__xnor2_1 _20067_ (.A(\hash.CA1.S1.X[13] ),
    .B(_06689_),
    .Y(_08086_));
 sky130_fd_sc_hd__xnor2_1 _20068_ (.A(\hash.CA1.S1.X[31] ),
    .B(_08086_),
    .Y(_14027_));
 sky130_fd_sc_hd__xnor2_1 _20069_ (.A(_14030_),
    .B(_07128_),
    .Y(_12598_));
 sky130_fd_sc_hd__nor2_1 _20070_ (.A(\hash.CA1.S1.X[0] ),
    .B(_06699_),
    .Y(_08087_));
 sky130_fd_sc_hd__a21oi_1 _20071_ (.A1(_13445_),
    .A2(_06699_),
    .B1(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__xnor2_1 _20072_ (.A(_06597_),
    .B(_08088_),
    .Y(_14035_));
 sky130_fd_sc_hd__mux2i_1 _20073_ (.A0(_12365_),
    .A1(_13854_),
    .S(_06707_),
    .Y(_08089_));
 sky130_fd_sc_hd__xnor2_1 _20074_ (.A(_06610_),
    .B(_08089_),
    .Y(_14044_));
 sky130_fd_sc_hd__inv_1 _20075_ (.A(_12606_),
    .Y(_14048_));
 sky130_fd_sc_hd__xnor2_1 _20076_ (.A(_06514_),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_08090_));
 sky130_fd_sc_hd__xnor2_2 _20077_ (.A(_06712_),
    .B(_08090_),
    .Y(_14054_));
 sky130_fd_sc_hd__inv_1 _20078_ (.A(_12611_),
    .Y(_14058_));
 sky130_fd_sc_hd__xor2_1 _20079_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06624_),
    .X(_08091_));
 sky130_fd_sc_hd__xnor2_1 _20080_ (.A(net1045),
    .B(_08091_),
    .Y(_14064_));
 sky130_fd_sc_hd__inv_1 _20081_ (.A(_12616_),
    .Y(_14068_));
 sky130_fd_sc_hd__xnor2_1 _20082_ (.A(_06524_),
    .B(_06634_),
    .Y(_08092_));
 sky130_fd_sc_hd__xnor2_2 _20083_ (.A(\hash.CA1.S1.X[31] ),
    .B(_08092_),
    .Y(_14074_));
 sky130_fd_sc_hd__inv_1 _20084_ (.A(_12621_),
    .Y(_14078_));
 sky130_fd_sc_hd__nor2_1 _20085_ (.A(_14072_),
    .B(_07093_),
    .Y(_08093_));
 sky130_fd_sc_hd__xnor2_2 _20086_ (.A(_14083_),
    .B(_08093_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand2_8 _20087_ (.A(_06528_),
    .B(_06530_),
    .Y(_08094_));
 sky130_fd_sc_hd__xnor2_1 _20088_ (.A(_13445_),
    .B(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__and2_4 _20089_ (.A(_06002_),
    .B(_08095_),
    .X(_08096_));
 sky130_fd_sc_hd__xnor2_2 _20090_ (.A(_06642_),
    .B(_08096_),
    .Y(_14084_));
 sky130_fd_sc_hd__xor2_1 _20091_ (.A(_14087_),
    .B(_07129_),
    .X(_12628_));
 sky130_fd_sc_hd__inv_1 _20092_ (.A(_12626_),
    .Y(_14088_));
 sky130_fd_sc_hd__mux2i_1 _20093_ (.A0(_12365_),
    .A1(_13854_),
    .S(\hash.CA1.S1.X[6] ),
    .Y(_08097_));
 sky130_fd_sc_hd__xnor2_2 _20094_ (.A(\hash.CA1.S1.X[20] ),
    .B(_08097_),
    .Y(_14093_));
 sky130_fd_sc_hd__xnor2_1 _20095_ (.A(\hash.CA1.S1.X[2] ),
    .B(\hash.CA1.S1.X[7] ),
    .Y(_08098_));
 sky130_fd_sc_hd__xnor2_1 _20096_ (.A(\hash.CA1.S1.X[21] ),
    .B(_08098_),
    .Y(_14102_));
 sky130_fd_sc_hd__inv_1 _20097_ (.A(_12636_),
    .Y(_14106_));
 sky130_fd_sc_hd__nor3_2 _20098_ (.A(_14072_),
    .B(_14082_),
    .C(_14091_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand2_1 _20099_ (.A(_14101_),
    .B(_07095_),
    .Y(_08100_));
 sky130_fd_sc_hd__a21oi_4 _20100_ (.A1(_07084_),
    .A2(_08099_),
    .B1(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__nor2_1 _20101_ (.A(_14100_),
    .B(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__xnor2_2 _20102_ (.A(_14111_),
    .B(_08102_),
    .Y(_12644_));
 sky130_fd_sc_hd__xnor2_1 _20103_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06552_),
    .Y(_08103_));
 sky130_fd_sc_hd__xnor2_1 _20104_ (.A(\hash.CA1.S1.X[22] ),
    .B(_08103_),
    .Y(_14112_));
 sky130_fd_sc_hd__xnor2_1 _20105_ (.A(_14115_),
    .B(_07134_),
    .Y(_12643_));
 sky130_fd_sc_hd__inv_1 _20106_ (.A(_12641_),
    .Y(_14116_));
 sky130_fd_sc_hd__or3_4 _20107_ (.A(_07107_),
    .B(_07109_),
    .C(_07110_),
    .X(_12870_));
 sky130_fd_sc_hd__xnor2_1 _20108_ (.A(_06524_),
    .B(_06559_),
    .Y(_08104_));
 sky130_fd_sc_hd__xnor2_1 _20109_ (.A(\hash.CA1.S1.X[23] ),
    .B(_08104_),
    .Y(_14121_));
 sky130_fd_sc_hd__inv_1 _20110_ (.A(_12663_),
    .Y(_14128_));
 sky130_fd_sc_hd__inv_1 _20111_ (.A(_12672_),
    .Y(_14132_));
 sky130_fd_sc_hd__clkinv_1 _20112_ (.A(_12677_),
    .Y(_14136_));
 sky130_fd_sc_hd__clkinv_1 _20113_ (.A(_12682_),
    .Y(_14140_));
 sky130_fd_sc_hd__clkinv_1 _20114_ (.A(_12689_),
    .Y(_14144_));
 sky130_fd_sc_hd__clkinv_1 _20115_ (.A(_12698_),
    .Y(_14148_));
 sky130_fd_sc_hd__inv_1 _20116_ (.A(_12706_),
    .Y(_14152_));
 sky130_fd_sc_hd__clkinv_1 _20117_ (.A(_12709_),
    .Y(_12718_));
 sky130_fd_sc_hd__inv_1 _20118_ (.A(_12711_),
    .Y(_14156_));
 sky130_fd_sc_hd__inv_2 _20119_ (.A(_12716_),
    .Y(_12726_));
 sky130_fd_sc_hd__inv_1 _20120_ (.A(_12753_),
    .Y(_12762_));
 sky130_fd_sc_hd__inv_1 _20121_ (.A(_12760_),
    .Y(_12770_));
 sky130_fd_sc_hd__inv_2 _20122_ (.A(_12795_),
    .Y(_12806_));
 sky130_fd_sc_hd__inv_1 _20123_ (.A(_12811_),
    .Y(_12822_));
 sky130_fd_sc_hd__inv_1 _20124_ (.A(_12827_),
    .Y(_12838_));
 sky130_fd_sc_hd__inv_2 _20125_ (.A(_06782_),
    .Y(_12842_));
 sky130_fd_sc_hd__a21oi_1 _20126_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_13235_),
    .B1(_12922_),
    .Y(_08105_));
 sky130_fd_sc_hd__nor2_1 _20127_ (.A(\hash.CA2.a_dash[0] ),
    .B(_13235_),
    .Y(_08106_));
 sky130_fd_sc_hd__o21ai_0 _20128_ (.A1(_08105_),
    .A2(_08106_),
    .B1(_06002_),
    .Y(_14202_));
 sky130_fd_sc_hd__clkinvlp_4 _20129_ (.A(\count_hash2[2] ),
    .Y(_12900_));
 sky130_fd_sc_hd__clkinvlp_4 _20130_ (.A(\count_hash1[2] ),
    .Y(_12910_));
 sky130_fd_sc_hd__inv_1 _20131_ (.A(_11583_),
    .Y(_12984_));
 sky130_fd_sc_hd__inv_1 _20132_ (.A(_11591_),
    .Y(_12987_));
 sky130_fd_sc_hd__inv_1 _20133_ (.A(_11599_),
    .Y(_12991_));
 sky130_fd_sc_hd__inv_1 _20134_ (.A(_11610_),
    .Y(_12995_));
 sky130_fd_sc_hd__inv_1 _20135_ (.A(_11618_),
    .Y(_12999_));
 sky130_fd_sc_hd__inv_1 _20136_ (.A(_11626_),
    .Y(_13003_));
 sky130_fd_sc_hd__inv_1 _20137_ (.A(_11634_),
    .Y(_13007_));
 sky130_fd_sc_hd__inv_1 _20138_ (.A(_11642_),
    .Y(_13011_));
 sky130_fd_sc_hd__inv_1 _20139_ (.A(_11650_),
    .Y(_13015_));
 sky130_fd_sc_hd__inv_1 _20140_ (.A(_11658_),
    .Y(_13019_));
 sky130_fd_sc_hd__inv_1 _20141_ (.A(_11666_),
    .Y(_13023_));
 sky130_fd_sc_hd__inv_1 _20142_ (.A(_11674_),
    .Y(_13027_));
 sky130_fd_sc_hd__inv_1 _20143_ (.A(_11682_),
    .Y(_13031_));
 sky130_fd_sc_hd__inv_1 _20144_ (.A(_11690_),
    .Y(_13035_));
 sky130_fd_sc_hd__inv_1 _20145_ (.A(_11698_),
    .Y(_13039_));
 sky130_fd_sc_hd__inv_1 _20146_ (.A(_11706_),
    .Y(_13043_));
 sky130_fd_sc_hd__inv_1 _20147_ (.A(_11714_),
    .Y(_13047_));
 sky130_fd_sc_hd__inv_1 _20148_ (.A(_11722_),
    .Y(_13051_));
 sky130_fd_sc_hd__inv_1 _20149_ (.A(_11730_),
    .Y(_13055_));
 sky130_fd_sc_hd__inv_1 _20150_ (.A(_11738_),
    .Y(_13059_));
 sky130_fd_sc_hd__inv_1 _20151_ (.A(_11746_),
    .Y(_13063_));
 sky130_fd_sc_hd__inv_1 _20152_ (.A(_11754_),
    .Y(_13067_));
 sky130_fd_sc_hd__inv_1 _20153_ (.A(_11762_),
    .Y(_13071_));
 sky130_fd_sc_hd__inv_1 _20154_ (.A(_11770_),
    .Y(_13075_));
 sky130_fd_sc_hd__inv_1 _20155_ (.A(_11778_),
    .Y(_13079_));
 sky130_fd_sc_hd__inv_1 _20156_ (.A(_11786_),
    .Y(_13083_));
 sky130_fd_sc_hd__inv_2 _20157_ (.A(_11794_),
    .Y(_13087_));
 sky130_fd_sc_hd__inv_1 _20158_ (.A(_11802_),
    .Y(_13091_));
 sky130_fd_sc_hd__inv_1 _20159_ (.A(_11810_),
    .Y(_13095_));
 sky130_fd_sc_hd__inv_2 _20160_ (.A(_11818_),
    .Y(_13099_));
 sky130_fd_sc_hd__inv_1 _20161_ (.A(_11826_),
    .Y(_13103_));
 sky130_fd_sc_hd__inv_1 _20162_ (.A(_11831_),
    .Y(_13107_));
 sky130_fd_sc_hd__clkinvlp_2 _20163_ (.A(_11839_),
    .Y(_13110_));
 sky130_fd_sc_hd__inv_1 _20164_ (.A(_11847_),
    .Y(_13114_));
 sky130_fd_sc_hd__inv_1 _20165_ (.A(_11858_),
    .Y(_13118_));
 sky130_fd_sc_hd__inv_1 _20166_ (.A(_11866_),
    .Y(_13122_));
 sky130_fd_sc_hd__inv_1 _20167_ (.A(_11874_),
    .Y(_13126_));
 sky130_fd_sc_hd__inv_1 _20168_ (.A(_11882_),
    .Y(_13130_));
 sky130_fd_sc_hd__inv_1 _20169_ (.A(_11890_),
    .Y(_13134_));
 sky130_fd_sc_hd__inv_1 _20170_ (.A(_11898_),
    .Y(_13138_));
 sky130_fd_sc_hd__clkinv_1 _20171_ (.A(_11906_),
    .Y(_13142_));
 sky130_fd_sc_hd__inv_1 _20172_ (.A(_11914_),
    .Y(_13146_));
 sky130_fd_sc_hd__inv_2 _20173_ (.A(_11922_),
    .Y(_13150_));
 sky130_fd_sc_hd__inv_1 _20174_ (.A(_11930_),
    .Y(_13154_));
 sky130_fd_sc_hd__inv_1 _20175_ (.A(_11938_),
    .Y(_13158_));
 sky130_fd_sc_hd__inv_1 _20176_ (.A(_11946_),
    .Y(_13162_));
 sky130_fd_sc_hd__inv_1 _20177_ (.A(_11954_),
    .Y(_13166_));
 sky130_fd_sc_hd__inv_1 _20178_ (.A(_11962_),
    .Y(_13170_));
 sky130_fd_sc_hd__inv_1 _20179_ (.A(_11970_),
    .Y(_13174_));
 sky130_fd_sc_hd__clkinv_1 _20180_ (.A(_11978_),
    .Y(_13178_));
 sky130_fd_sc_hd__clkinv_1 _20181_ (.A(_11986_),
    .Y(_13182_));
 sky130_fd_sc_hd__inv_1 _20182_ (.A(_11994_),
    .Y(_13186_));
 sky130_fd_sc_hd__inv_1 _20183_ (.A(_12002_),
    .Y(_13190_));
 sky130_fd_sc_hd__inv_1 _20184_ (.A(_12010_),
    .Y(_13194_));
 sky130_fd_sc_hd__inv_1 _20185_ (.A(_12018_),
    .Y(_13198_));
 sky130_fd_sc_hd__inv_1 _20186_ (.A(_12026_),
    .Y(_13202_));
 sky130_fd_sc_hd__inv_1 _20187_ (.A(_12034_),
    .Y(_13206_));
 sky130_fd_sc_hd__inv_1 _20188_ (.A(_12042_),
    .Y(_13210_));
 sky130_fd_sc_hd__inv_1 _20189_ (.A(_12050_),
    .Y(_13214_));
 sky130_fd_sc_hd__inv_1 _20190_ (.A(_12058_),
    .Y(_13218_));
 sky130_fd_sc_hd__inv_1 _20191_ (.A(_12066_),
    .Y(_13222_));
 sky130_fd_sc_hd__inv_1 _20192_ (.A(_12074_),
    .Y(_13226_));
 sky130_fd_sc_hd__inv_1 _20193_ (.A(_12079_),
    .Y(_13233_));
 sky130_fd_sc_hd__inv_1 _20194_ (.A(_12091_),
    .Y(_12093_));
 sky130_fd_sc_hd__xnor2_1 _20195_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[27] ),
    .Y(_08107_));
 sky130_fd_sc_hd__xnor2_2 _20196_ (.A(\hash.CA2.S1.X[13] ),
    .B(_08107_),
    .Y(_13243_));
 sky130_fd_sc_hd__inv_1 _20197_ (.A(_12100_),
    .Y(_12102_));
 sky130_fd_sc_hd__xnor2_1 _20198_ (.A(\hash.CA2.S1.X[9] ),
    .B(\hash.CA2.S1.X[28] ),
    .Y(_08108_));
 sky130_fd_sc_hd__xnor2_2 _20199_ (.A(\hash.CA2.S1.X[14] ),
    .B(_08108_),
    .Y(_13250_));
 sky130_fd_sc_hd__inv_1 _20200_ (.A(_12114_),
    .Y(_12116_));
 sky130_fd_sc_hd__xnor2_2 _20201_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA2.S1.X[29] ),
    .Y(_08109_));
 sky130_fd_sc_hd__xnor2_2 _20202_ (.A(\hash.CA2.S1.X[15] ),
    .B(_08109_),
    .Y(_13257_));
 sky130_fd_sc_hd__inv_1 _20203_ (.A(_12123_),
    .Y(_12125_));
 sky130_fd_sc_hd__xnor2_1 _20204_ (.A(\hash.CA2.S1.X[16] ),
    .B(\hash.CA2.S1.X[30] ),
    .Y(_08110_));
 sky130_fd_sc_hd__xnor2_1 _20205_ (.A(\hash.CA2.S1.X[11] ),
    .B(_08110_),
    .Y(_13264_));
 sky130_fd_sc_hd__inv_1 _20206_ (.A(_12132_),
    .Y(_12134_));
 sky130_fd_sc_hd__xnor2_1 _20207_ (.A(\hash.CA2.S1.X[12] ),
    .B(\hash.CA2.S1.X[17] ),
    .Y(_08111_));
 sky130_fd_sc_hd__xnor2_1 _20208_ (.A(\hash.CA2.S1.X[31] ),
    .B(_08111_),
    .Y(_13271_));
 sky130_fd_sc_hd__inv_1 _20209_ (.A(_12141_),
    .Y(_12143_));
 sky130_fd_sc_hd__xnor2_1 _20210_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA2.S1.X[18] ),
    .Y(_08112_));
 sky130_fd_sc_hd__xnor2_1 _20211_ (.A(\hash.CA2.S1.X[0] ),
    .B(_08112_),
    .Y(_13278_));
 sky130_fd_sc_hd__inv_1 _20212_ (.A(_12150_),
    .Y(_12152_));
 sky130_fd_sc_hd__xnor2_1 _20213_ (.A(\hash.CA2.S1.X[14] ),
    .B(\hash.CA2.S1.X[19] ),
    .Y(_08113_));
 sky130_fd_sc_hd__xnor2_1 _20214_ (.A(\hash.CA2.S1.X[1] ),
    .B(_08113_),
    .Y(_13285_));
 sky130_fd_sc_hd__inv_2 _20215_ (.A(_12159_),
    .Y(_12161_));
 sky130_fd_sc_hd__xnor2_1 _20216_ (.A(\hash.CA2.S1.X[15] ),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08114_));
 sky130_fd_sc_hd__xnor2_1 _20217_ (.A(\hash.CA2.S1.X[2] ),
    .B(_08114_),
    .Y(_13292_));
 sky130_fd_sc_hd__inv_1 _20218_ (.A(_12168_),
    .Y(_12170_));
 sky130_fd_sc_hd__xnor2_1 _20219_ (.A(\hash.CA2.S1.X[16] ),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08115_));
 sky130_fd_sc_hd__xnor2_1 _20220_ (.A(\hash.CA2.S1.X[3] ),
    .B(_08115_),
    .Y(_13299_));
 sky130_fd_sc_hd__inv_1 _20221_ (.A(_12177_),
    .Y(_12179_));
 sky130_fd_sc_hd__xnor2_1 _20222_ (.A(\hash.CA2.S1.X[17] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08116_));
 sky130_fd_sc_hd__xnor2_1 _20223_ (.A(\hash.CA2.S1.X[4] ),
    .B(_08116_),
    .Y(_13306_));
 sky130_fd_sc_hd__inv_1 _20224_ (.A(_12186_),
    .Y(_12188_));
 sky130_fd_sc_hd__xnor2_1 _20225_ (.A(\hash.CA2.S1.X[18] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08117_));
 sky130_fd_sc_hd__xnor2_1 _20226_ (.A(\hash.CA2.S1.X[5] ),
    .B(_08117_),
    .Y(_13313_));
 sky130_fd_sc_hd__inv_1 _20227_ (.A(_12195_),
    .Y(_12197_));
 sky130_fd_sc_hd__xnor2_1 _20228_ (.A(\hash.CA2.S1.X[19] ),
    .B(\hash.CA2.S1.X[24] ),
    .Y(_08118_));
 sky130_fd_sc_hd__xnor2_1 _20229_ (.A(\hash.CA2.S1.X[6] ),
    .B(_08118_),
    .Y(_13320_));
 sky130_fd_sc_hd__inv_1 _20230_ (.A(_12204_),
    .Y(_12206_));
 sky130_fd_sc_hd__xnor2_1 _20231_ (.A(net1062),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08119_));
 sky130_fd_sc_hd__xnor2_1 _20232_ (.A(net1072),
    .B(_08119_),
    .Y(_13327_));
 sky130_fd_sc_hd__inv_1 _20233_ (.A(_12213_),
    .Y(_12215_));
 sky130_fd_sc_hd__xnor2_1 _20234_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08120_));
 sky130_fd_sc_hd__xnor2_1 _20235_ (.A(net1063),
    .B(_08120_),
    .Y(_13334_));
 sky130_fd_sc_hd__inv_1 _20236_ (.A(_12222_),
    .Y(_12224_));
 sky130_fd_sc_hd__xnor2_1 _20237_ (.A(\hash.CA2.S1.X[9] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08121_));
 sky130_fd_sc_hd__xnor2_1 _20238_ (.A(\hash.CA2.S1.X[27] ),
    .B(_08121_),
    .Y(_13341_));
 sky130_fd_sc_hd__inv_1 _20239_ (.A(_12231_),
    .Y(_12233_));
 sky130_fd_sc_hd__xnor2_1 _20240_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08122_));
 sky130_fd_sc_hd__xnor2_1 _20241_ (.A(\hash.CA2.S1.X[28] ),
    .B(_08122_),
    .Y(_13348_));
 sky130_fd_sc_hd__inv_1 _20242_ (.A(_12240_),
    .Y(_12242_));
 sky130_fd_sc_hd__xnor2_1 _20243_ (.A(\hash.CA2.S1.X[29] ),
    .B(\hash.CA2.S1.X[24] ),
    .Y(_08123_));
 sky130_fd_sc_hd__xnor2_1 _20244_ (.A(\hash.CA2.S1.X[11] ),
    .B(_08123_),
    .Y(_13355_));
 sky130_fd_sc_hd__inv_1 _20245_ (.A(_12249_),
    .Y(_12251_));
 sky130_fd_sc_hd__xnor2_1 _20246_ (.A(\hash.CA2.S1.X[12] ),
    .B(\hash.CA2.S1.X[30] ),
    .Y(_08124_));
 sky130_fd_sc_hd__xnor2_1 _20247_ (.A(\hash.CA2.S1.X[25] ),
    .B(_08124_),
    .Y(_13362_));
 sky130_fd_sc_hd__inv_1 _20248_ (.A(_12258_),
    .Y(_12260_));
 sky130_fd_sc_hd__xnor2_1 _20249_ (.A(\hash.CA2.S1.X[26] ),
    .B(\hash.CA2.S1.X[13] ),
    .Y(_08125_));
 sky130_fd_sc_hd__xnor2_1 _20250_ (.A(\hash.CA2.S1.X[31] ),
    .B(_08125_),
    .Y(_13369_));
 sky130_fd_sc_hd__inv_1 _20251_ (.A(_12267_),
    .Y(_12269_));
 sky130_fd_sc_hd__xnor2_1 _20252_ (.A(\hash.CA2.S1.X[27] ),
    .B(\hash.CA2.S1.X[14] ),
    .Y(_08126_));
 sky130_fd_sc_hd__xnor2_1 _20253_ (.A(\hash.CA2.S1.X[0] ),
    .B(_08126_),
    .Y(_13376_));
 sky130_fd_sc_hd__inv_1 _20254_ (.A(_12276_),
    .Y(_12278_));
 sky130_fd_sc_hd__xnor2_1 _20255_ (.A(\hash.CA2.S1.X[28] ),
    .B(\hash.CA2.S1.X[15] ),
    .Y(_08127_));
 sky130_fd_sc_hd__xnor2_1 _20256_ (.A(\hash.CA2.S1.X[1] ),
    .B(_08127_),
    .Y(_13383_));
 sky130_fd_sc_hd__inv_1 _20257_ (.A(_12285_),
    .Y(_12287_));
 sky130_fd_sc_hd__xnor2_1 _20258_ (.A(\hash.CA2.S1.X[29] ),
    .B(\hash.CA2.S1.X[16] ),
    .Y(_08128_));
 sky130_fd_sc_hd__xnor2_1 _20259_ (.A(\hash.CA2.S1.X[2] ),
    .B(_08128_),
    .Y(_13390_));
 sky130_fd_sc_hd__inv_1 _20260_ (.A(_12294_),
    .Y(_12296_));
 sky130_fd_sc_hd__xnor2_1 _20261_ (.A(\hash.CA2.S1.X[30] ),
    .B(\hash.CA2.S1.X[17] ),
    .Y(_08129_));
 sky130_fd_sc_hd__xnor2_1 _20262_ (.A(\hash.CA2.S1.X[3] ),
    .B(_08129_),
    .Y(_13397_));
 sky130_fd_sc_hd__inv_1 _20263_ (.A(_12303_),
    .Y(_12305_));
 sky130_fd_sc_hd__xnor2_1 _20264_ (.A(\hash.CA2.S1.X[4] ),
    .B(\hash.CA2.S1.X[18] ),
    .Y(_08130_));
 sky130_fd_sc_hd__xnor2_1 _20265_ (.A(\hash.CA2.S1.X[31] ),
    .B(_08130_),
    .Y(_13404_));
 sky130_fd_sc_hd__inv_1 _20266_ (.A(_12312_),
    .Y(_12314_));
 sky130_fd_sc_hd__xnor2_1 _20267_ (.A(\hash.CA2.S1.X[5] ),
    .B(\hash.CA2.S1.X[19] ),
    .Y(_08131_));
 sky130_fd_sc_hd__xnor2_1 _20268_ (.A(\hash.CA2.S1.X[0] ),
    .B(_08131_),
    .Y(_13411_));
 sky130_fd_sc_hd__inv_1 _20269_ (.A(_12321_),
    .Y(_12323_));
 sky130_fd_sc_hd__xnor2_1 _20270_ (.A(\hash.CA2.S1.X[1] ),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08132_));
 sky130_fd_sc_hd__xnor2_1 _20271_ (.A(\hash.CA2.S1.X[6] ),
    .B(_08132_),
    .Y(_13418_));
 sky130_fd_sc_hd__inv_1 _20272_ (.A(_12330_),
    .Y(_12332_));
 sky130_fd_sc_hd__xnor2_1 _20273_ (.A(\hash.CA2.S1.X[2] ),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08133_));
 sky130_fd_sc_hd__xnor2_1 _20274_ (.A(net1059),
    .B(_08133_),
    .Y(_13425_));
 sky130_fd_sc_hd__inv_1 _20275_ (.A(_12339_),
    .Y(_12341_));
 sky130_fd_sc_hd__xnor2_1 _20276_ (.A(\hash.CA2.S1.X[3] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08134_));
 sky130_fd_sc_hd__xnor2_1 _20277_ (.A(\hash.CA2.S1.X[8] ),
    .B(_08134_),
    .Y(_13432_));
 sky130_fd_sc_hd__inv_1 _20278_ (.A(_12348_),
    .Y(_12350_));
 sky130_fd_sc_hd__xnor2_1 _20279_ (.A(\hash.CA2.S1.X[4] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08135_));
 sky130_fd_sc_hd__xnor2_1 _20280_ (.A(\hash.CA2.S1.X[9] ),
    .B(_08135_),
    .Y(_13439_));
 sky130_fd_sc_hd__inv_1 _20281_ (.A(_12357_),
    .Y(_12359_));
 sky130_fd_sc_hd__inv_1 _20282_ (.A(_12087_),
    .Y(_12363_));
 sky130_fd_sc_hd__xnor2_1 _20283_ (.A(_13427_),
    .B(_04760_),
    .Y(_13428_));
 sky130_fd_sc_hd__xor2_1 _20284_ (.A(_13441_),
    .B(_04777_),
    .X(_13442_));
 sky130_fd_sc_hd__inv_2 _20285_ (.A(\count_1[2] ),
    .Y(_13527_));
 sky130_fd_sc_hd__inv_2 _20286_ (.A(\count_2[2] ),
    .Y(_13535_));
 sky130_fd_sc_hd__xnor2_1 _20287_ (.A(_06010_),
    .B(\hash.CA1.S0.X[15] ),
    .Y(_08136_));
 sky130_fd_sc_hd__xnor2_4 _20288_ (.A(_08136_),
    .B(_06179_),
    .Y(_13552_));
 sky130_fd_sc_hd__xnor2_1 _20289_ (.A(_06016_),
    .B(_06108_),
    .Y(_08137_));
 sky130_fd_sc_hd__xnor2_2 _20290_ (.A(\hash.CA1.S0.X[25] ),
    .B(_08137_),
    .Y(_13556_));
 sky130_fd_sc_hd__xnor2_1 _20291_ (.A(\hash.CA1.S0.X[6] ),
    .B(\hash.CA1.S0.X[17] ),
    .Y(_08138_));
 sky130_fd_sc_hd__xnor2_1 _20292_ (.A(net1094),
    .B(_08138_),
    .Y(_13560_));
 sky130_fd_sc_hd__xnor2_1 _20293_ (.A(\hash.CA1.S0.X[7] ),
    .B(\hash.CA1.S0.X[18] ),
    .Y(_08139_));
 sky130_fd_sc_hd__xnor2_1 _20294_ (.A(_06211_),
    .B(_08139_),
    .Y(_13564_));
 sky130_fd_sc_hd__xnor2_1 _20295_ (.A(_06043_),
    .B(_06133_),
    .Y(_08140_));
 sky130_fd_sc_hd__xnor2_2 _20296_ (.A(_06218_),
    .B(_08140_),
    .Y(_13568_));
 sky130_fd_sc_hd__xor2_1 _20297_ (.A(\hash.CA1.S0.X[9] ),
    .B(_06148_),
    .X(_08141_));
 sky130_fd_sc_hd__xnor2_1 _20298_ (.A(_06226_),
    .B(_08141_),
    .Y(_13572_));
 sky130_fd_sc_hd__xnor2_1 _20299_ (.A(\hash.CA1.S0.X[10] ),
    .B(_06156_),
    .Y(_08142_));
 sky130_fd_sc_hd__xnor2_4 _20300_ (.A(_06234_),
    .B(_08142_),
    .Y(_13576_));
 sky130_fd_sc_hd__xnor2_1 _20301_ (.A(_06066_),
    .B(\hash.CA1.S0.X[22] ),
    .Y(_08143_));
 sky130_fd_sc_hd__xnor2_2 _20302_ (.A(_06269_),
    .B(_08143_),
    .Y(_13580_));
 sky130_fd_sc_hd__xnor2_1 _20303_ (.A(_13235_),
    .B(_06073_),
    .Y(_08144_));
 sky130_fd_sc_hd__nor2_1 _20304_ (.A(net349),
    .B(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__xor2_1 _20305_ (.A(_06172_),
    .B(_08145_),
    .X(_13584_));
 sky130_fd_sc_hd__xor2_1 _20306_ (.A(_13241_),
    .B(_06079_),
    .X(_08146_));
 sky130_fd_sc_hd__xnor2_1 _20307_ (.A(_07935_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__nor2_1 _20308_ (.A(net349),
    .B(_08147_),
    .Y(_13588_));
 sky130_fd_sc_hd__xnor2_1 _20309_ (.A(_05998_),
    .B(_06091_),
    .Y(_08148_));
 sky130_fd_sc_hd__xnor2_1 _20310_ (.A(_06212_),
    .B(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand2_1 _20311_ (.A(_06002_),
    .B(_08149_),
    .Y(_13592_));
 sky130_fd_sc_hd__xnor2_1 _20312_ (.A(\hash.CA1.S0.X[3] ),
    .B(\hash.CA1.S0.X[15] ),
    .Y(_08150_));
 sky130_fd_sc_hd__xnor2_1 _20313_ (.A(net1094),
    .B(_08150_),
    .Y(_13596_));
 sky130_fd_sc_hd__xnor2_1 _20314_ (.A(_06010_),
    .B(\hash.CA1.S0.X[16] ),
    .Y(_08151_));
 sky130_fd_sc_hd__xnor2_1 _20315_ (.A(_06211_),
    .B(_08151_),
    .Y(_13600_));
 sky130_fd_sc_hd__xnor2_1 _20316_ (.A(_06016_),
    .B(\hash.CA1.S0.X[17] ),
    .Y(_08152_));
 sky130_fd_sc_hd__xnor2_1 _20317_ (.A(_06218_),
    .B(_08152_),
    .Y(_13604_));
 sky130_fd_sc_hd__xnor2_1 _20318_ (.A(_06024_),
    .B(\hash.CA1.S0.X[18] ),
    .Y(_08153_));
 sky130_fd_sc_hd__xnor2_1 _20319_ (.A(_06226_),
    .B(_08153_),
    .Y(_13608_));
 sky130_fd_sc_hd__xnor2_1 _20320_ (.A(_06032_),
    .B(_06133_),
    .Y(_08154_));
 sky130_fd_sc_hd__xnor2_1 _20321_ (.A(_06234_),
    .B(_08154_),
    .Y(_13612_));
 sky130_fd_sc_hd__xor2_1 _20322_ (.A(_06043_),
    .B(_06148_),
    .X(_08155_));
 sky130_fd_sc_hd__xnor2_4 _20323_ (.A(_06269_),
    .B(_08155_),
    .Y(_13616_));
 sky130_fd_sc_hd__xnor2_1 _20324_ (.A(_13235_),
    .B(_06155_),
    .Y(_08156_));
 sky130_fd_sc_hd__nand2_1 _20325_ (.A(_06002_),
    .B(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__xor2_1 _20326_ (.A(\hash.CA1.S0.X[9] ),
    .B(_08157_),
    .X(_13620_));
 sky130_fd_sc_hd__xnor2_1 _20327_ (.A(_13241_),
    .B(_06164_),
    .Y(_08158_));
 sky130_fd_sc_hd__nor2_2 _20328_ (.A(net349),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__xnor2_1 _20329_ (.A(\hash.CA1.S0.X[10] ),
    .B(_08159_),
    .Y(_13624_));
 sky130_fd_sc_hd__nor2_1 _20330_ (.A(_12109_),
    .B(_06172_),
    .Y(_08160_));
 sky130_fd_sc_hd__a21oi_2 _20331_ (.A1(_05999_),
    .A2(_06172_),
    .B1(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__xnor2_2 _20332_ (.A(_06066_),
    .B(_08161_),
    .Y(_13628_));
 sky130_fd_sc_hd__xnor2_1 _20333_ (.A(\hash.CA1.S0.X[3] ),
    .B(\hash.CA1.S0.X[12] ),
    .Y(_08162_));
 sky130_fd_sc_hd__xnor2_1 _20334_ (.A(_06179_),
    .B(_08162_),
    .Y(_13632_));
 sky130_fd_sc_hd__xor2_1 _20335_ (.A(_06010_),
    .B(_06080_),
    .X(_08163_));
 sky130_fd_sc_hd__xnor2_1 _20336_ (.A(\hash.CA1.S0.X[25] ),
    .B(_08163_),
    .Y(_13636_));
 sky130_fd_sc_hd__xnor2_2 _20337_ (.A(\hash.CA1.S0.X[5] ),
    .B(\hash.CA1.S0.X[14] ),
    .Y(_08164_));
 sky130_fd_sc_hd__xnor2_1 _20338_ (.A(net1094),
    .B(_08164_),
    .Y(_13640_));
 sky130_fd_sc_hd__xnor2_1 _20339_ (.A(\hash.CA1.S0.X[6] ),
    .B(\hash.CA1.S0.X[15] ),
    .Y(_08165_));
 sky130_fd_sc_hd__xnor2_1 _20340_ (.A(_06211_),
    .B(_08165_),
    .Y(_13644_));
 sky130_fd_sc_hd__xnor2_1 _20341_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06108_),
    .Y(_08166_));
 sky130_fd_sc_hd__xnor2_1 _20342_ (.A(_06218_),
    .B(_08166_),
    .Y(_13648_));
 sky130_fd_sc_hd__xor2_1 _20343_ (.A(_06043_),
    .B(\hash.CA1.S0.X[17] ),
    .X(_08167_));
 sky130_fd_sc_hd__xnor2_1 _20344_ (.A(_06226_),
    .B(_08167_),
    .Y(_13652_));
 sky130_fd_sc_hd__xnor2_1 _20345_ (.A(\hash.CA1.S0.X[9] ),
    .B(\hash.CA1.S0.X[18] ),
    .Y(_08168_));
 sky130_fd_sc_hd__xnor2_1 _20346_ (.A(_06234_),
    .B(_08168_),
    .Y(_13656_));
 sky130_fd_sc_hd__xnor2_1 _20347_ (.A(\hash.CA1.S0.X[10] ),
    .B(_06133_),
    .Y(_08169_));
 sky130_fd_sc_hd__xnor2_1 _20348_ (.A(_06269_),
    .B(_08169_),
    .Y(_13660_));
 sky130_fd_sc_hd__mux2i_2 _20349_ (.A0(_13235_),
    .A1(_00658_),
    .S(_06066_),
    .Y(_08170_));
 sky130_fd_sc_hd__xor2_1 _20350_ (.A(_06148_),
    .B(_08170_),
    .X(_13664_));
 sky130_fd_sc_hd__inv_1 _20351_ (.A(_12370_),
    .Y(_13668_));
 sky130_fd_sc_hd__inv_1 _20352_ (.A(_12385_),
    .Y(_13676_));
 sky130_fd_sc_hd__inv_1 _20353_ (.A(_12393_),
    .Y(_13688_));
 sky130_fd_sc_hd__clkinv_2 _20354_ (.A(_12401_),
    .Y(_13700_));
 sky130_fd_sc_hd__inv_1 _20355_ (.A(_06800_),
    .Y(_13703_));
 sky130_fd_sc_hd__inv_1 _20356_ (.A(_12406_),
    .Y(_13707_));
 sky130_fd_sc_hd__inv_1 _20357_ (.A(_12417_),
    .Y(_13724_));
 sky130_fd_sc_hd__nor2b_1 _20358_ (.A(net350),
    .B_N(\hash.CA2.a_dash[11] ),
    .Y(_13727_));
 sky130_fd_sc_hd__clkinv_1 _20359_ (.A(_12422_),
    .Y(_13731_));
 sky130_fd_sc_hd__inv_1 _20360_ (.A(_12430_),
    .Y(_13743_));
 sky130_fd_sc_hd__inv_1 _20361_ (.A(_12435_),
    .Y(_13750_));
 sky130_fd_sc_hd__inv_1 _20362_ (.A(_12440_),
    .Y(_13757_));
 sky130_fd_sc_hd__inv_1 _20363_ (.A(_12445_),
    .Y(_13764_));
 sky130_fd_sc_hd__inv_1 _20364_ (.A(_12465_),
    .Y(_13796_));
 sky130_fd_sc_hd__inv_1 _20365_ (.A(_12470_),
    .Y(_13803_));
 sky130_fd_sc_hd__nor2b_1 _20366_ (.A(net351),
    .B_N(\hash.CA2.a_dash[24] ),
    .Y(_13806_));
 sky130_fd_sc_hd__inv_1 _20367_ (.A(_12475_),
    .Y(_13810_));
 sky130_fd_sc_hd__nor2_1 _20368_ (.A(net351),
    .B(_04734_),
    .Y(_13813_));
 sky130_fd_sc_hd__clkinv_1 _20369_ (.A(_12480_),
    .Y(_13817_));
 sky130_fd_sc_hd__inv_1 _20370_ (.A(_12485_),
    .Y(_13824_));
 sky130_fd_sc_hd__inv_1 _20371_ (.A(_12490_),
    .Y(_13831_));
 sky130_fd_sc_hd__mux2i_1 _20372_ (.A0(\hash.CA2.e_dash[2] ),
    .A1(\hash.CA2.S1.X[2] ),
    .S(_06513_),
    .Y(_08171_));
 sky130_fd_sc_hd__nand2_1 _20373_ (.A(_06002_),
    .B(_08171_),
    .Y(_13870_));
 sky130_fd_sc_hd__inv_1 _20374_ (.A(_12517_),
    .Y(_13881_));
 sky130_fd_sc_hd__mux2_4 _20375_ (.A0(\hash.CA1.f[4] ),
    .A1(\hash.CA2.e_dash[4] ),
    .S(_06524_),
    .X(_13887_));
 sky130_fd_sc_hd__inv_1 _20376_ (.A(_12522_),
    .Y(_13891_));
 sky130_fd_sc_hd__nand2_1 _20377_ (.A(\hash.CA2.e_dash[5] ),
    .B(_06531_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_1 _20378_ (.A(\hash.CA1.f[5] ),
    .B(\hash.CA1.S1.X[5] ),
    .Y(_08173_));
 sky130_fd_sc_hd__nand2_1 _20379_ (.A(_08172_),
    .B(_08173_),
    .Y(_13897_));
 sky130_fd_sc_hd__mux2i_2 _20380_ (.A0(_12399_),
    .A1(_06428_),
    .S(\hash.CA1.S1.X[7] ),
    .Y(_13914_));
 sky130_fd_sc_hd__nor3_1 _20381_ (.A(net354),
    .B(\hash.CA2.e_dash[8] ),
    .C(_06551_),
    .Y(_08174_));
 sky130_fd_sc_hd__a21oi_4 _20382_ (.A1(_06433_),
    .A2(_06552_),
    .B1(_08174_),
    .Y(_13922_));
 sky130_fd_sc_hd__inv_1 _20383_ (.A(_12542_),
    .Y(_13925_));
 sky130_fd_sc_hd__nand2_1 _20384_ (.A(\hash.CA2.e_dash[9] ),
    .B(_06559_),
    .Y(_08175_));
 sky130_fd_sc_hd__nand2_1 _20385_ (.A(_06438_),
    .B(\hash.CA1.S1.X[9] ),
    .Y(_08176_));
 sky130_fd_sc_hd__nand2_2 _20386_ (.A(_08175_),
    .B(_08176_),
    .Y(_13931_));
 sky130_fd_sc_hd__nand2_2 _20387_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA1.S1.X[10] ),
    .Y(_08177_));
 sky130_fd_sc_hd__nand2_2 _20388_ (.A(_12410_),
    .B(_06568_),
    .Y(_08178_));
 sky130_fd_sc_hd__nand2_2 _20389_ (.A(_08177_),
    .B(_08178_),
    .Y(_13940_));
 sky130_fd_sc_hd__inv_1 _20390_ (.A(_12552_),
    .Y(_13943_));
 sky130_fd_sc_hd__inv_2 _20391_ (.A(_12557_),
    .Y(_13953_));
 sky130_fd_sc_hd__nand2_1 _20392_ (.A(\hash.CA2.e_dash[12] ),
    .B(_06581_),
    .Y(_08179_));
 sky130_fd_sc_hd__nand2_1 _20393_ (.A(\hash.CA1.f[12] ),
    .B(\hash.CA1.S1.X[12] ),
    .Y(_08180_));
 sky130_fd_sc_hd__nand2_1 _20394_ (.A(_08179_),
    .B(_08180_),
    .Y(_13959_));
 sky130_fd_sc_hd__nand2_1 _20395_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_08181_));
 sky130_fd_sc_hd__nand2_1 _20396_ (.A(_12423_),
    .B(_06589_),
    .Y(_08182_));
 sky130_fd_sc_hd__nand2_2 _20397_ (.A(_08181_),
    .B(_08182_),
    .Y(_13968_));
 sky130_fd_sc_hd__inv_1 _20398_ (.A(_12572_),
    .Y(_13979_));
 sky130_fd_sc_hd__clkinv_1 _20399_ (.A(\hash.CA2.S1.X[15] ),
    .Y(_08183_));
 sky130_fd_sc_hd__nor3_2 _20400_ (.A(net351),
    .B(\hash.CA2.e_dash[15] ),
    .C(_06610_),
    .Y(_08184_));
 sky130_fd_sc_hd__a21oi_4 _20401_ (.A1(_08183_),
    .A2(_06610_),
    .B1(_08184_),
    .Y(_13985_));
 sky130_fd_sc_hd__inv_1 _20402_ (.A(_12577_),
    .Y(_13989_));
 sky130_fd_sc_hd__mux2_4 _20403_ (.A0(\hash.CA1.f[17] ),
    .A1(\hash.CA2.e_dash[17] ),
    .S(_06624_),
    .X(_14004_));
 sky130_fd_sc_hd__mux2_1 _20404_ (.A0(\hash.CA1.f[19] ),
    .A1(\hash.CA2.e_dash[19] ),
    .S(_06642_),
    .X(_14020_));
 sky130_fd_sc_hd__mux2_1 _20405_ (.A0(_12452_),
    .A1(\hash.CA2.S1.X[20] ),
    .S(\hash.CA1.S1.X[20] ),
    .X(_14028_));
 sky130_fd_sc_hd__mux2_1 _20406_ (.A0(_12455_),
    .A1(\hash.CA2.S1.X[21] ),
    .S(\hash.CA1.S1.X[21] ),
    .X(_14036_));
 sky130_fd_sc_hd__inv_1 _20407_ (.A(_12607_),
    .Y(_14039_));
 sky130_fd_sc_hd__mux2_1 _20408_ (.A0(_12458_),
    .A1(\hash.CA2.S1.X[22] ),
    .S(\hash.CA1.S1.X[22] ),
    .X(_14045_));
 sky130_fd_sc_hd__inv_1 _20409_ (.A(_12612_),
    .Y(_14049_));
 sky130_fd_sc_hd__nor2_1 _20410_ (.A(\hash.CA2.S1.X[23] ),
    .B(_06665_),
    .Y(_08185_));
 sky130_fd_sc_hd__a21oi_2 _20411_ (.A1(_12463_),
    .A2(_06665_),
    .B1(_08185_),
    .Y(_14055_));
 sky130_fd_sc_hd__inv_1 _20412_ (.A(_12617_),
    .Y(_14059_));
 sky130_fd_sc_hd__inv_1 _20413_ (.A(_12622_),
    .Y(_14069_));
 sky130_fd_sc_hd__inv_1 _20414_ (.A(_12627_),
    .Y(_14079_));
 sky130_fd_sc_hd__inv_1 _20415_ (.A(\hash.CA2.S1.X[26] ),
    .Y(_08186_));
 sky130_fd_sc_hd__nor3_1 _20416_ (.A(net352),
    .B(\hash.CA2.e_dash[26] ),
    .C(_06689_),
    .Y(_08187_));
 sky130_fd_sc_hd__a21oi_4 _20417_ (.A1(_08186_),
    .A2(_06689_),
    .B1(_08187_),
    .Y(_14085_));
 sky130_fd_sc_hd__inv_1 _20418_ (.A(_12637_),
    .Y(_14097_));
 sky130_fd_sc_hd__inv_1 _20419_ (.A(_12642_),
    .Y(_14107_));
 sky130_fd_sc_hd__mux2_8 _20420_ (.A0(\hash.CA2.S1.X[29] ),
    .A1(_12491_),
    .S(_06712_),
    .X(_14113_));
 sky130_fd_sc_hd__mux2_8 _20421_ (.A0(\hash.CA2.e_dash[30] ),
    .A1(\hash.CA1.f[30] ),
    .S(net1047),
    .X(_14122_));
 sky130_fd_sc_hd__inv_1 _20422_ (.A(_12652_),
    .Y(_14125_));
 sky130_fd_sc_hd__inv_1 _20423_ (.A(_12673_),
    .Y(_14129_));
 sky130_fd_sc_hd__inv_1 _20424_ (.A(_12678_),
    .Y(_14133_));
 sky130_fd_sc_hd__inv_1 _20425_ (.A(_12683_),
    .Y(_14137_));
 sky130_fd_sc_hd__inv_1 _20426_ (.A(_12690_),
    .Y(_14141_));
 sky130_fd_sc_hd__clkinv_1 _20427_ (.A(_12699_),
    .Y(_14145_));
 sky130_fd_sc_hd__clkinv_1 _20428_ (.A(_12707_),
    .Y(_14149_));
 sky130_fd_sc_hd__inv_1 _20429_ (.A(_12712_),
    .Y(_14153_));
 sky130_fd_sc_hd__inv_1 _20430_ (.A(_12717_),
    .Y(_12719_));
 sky130_fd_sc_hd__inv_1 _20431_ (.A(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__inv_1 _20432_ (.A(_12761_),
    .Y(_12763_));
 sky130_fd_sc_hd__clkinv_2 _20433_ (.A(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__clkinv_1 _20434_ (.A(_12812_),
    .Y(_12813_));
 sky130_fd_sc_hd__inv_1 _20435_ (.A(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__inv_1 _20436_ (.A(_12878_),
    .Y(_14199_));
 sky130_fd_sc_hd__xnor2_1 _20437_ (.A(_05998_),
    .B(_06079_),
    .Y(_08188_));
 sky130_fd_sc_hd__xnor2_2 _20438_ (.A(_08188_),
    .B(_06164_),
    .Y(_08189_));
 sky130_fd_sc_hd__nor2_2 _20439_ (.A(_08189_),
    .B(net349),
    .Y(_14203_));
 sky130_fd_sc_hd__inv_1 _20440_ (.A(_12664_),
    .Y(_14206_));
 sky130_fd_sc_hd__inv_1 _20441_ (.A(_12374_),
    .Y(\hash.CA1.p4[0] ));
 sky130_fd_sc_hd__inv_4 _20442_ (.A(_13232_),
    .Y(_12076_));
 sky130_fd_sc_hd__inv_1 _20443_ (.A(_13856_),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_1 _20444_ (.A(_13545_),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_1 _20445_ (.A(\hash.CA1.p4[1] ),
    .Y(_12895_));
 sky130_fd_sc_hd__inv_1 _20446_ (.A(_13850_),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_1 _20447_ (.A(_13853_),
    .Y(_00824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_983 ();
 sky130_fd_sc_hd__nor2_1 _20449_ (.A(net1044),
    .B(\count15_1[1] ),
    .Y(_00907_));
 sky130_fd_sc_hd__nor2b_1 _20450_ (.A(net1043),
    .B_N(_00644_),
    .Y(_00908_));
 sky130_fd_sc_hd__xnor2_1 _20451_ (.A(net524),
    .B(_13521_),
    .Y(_08191_));
 sky130_fd_sc_hd__nor2_1 _20452_ (.A(net1043),
    .B(_08191_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand3_1 _20453_ (.A(net537),
    .B(\count15_1[2] ),
    .C(net524),
    .Y(_08192_));
 sky130_fd_sc_hd__xor2_1 _20454_ (.A(net521),
    .B(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__nor2_1 _20455_ (.A(net1043),
    .B(_08193_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand3_1 _20456_ (.A(net524),
    .B(net521),
    .C(_13521_),
    .Y(_08194_));
 sky130_fd_sc_hd__xor2_1 _20457_ (.A(net558),
    .B(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__nor2_1 _20458_ (.A(net1043),
    .B(_08195_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _20459_ (.A(_09731_),
    .B(net517),
    .Y(_00912_));
 sky130_fd_sc_hd__nor2b_1 _20460_ (.A(net784),
    .B_N(_00648_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_1 _20461_ (.A(net504),
    .B(_13525_),
    .Y(_08196_));
 sky130_fd_sc_hd__nor2_1 _20462_ (.A(net784),
    .B(_08196_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand3_1 _20463_ (.A(net516),
    .B(net511),
    .C(\count15_2[3] ),
    .Y(_08197_));
 sky130_fd_sc_hd__xor2_1 _20464_ (.A(net501),
    .B(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__nor2_1 _20465_ (.A(net1043),
    .B(_08198_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand3_2 _20466_ (.A(\count15_2[3] ),
    .B(net501),
    .C(_13525_),
    .Y(_08199_));
 sky130_fd_sc_hd__xor2_1 _20467_ (.A(\count15_2[5] ),
    .B(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__nor2_1 _20468_ (.A(net1043),
    .B(_08200_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_1 _20469_ (.A(net784),
    .B(net496),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2b_1 _20470_ (.A(net1043),
    .B_N(_00645_),
    .Y(_00918_));
 sky130_fd_sc_hd__xnor2_1 _20471_ (.A(net484),
    .B(_13522_),
    .Y(_08201_));
 sky130_fd_sc_hd__nor2_1 _20472_ (.A(net1043),
    .B(_08201_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand3_1 _20473_ (.A(net556),
    .B(net491),
    .C(\count16_1[3] ),
    .Y(_08202_));
 sky130_fd_sc_hd__xor2_1 _20474_ (.A(\count16_1[4] ),
    .B(_08202_),
    .X(_08203_));
 sky130_fd_sc_hd__nor2_1 _20475_ (.A(net1043),
    .B(_08203_),
    .Y(_00920_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_982 ();
 sky130_fd_sc_hd__nand3_1 _20477_ (.A(net484),
    .B(\count16_1[4] ),
    .C(_13522_),
    .Y(_08205_));
 sky130_fd_sc_hd__xor2_1 _20478_ (.A(\count16_1[5] ),
    .B(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__nor2_1 _20479_ (.A(net1043),
    .B(_08206_),
    .Y(_00921_));
 sky130_fd_sc_hd__nor2_1 _20480_ (.A(net1044),
    .B(net553),
    .Y(_00922_));
 sky130_fd_sc_hd__nor2b_1 _20481_ (.A(net1043),
    .B_N(_00649_),
    .Y(_00923_));
 sky130_fd_sc_hd__xnor2_1 _20482_ (.A(net464),
    .B(_13526_),
    .Y(_08207_));
 sky130_fd_sc_hd__nor2_1 _20483_ (.A(net1043),
    .B(_08207_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand3_1 _20484_ (.A(net477),
    .B(net471),
    .C(net464),
    .Y(_08208_));
 sky130_fd_sc_hd__xor2_1 _20485_ (.A(\count16_2[4] ),
    .B(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__nor2_1 _20486_ (.A(net1044),
    .B(_08209_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand3_1 _20487_ (.A(net464),
    .B(\count16_2[4] ),
    .C(_13526_),
    .Y(_08210_));
 sky130_fd_sc_hd__xor2_1 _20488_ (.A(\count16_2[5] ),
    .B(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__nor2_1 _20489_ (.A(net1043),
    .B(_08211_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_1 _20490_ (.A(_09731_),
    .B(\count2_1[1] ),
    .Y(_00927_));
 sky130_fd_sc_hd__or2_0 _20491_ (.A(net1043),
    .B(_00642_),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_1 _20492_ (.A(\count2_1[3] ),
    .B(_13546_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand2_1 _20493_ (.A(_09731_),
    .B(_08212_),
    .Y(_00929_));
 sky130_fd_sc_hd__nand3_1 _20494_ (.A(net456),
    .B(net551),
    .C(net443),
    .Y(_08213_));
 sky130_fd_sc_hd__xor2_1 _20495_ (.A(\count2_1[4] ),
    .B(_08213_),
    .X(_08214_));
 sky130_fd_sc_hd__nor2_1 _20496_ (.A(net1043),
    .B(_08214_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand3_1 _20497_ (.A(\count2_1[3] ),
    .B(\count2_1[4] ),
    .C(_13546_),
    .Y(_08215_));
 sky130_fd_sc_hd__xor2_1 _20498_ (.A(\count2_1[5] ),
    .B(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__nor2_1 _20499_ (.A(net1043),
    .B(_08216_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _20500_ (.A(_09731_),
    .B(net436),
    .Y(_00932_));
 sky130_fd_sc_hd__or2_0 _20501_ (.A(net1044),
    .B(_00646_),
    .X(_00933_));
 sky130_fd_sc_hd__xnor2_1 _20502_ (.A(\count2_2[3] ),
    .B(_13523_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_1 _20503_ (.A(_09731_),
    .B(_08217_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand3_1 _20504_ (.A(net433),
    .B(net430),
    .C(net423),
    .Y(_08218_));
 sky130_fd_sc_hd__xor2_1 _20505_ (.A(\count2_2[4] ),
    .B(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__nor2_1 _20506_ (.A(net1043),
    .B(_08219_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand3_1 _20507_ (.A(\count2_2[3] ),
    .B(net548),
    .C(_13523_),
    .Y(_08220_));
 sky130_fd_sc_hd__xor2_1 _20508_ (.A(\count2_2[5] ),
    .B(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__nor2_1 _20509_ (.A(net1044),
    .B(_08221_),
    .Y(_00936_));
 sky130_fd_sc_hd__nor2_1 _20510_ (.A(net1044),
    .B(net547),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2b_1 _20511_ (.A(net1043),
    .B_N(_00643_),
    .Y(_00938_));
 sky130_fd_sc_hd__xnor2_1 _20512_ (.A(\count7_1[3] ),
    .B(_13520_),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2_1 _20513_ (.A(_09731_),
    .B(_08222_),
    .Y(_00939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_981 ();
 sky130_fd_sc_hd__nand3_1 _20515_ (.A(net417),
    .B(\count7_1[2] ),
    .C(net546),
    .Y(_08224_));
 sky130_fd_sc_hd__xor2_1 _20516_ (.A(net402),
    .B(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__nor2_1 _20517_ (.A(net1043),
    .B(_08225_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand3_1 _20518_ (.A(net546),
    .B(net402),
    .C(_13520_),
    .Y(_08226_));
 sky130_fd_sc_hd__xor2_1 _20519_ (.A(\count7_1[5] ),
    .B(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__nor2_1 _20520_ (.A(net1043),
    .B(_08227_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_1 _20521_ (.A(_09731_),
    .B(\count7_2[1] ),
    .Y(_00942_));
 sky130_fd_sc_hd__nor2b_1 _20522_ (.A(net1044),
    .B_N(_00647_),
    .Y(_00943_));
 sky130_fd_sc_hd__xnor2_1 _20523_ (.A(\count7_2[3] ),
    .B(_13524_),
    .Y(_08228_));
 sky130_fd_sc_hd__nand2_1 _20524_ (.A(_09731_),
    .B(_08228_),
    .Y(_00944_));
 sky130_fd_sc_hd__nand3_1 _20525_ (.A(net544),
    .B(net393),
    .C(net385),
    .Y(_08229_));
 sky130_fd_sc_hd__xor2_1 _20526_ (.A(net383),
    .B(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__nor2_1 _20527_ (.A(net1043),
    .B(_08230_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand3_1 _20528_ (.A(net386),
    .B(net383),
    .C(_13524_),
    .Y(_08231_));
 sky130_fd_sc_hd__xor2_1 _20529_ (.A(\count7_2[5] ),
    .B(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__nor2_1 _20530_ (.A(net1043),
    .B(_08232_),
    .Y(_00946_));
 sky130_fd_sc_hd__xnor2_1 _20531_ (.A(_00650_),
    .B(_00128_),
    .Y(_08233_));
 sky130_fd_sc_hd__nor2_1 _20532_ (.A(net1044),
    .B(_08233_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _20533_ (.A(\count_1[2] ),
    .B(_00128_),
    .Y(_08234_));
 sky130_fd_sc_hd__nand2_1 _20534_ (.A(_00651_),
    .B(_09727_),
    .Y(_08235_));
 sky130_fd_sc_hd__a21oi_1 _20535_ (.A1(_08234_),
    .A2(_08235_),
    .B1(net1044),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _20536_ (.A(_13533_),
    .B(_09727_),
    .Y(_08236_));
 sky130_fd_sc_hd__xor2_1 _20537_ (.A(\count_1[3] ),
    .B(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__nor2_1 _20538_ (.A(net1044),
    .B(_08237_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand4_1 _20539_ (.A(\count_1[3] ),
    .B(\count_1[2] ),
    .C(\count_1[1] ),
    .D(_09727_),
    .Y(_08238_));
 sky130_fd_sc_hd__xor2_1 _20540_ (.A(\count_1[4] ),
    .B(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__nand2_1 _20541_ (.A(_09731_),
    .B(_08239_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand4_1 _20542_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C(_13533_),
    .D(_09727_),
    .Y(_08240_));
 sky130_fd_sc_hd__xor2_1 _20543_ (.A(\count_1[5] ),
    .B(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__nor2_1 _20544_ (.A(net1044),
    .B(_08241_),
    .Y(_00951_));
 sky130_fd_sc_hd__xnor2_1 _20545_ (.A(_00652_),
    .B(_00128_),
    .Y(_08242_));
 sky130_fd_sc_hd__nor2_1 _20546_ (.A(net1044),
    .B(_08242_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand2_1 _20547_ (.A(\count_2[2] ),
    .B(_00128_),
    .Y(_08243_));
 sky130_fd_sc_hd__nand2_1 _20548_ (.A(_00653_),
    .B(_09727_),
    .Y(_08244_));
 sky130_fd_sc_hd__a21oi_1 _20549_ (.A1(_08243_),
    .A2(_08244_),
    .B1(net1044),
    .Y(_00953_));
 sky130_fd_sc_hd__xnor2_1 _20550_ (.A(\count_2[3] ),
    .B(_13541_),
    .Y(_08245_));
 sky130_fd_sc_hd__a21oi_1 _20551_ (.A1(_09727_),
    .A2(_08245_),
    .B1(net1043),
    .Y(_00954_));
 sky130_fd_sc_hd__nand3_1 _20552_ (.A(\count_2[3] ),
    .B(\count_2[2] ),
    .C(\count_2[1] ),
    .Y(_08246_));
 sky130_fd_sc_hd__xor2_1 _20553_ (.A(\count_2[4] ),
    .B(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__nand3_1 _20554_ (.A(_09731_),
    .B(_09727_),
    .C(_08247_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand3_1 _20555_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_13541_),
    .Y(_08248_));
 sky130_fd_sc_hd__nand2_1 _20556_ (.A(\count_2[6] ),
    .B(\count_2[5] ),
    .Y(_08249_));
 sky130_fd_sc_hd__nor2_1 _20557_ (.A(_08248_),
    .B(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__a211oi_1 _20558_ (.A1(_09802_),
    .A2(_08248_),
    .B1(_08250_),
    .C1(net1043),
    .Y(_00956_));
 sky130_fd_sc_hd__nor2b_1 _20559_ (.A(\count_2[6] ),
    .B_N(_09726_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_1 _20560_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .Y(_08252_));
 sky130_fd_sc_hd__nor2_1 _20561_ (.A(_08246_),
    .B(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__mux2i_1 _20562_ (.A0(\count_2[6] ),
    .A1(_08251_),
    .S(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__nor2_1 _20563_ (.A(net1043),
    .B(_08254_),
    .Y(_00957_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_980 ();
 sky130_fd_sc_hd__nand3_2 _20565_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(\count_hash1[5] ),
    .Y(_08256_));
 sky130_fd_sc_hd__nor2_4 _20566_ (.A(\count_hash1[6] ),
    .B(_08256_),
    .Y(_08257_));
 sky130_fd_sc_hd__nand2_8 _20567_ (.A(_12920_),
    .B(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__xnor2_1 _20568_ (.A(\count_hash1[1] ),
    .B(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__nor2_1 _20569_ (.A(net540),
    .B(_08259_),
    .Y(_00958_));
 sky130_fd_sc_hd__nor2_1 _20570_ (.A(_12910_),
    .B(_08258_),
    .Y(_08260_));
 sky130_fd_sc_hd__a21oi_1 _20571_ (.A1(_00655_),
    .A2(_08258_),
    .B1(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__nor2_1 _20572_ (.A(net540),
    .B(_08261_),
    .Y(_00959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_978 ();
 sky130_fd_sc_hd__nor2_1 _20575_ (.A(_10348_),
    .B(_08257_),
    .Y(_08264_));
 sky130_fd_sc_hd__nor2_1 _20576_ (.A(net540),
    .B(_08264_),
    .Y(_00960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_977 ();
 sky130_fd_sc_hd__a21oi_1 _20578_ (.A1(_10352_),
    .A2(_08258_),
    .B1(net540),
    .Y(_00961_));
 sky130_fd_sc_hd__xor2_4 _20579_ (.A(\count_hash1[5] ),
    .B(_10372_),
    .X(_08266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_974 ();
 sky130_fd_sc_hd__a21oi_1 _20583_ (.A1(_08266_),
    .A2(_08258_),
    .B1(net540),
    .Y(_00962_));
 sky130_fd_sc_hd__or4_1 _20584_ (.A(_12920_),
    .B(_00654_),
    .C(\count_hash1[6] ),
    .D(_09873_),
    .X(_08270_));
 sky130_fd_sc_hd__o21ai_0 _20585_ (.A1(_00654_),
    .A2(_09873_),
    .B1(\count_hash1[6] ),
    .Y(_08271_));
 sky130_fd_sc_hd__a21oi_1 _20586_ (.A1(_08270_),
    .A2(_08271_),
    .B1(net540),
    .Y(_00963_));
 sky130_fd_sc_hd__xnor2_1 _20587_ (.A(\count_hash2[1] ),
    .B(_08258_),
    .Y(_08272_));
 sky130_fd_sc_hd__nor2_1 _20588_ (.A(net540),
    .B(_08272_),
    .Y(_00964_));
 sky130_fd_sc_hd__nor2_1 _20589_ (.A(_12900_),
    .B(_08258_),
    .Y(_08273_));
 sky130_fd_sc_hd__a21oi_1 _20590_ (.A1(_00657_),
    .A2(_08258_),
    .B1(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__nor2_1 _20591_ (.A(net540),
    .B(_08274_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _20592_ (.A(_12908_),
    .B(_08258_),
    .Y(_08275_));
 sky130_fd_sc_hd__xor2_1 _20593_ (.A(\count_hash2[3] ),
    .B(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__nor2_1 _20594_ (.A(net540),
    .B(_08276_),
    .Y(_00966_));
 sky130_fd_sc_hd__a21oi_1 _20595_ (.A1(_12920_),
    .A2(_08257_),
    .B1(_09856_),
    .Y(_08277_));
 sky130_fd_sc_hd__xnor2_1 _20596_ (.A(\count_hash2[4] ),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__nor2_1 _20597_ (.A(net540),
    .B(_08278_),
    .Y(_00967_));
 sky130_fd_sc_hd__a21oi_1 _20598_ (.A1(_12920_),
    .A2(_08257_),
    .B1(_09866_),
    .Y(_08279_));
 sky130_fd_sc_hd__xnor2_1 _20599_ (.A(\count_hash2[5] ),
    .B(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__nor2_1 _20600_ (.A(net540),
    .B(_08280_),
    .Y(_00968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_972 ();
 sky130_fd_sc_hd__xnor2_4 _20603_ (.A(\count_hash1[3] ),
    .B(_12920_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand2_8 _20604_ (.A(net322),
    .B(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_969 ();
 sky130_fd_sc_hd__nor2_1 _20608_ (.A(_12912_),
    .B(net325),
    .Y(_08288_));
 sky130_fd_sc_hd__nor2_1 _20609_ (.A(net332),
    .B(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_965 ();
 sky130_fd_sc_hd__nor2_4 _20614_ (.A(_10352_),
    .B(_08283_),
    .Y(_08294_));
 sky130_fd_sc_hd__nor2_1 _20615_ (.A(_08266_),
    .B(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__o221ai_1 _20616_ (.A1(_12918_),
    .A2(_08284_),
    .B1(_08289_),
    .B2(_12916_),
    .C1(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__xnor2_4 _20617_ (.A(\count_hash1[4] ),
    .B(_10351_),
    .Y(_08297_));
 sky130_fd_sc_hd__nand2_8 _20618_ (.A(_08297_),
    .B(_08266_),
    .Y(_08298_));
 sky130_fd_sc_hd__nor2_4 _20619_ (.A(net331),
    .B(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_964 ();
 sky130_fd_sc_hd__nand2_2 _20621_ (.A(net332),
    .B(_10373_),
    .Y(_08301_));
 sky130_fd_sc_hd__o22ai_2 _20622_ (.A1(_08297_),
    .A2(_08301_),
    .B1(_08298_),
    .B2(net332),
    .Y(_08302_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_963 ();
 sky130_fd_sc_hd__nand2_8 _20624_ (.A(_10352_),
    .B(_10348_),
    .Y(_08304_));
 sky130_fd_sc_hd__nand2_1 _20625_ (.A(_12912_),
    .B(net295),
    .Y(_08305_));
 sky130_fd_sc_hd__nor2_2 _20626_ (.A(_08304_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__a221oi_4 _20627_ (.A1(_12916_),
    .A2(_08299_),
    .B1(_08302_),
    .B2(_12918_),
    .C1(_08306_),
    .Y(_08307_));
 sky130_fd_sc_hd__nand2_2 _20628_ (.A(net323),
    .B(_08266_),
    .Y(_08308_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_962 ();
 sky130_fd_sc_hd__nor2_4 _20630_ (.A(_12911_),
    .B(_12916_),
    .Y(_08310_));
 sky130_fd_sc_hd__nor3_1 _20631_ (.A(net331),
    .B(_08308_),
    .C(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_961 ();
 sky130_fd_sc_hd__nor2_4 _20633_ (.A(net325),
    .B(net296),
    .Y(_08313_));
 sky130_fd_sc_hd__nand2_1 _20634_ (.A(_12916_),
    .B(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__nand2_4 _20635_ (.A(net325),
    .B(net296),
    .Y(_08315_));
 sky130_fd_sc_hd__nand2_1 _20636_ (.A(_12912_),
    .B(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_960 ();
 sky130_fd_sc_hd__a21oi_1 _20638_ (.A1(_08314_),
    .A2(_08316_),
    .B1(_08283_),
    .Y(_08318_));
 sky130_fd_sc_hd__nor2_1 _20639_ (.A(_08311_),
    .B(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__or2_4 _20640_ (.A(\count_hash1[6] ),
    .B(_09874_),
    .X(_08320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_959 ();
 sky130_fd_sc_hd__nor2_4 _20642_ (.A(net540),
    .B(_08320_),
    .Y(_08322_));
 sky130_fd_sc_hd__nor2_4 _20643_ (.A(_12911_),
    .B(_12918_),
    .Y(_08323_));
 sky130_fd_sc_hd__or3_1 _20644_ (.A(_12911_),
    .B(_12912_),
    .C(_12916_),
    .X(_08324_));
 sky130_fd_sc_hd__nor2_4 _20645_ (.A(net332),
    .B(_10373_),
    .Y(_08325_));
 sky130_fd_sc_hd__nand2_1 _20646_ (.A(_08324_),
    .B(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__o21ai_2 _20647_ (.A1(_08283_),
    .A2(_08323_),
    .B1(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__nand2_4 _20648_ (.A(_10352_),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__nor2_2 _20649_ (.A(_12911_),
    .B(_12912_),
    .Y(_08329_));
 sky130_fd_sc_hd__nor2_4 _20650_ (.A(_12916_),
    .B(_12918_),
    .Y(_08330_));
 sky130_fd_sc_hd__nand2_4 _20651_ (.A(_08329_),
    .B(_08330_),
    .Y(_08331_));
 sky130_fd_sc_hd__nor2_4 _20652_ (.A(_08297_),
    .B(_10373_),
    .Y(_08332_));
 sky130_fd_sc_hd__nor2_4 _20653_ (.A(_12912_),
    .B(_12916_),
    .Y(_08333_));
 sky130_fd_sc_hd__a21oi_2 _20654_ (.A1(net333),
    .A2(_08333_),
    .B1(_08325_),
    .Y(_08334_));
 sky130_fd_sc_hd__o22ai_4 _20655_ (.A1(_08331_),
    .A2(_08332_),
    .B1(_08334_),
    .B2(_08297_),
    .Y(_08335_));
 sky130_fd_sc_hd__nand2_8 _20656_ (.A(_08328_),
    .B(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__nand2_8 _20657_ (.A(_08322_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_958 ();
 sky130_fd_sc_hd__a31oi_1 _20659_ (.A1(_08296_),
    .A2(_08307_),
    .A3(_08319_),
    .B1(_08337_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_2 _20660_ (.A(_08297_),
    .B(net332),
    .Y(_08339_));
 sky130_fd_sc_hd__nand2_4 _20661_ (.A(_12911_),
    .B(_08266_),
    .Y(_08340_));
 sky130_fd_sc_hd__o21ai_2 _20662_ (.A1(_08339_),
    .A2(_08340_),
    .B1(_08336_),
    .Y(_08341_));
 sky130_fd_sc_hd__a21oi_1 _20663_ (.A1(_12916_),
    .A2(_10373_),
    .B1(_08339_),
    .Y(_08342_));
 sky130_fd_sc_hd__nor2_4 _20664_ (.A(_08297_),
    .B(_08266_),
    .Y(_08343_));
 sky130_fd_sc_hd__a21oi_1 _20665_ (.A1(net332),
    .A2(_08343_),
    .B1(_08310_),
    .Y(_08344_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_957 ();
 sky130_fd_sc_hd__a21oi_1 _20667_ (.A1(_12916_),
    .A2(_08297_),
    .B1(_12911_),
    .Y(_08346_));
 sky130_fd_sc_hd__o21ai_0 _20668_ (.A1(_08332_),
    .A2(_08346_),
    .B1(_08283_),
    .Y(_08347_));
 sky130_fd_sc_hd__o21ai_0 _20669_ (.A1(_12912_),
    .A2(_08344_),
    .B1(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nor2_1 _20670_ (.A(_08342_),
    .B(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__nor2_4 _20671_ (.A(\count_hash1[6] ),
    .B(_09874_),
    .Y(_08350_));
 sky130_fd_sc_hd__o21ai_0 _20672_ (.A1(_08341_),
    .A2(_08349_),
    .B1(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__nand2b_1 _20673_ (.A_N(net540),
    .B(_08351_),
    .Y(_00970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_956 ();
 sky130_fd_sc_hd__and2_4 _20675_ (.A(_12918_),
    .B(net333),
    .X(_08353_));
 sky130_fd_sc_hd__a21oi_1 _20676_ (.A1(_12912_),
    .A2(_08283_),
    .B1(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__nor2_4 _20677_ (.A(_08297_),
    .B(net332),
    .Y(_08355_));
 sky130_fd_sc_hd__nor2_4 _20678_ (.A(_08283_),
    .B(_08266_),
    .Y(_08356_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_955 ();
 sky130_fd_sc_hd__o21ai_0 _20680_ (.A1(_08355_),
    .A2(_08356_),
    .B1(_12911_),
    .Y(_08358_));
 sky130_fd_sc_hd__nor2_4 _20681_ (.A(net323),
    .B(net331),
    .Y(_08359_));
 sky130_fd_sc_hd__nor2_4 _20682_ (.A(_08297_),
    .B(_08283_),
    .Y(_08360_));
 sky130_fd_sc_hd__nor2_4 _20683_ (.A(_08359_),
    .B(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__nand2_4 _20684_ (.A(_08297_),
    .B(net294),
    .Y(_08362_));
 sky130_fd_sc_hd__a21oi_1 _20685_ (.A1(_08283_),
    .A2(_08362_),
    .B1(_12916_),
    .Y(_08363_));
 sky130_fd_sc_hd__a21oi_1 _20686_ (.A1(_08324_),
    .A2(_08284_),
    .B1(_12918_),
    .Y(_08364_));
 sky130_fd_sc_hd__a211o_1 _20687_ (.A1(_08266_),
    .A2(_08361_),
    .B1(_08363_),
    .C1(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__nor2_4 _20688_ (.A(_08283_),
    .B(net295),
    .Y(_08366_));
 sky130_fd_sc_hd__nor2_4 _20689_ (.A(net331),
    .B(_08266_),
    .Y(_08367_));
 sky130_fd_sc_hd__a22oi_1 _20690_ (.A1(_12916_),
    .A2(_08366_),
    .B1(_08367_),
    .B2(_12912_),
    .Y(_08368_));
 sky130_fd_sc_hd__nor2_2 _20691_ (.A(net325),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__and2_4 _20692_ (.A(_08328_),
    .B(_08335_),
    .X(_08370_));
 sky130_fd_sc_hd__a211oi_2 _20693_ (.A1(_08332_),
    .A2(_08353_),
    .B1(_08369_),
    .C1(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__o2111ai_1 _20694_ (.A1(_08315_),
    .A2(_08354_),
    .B1(_08358_),
    .C1(_08365_),
    .D1(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_954 ();
 sky130_fd_sc_hd__a21o_1 _20696_ (.A1(_08350_),
    .A2(_08372_),
    .B1(net540),
    .X(_00971_));
 sky130_fd_sc_hd__nor2_4 _20697_ (.A(_08366_),
    .B(_08367_),
    .Y(_08374_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_953 ();
 sky130_fd_sc_hd__o22ai_1 _20699_ (.A1(_08283_),
    .A2(_08362_),
    .B1(_08374_),
    .B2(_08297_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand2_4 _20700_ (.A(net331),
    .B(_08266_),
    .Y(_08377_));
 sky130_fd_sc_hd__nand2_4 _20701_ (.A(_12918_),
    .B(_08297_),
    .Y(_08378_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_952 ();
 sky130_fd_sc_hd__o22ai_1 _20703_ (.A1(net295),
    .A2(_08284_),
    .B1(_08362_),
    .B2(_08283_),
    .Y(_08380_));
 sky130_fd_sc_hd__nand2_1 _20704_ (.A(_12911_),
    .B(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__o21ai_0 _20705_ (.A1(_08377_),
    .A2(_08378_),
    .B1(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__a21oi_1 _20706_ (.A1(_12916_),
    .A2(_08376_),
    .B1(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__a21oi_1 _20707_ (.A1(_12911_),
    .A2(_08359_),
    .B1(_08306_),
    .Y(_08384_));
 sky130_fd_sc_hd__a21oi_1 _20708_ (.A1(_08383_),
    .A2(_08384_),
    .B1(_08337_),
    .Y(_00972_));
 sky130_fd_sc_hd__o21ai_0 _20709_ (.A1(_08299_),
    .A2(_08360_),
    .B1(_12918_),
    .Y(_08385_));
 sky130_fd_sc_hd__o21ai_0 _20710_ (.A1(_08356_),
    .A2(_08313_),
    .B1(_12912_),
    .Y(_08386_));
 sky130_fd_sc_hd__nor2_1 _20711_ (.A(net325),
    .B(_08266_),
    .Y(_08387_));
 sky130_fd_sc_hd__o21ai_0 _20712_ (.A1(_08355_),
    .A2(_08387_),
    .B1(_12911_),
    .Y(_08388_));
 sky130_fd_sc_hd__nor2_1 _20713_ (.A(_08266_),
    .B(_08359_),
    .Y(_08389_));
 sky130_fd_sc_hd__o21ai_0 _20714_ (.A1(_08299_),
    .A2(_08389_),
    .B1(_12916_),
    .Y(_08390_));
 sky130_fd_sc_hd__nand4_1 _20715_ (.A(_08385_),
    .B(_08386_),
    .C(_08388_),
    .D(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__o21ai_0 _20716_ (.A1(_08341_),
    .A2(_08391_),
    .B1(_08350_),
    .Y(_08392_));
 sky130_fd_sc_hd__nand2b_1 _20717_ (.A_N(net540),
    .B(_08392_),
    .Y(_00973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_951 ();
 sky130_fd_sc_hd__nand2_2 _20719_ (.A(_08283_),
    .B(net295),
    .Y(_08394_));
 sky130_fd_sc_hd__o21ai_0 _20720_ (.A1(_08283_),
    .A2(_08298_),
    .B1(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__a22o_1 _20721_ (.A1(_12918_),
    .A2(_08356_),
    .B1(_08374_),
    .B2(_12916_),
    .X(_08396_));
 sky130_fd_sc_hd__nand2_1 _20722_ (.A(_12911_),
    .B(_10373_),
    .Y(_08397_));
 sky130_fd_sc_hd__a21oi_1 _20723_ (.A1(_08378_),
    .A2(_08397_),
    .B1(net332),
    .Y(_08398_));
 sky130_fd_sc_hd__a221oi_1 _20724_ (.A1(_12912_),
    .A2(_08395_),
    .B1(_08396_),
    .B2(net325),
    .C1(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__a21oi_2 _20725_ (.A1(_08383_),
    .A2(_08399_),
    .B1(_08337_),
    .Y(_00974_));
 sky130_fd_sc_hd__nor2_1 _20726_ (.A(_08283_),
    .B(_08330_),
    .Y(_08400_));
 sky130_fd_sc_hd__o221ai_1 _20727_ (.A1(_12916_),
    .A2(_08304_),
    .B1(_08400_),
    .B2(_12912_),
    .C1(_08389_),
    .Y(_08401_));
 sky130_fd_sc_hd__nand2_1 _20728_ (.A(_12918_),
    .B(_10373_),
    .Y(_08402_));
 sky130_fd_sc_hd__nand2_2 _20729_ (.A(_08340_),
    .B(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__o21ai_4 _20730_ (.A1(_12912_),
    .A2(_08403_),
    .B1(_08359_),
    .Y(_08404_));
 sky130_fd_sc_hd__a31oi_1 _20731_ (.A1(_08328_),
    .A2(_08401_),
    .A3(_08404_),
    .B1(_08337_),
    .Y(_00975_));
 sky130_fd_sc_hd__and2_4 _20732_ (.A(_12918_),
    .B(net295),
    .X(_08405_));
 sky130_fd_sc_hd__a21oi_1 _20733_ (.A1(_12912_),
    .A2(_08266_),
    .B1(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__o21ai_0 _20734_ (.A1(_08297_),
    .A2(_08406_),
    .B1(_08314_),
    .Y(_08407_));
 sky130_fd_sc_hd__nand2_1 _20735_ (.A(_08283_),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__nor2_1 _20736_ (.A(_12912_),
    .B(_12918_),
    .Y(_08409_));
 sky130_fd_sc_hd__a21oi_1 _20737_ (.A1(_08297_),
    .A2(_08409_),
    .B1(_08283_),
    .Y(_08410_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_950 ();
 sky130_fd_sc_hd__nor2_1 _20739_ (.A(_12918_),
    .B(net331),
    .Y(_08412_));
 sky130_fd_sc_hd__a21oi_1 _20740_ (.A1(net332),
    .A2(_08313_),
    .B1(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__o21ai_1 _20741_ (.A1(_08283_),
    .A2(_08323_),
    .B1(_10352_),
    .Y(_08414_));
 sky130_fd_sc_hd__o221ai_1 _20742_ (.A1(_08266_),
    .A2(_08410_),
    .B1(_08413_),
    .B2(_12911_),
    .C1(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__a21oi_1 _20743_ (.A1(_08408_),
    .A2(_08415_),
    .B1(_08337_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_1 _20744_ (.A(net325),
    .B(_08377_),
    .Y(_08416_));
 sky130_fd_sc_hd__o21ai_0 _20745_ (.A1(_08283_),
    .A2(_08298_),
    .B1(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__nand2_1 _20746_ (.A(_08315_),
    .B(_08298_),
    .Y(_08418_));
 sky130_fd_sc_hd__nor3_1 _20747_ (.A(_08266_),
    .B(_08330_),
    .C(_08284_),
    .Y(_08419_));
 sky130_fd_sc_hd__a31oi_2 _20748_ (.A1(_12911_),
    .A2(net332),
    .A3(_08418_),
    .B1(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__o21ai_0 _20749_ (.A1(_08332_),
    .A2(_08356_),
    .B1(_12916_),
    .Y(_08421_));
 sky130_fd_sc_hd__o21ai_0 _20750_ (.A1(net332),
    .A2(_08313_),
    .B1(_12918_),
    .Y(_08422_));
 sky130_fd_sc_hd__nand4_1 _20751_ (.A(_08336_),
    .B(_08420_),
    .C(_08421_),
    .D(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__a21oi_1 _20752_ (.A1(_12912_),
    .A2(_08417_),
    .B1(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__o21bai_1 _20753_ (.A1(_08320_),
    .A2(_08424_),
    .B1_N(net540),
    .Y(_00977_));
 sky130_fd_sc_hd__nor2_1 _20754_ (.A(_08343_),
    .B(_08313_),
    .Y(_08425_));
 sky130_fd_sc_hd__nand2_1 _20755_ (.A(_08323_),
    .B(_08343_),
    .Y(_08426_));
 sky130_fd_sc_hd__o21ai_0 _20756_ (.A1(_12912_),
    .A2(_10373_),
    .B1(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__or2_4 _20757_ (.A(_12912_),
    .B(_12918_),
    .X(_08428_));
 sky130_fd_sc_hd__o22ai_1 _20758_ (.A1(net325),
    .A2(_08367_),
    .B1(_08428_),
    .B2(_08355_),
    .Y(_08429_));
 sky130_fd_sc_hd__a21oi_1 _20759_ (.A1(_08283_),
    .A2(_08427_),
    .B1(_08429_),
    .Y(_08430_));
 sky130_fd_sc_hd__a221oi_1 _20760_ (.A1(_12918_),
    .A2(_08294_),
    .B1(_08425_),
    .B2(_12916_),
    .C1(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__nor2_1 _20761_ (.A(_08337_),
    .B(_08431_),
    .Y(_00978_));
 sky130_fd_sc_hd__a21oi_1 _20762_ (.A1(_12912_),
    .A2(_08297_),
    .B1(_12916_),
    .Y(_08432_));
 sky130_fd_sc_hd__nor2_1 _20763_ (.A(net333),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__a211oi_1 _20764_ (.A1(_12911_),
    .A2(_08339_),
    .B1(_08433_),
    .C1(_08266_),
    .Y(_08434_));
 sky130_fd_sc_hd__a221oi_1 _20765_ (.A1(_12918_),
    .A2(_08294_),
    .B1(_08361_),
    .B2(_12912_),
    .C1(_10373_),
    .Y(_08435_));
 sky130_fd_sc_hd__nor2_1 _20766_ (.A(_10373_),
    .B(_08333_),
    .Y(_08436_));
 sky130_fd_sc_hd__a21oi_1 _20767_ (.A1(_08328_),
    .A2(_08333_),
    .B1(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand2_1 _20768_ (.A(_08266_),
    .B(_08328_),
    .Y(_08438_));
 sky130_fd_sc_hd__o21ai_0 _20769_ (.A1(_08283_),
    .A2(_08437_),
    .B1(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__o21ai_0 _20770_ (.A1(_08283_),
    .A2(_08362_),
    .B1(_08331_),
    .Y(_08440_));
 sky130_fd_sc_hd__a21oi_2 _20771_ (.A1(net325),
    .A2(_08439_),
    .B1(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__o211ai_1 _20772_ (.A1(_08434_),
    .A2(_08435_),
    .B1(_08307_),
    .C1(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a21o_4 _20773_ (.A1(_08350_),
    .A2(_08442_),
    .B1(net540),
    .X(_00979_));
 sky130_fd_sc_hd__o21ai_0 _20774_ (.A1(net295),
    .A2(_08304_),
    .B1(_08394_),
    .Y(_08443_));
 sky130_fd_sc_hd__nand2_2 _20775_ (.A(_12912_),
    .B(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__nand2_1 _20776_ (.A(_08359_),
    .B(_08405_),
    .Y(_08445_));
 sky130_fd_sc_hd__a21oi_1 _20777_ (.A1(net332),
    .A2(_08428_),
    .B1(_12916_),
    .Y(_08446_));
 sky130_fd_sc_hd__nor2_2 _20778_ (.A(_08362_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__a31oi_4 _20779_ (.A1(_12911_),
    .A2(net325),
    .A3(_08366_),
    .B1(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__nor2_2 _20780_ (.A(_12911_),
    .B(net331),
    .Y(_08449_));
 sky130_fd_sc_hd__nor2_1 _20781_ (.A(_12918_),
    .B(_08283_),
    .Y(_08450_));
 sky130_fd_sc_hd__nor2_1 _20782_ (.A(_08449_),
    .B(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__o211ai_1 _20783_ (.A1(_12916_),
    .A2(_08451_),
    .B1(_08304_),
    .C1(_08266_),
    .Y(_08452_));
 sky130_fd_sc_hd__a41oi_2 _20784_ (.A1(_08444_),
    .A2(_08445_),
    .A3(_08448_),
    .A4(_08452_),
    .B1(_08337_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _20785_ (.A(_12918_),
    .B(_08266_),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_1 _20786_ (.A(_12912_),
    .B(_08374_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand2_2 _20787_ (.A(_12916_),
    .B(_08356_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand3_1 _20788_ (.A(_08453_),
    .B(_08454_),
    .C(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__nand2_2 _20789_ (.A(_08297_),
    .B(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__a21oi_1 _20790_ (.A1(_08340_),
    .A2(_08402_),
    .B1(_08283_),
    .Y(_08458_));
 sky130_fd_sc_hd__o21ai_1 _20791_ (.A1(_08436_),
    .A2(_08458_),
    .B1(net325),
    .Y(_08459_));
 sky130_fd_sc_hd__a31oi_1 _20792_ (.A1(_08296_),
    .A2(_08457_),
    .A3(_08459_),
    .B1(_08337_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_1 _20793_ (.A(_08305_),
    .B(_08453_),
    .Y(_08460_));
 sky130_fd_sc_hd__o21ai_0 _20794_ (.A1(_12916_),
    .A2(_08460_),
    .B1(_08294_),
    .Y(_08461_));
 sky130_fd_sc_hd__o31ai_1 _20795_ (.A1(net295),
    .A2(_08304_),
    .A3(_08310_),
    .B1(_08445_),
    .Y(_08462_));
 sky130_fd_sc_hd__a221oi_1 _20796_ (.A1(_12912_),
    .A2(_08299_),
    .B1(_08451_),
    .B2(_08343_),
    .C1(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__a31oi_1 _20797_ (.A1(_08408_),
    .A2(_08461_),
    .A3(_08463_),
    .B1(_08337_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _20798_ (.A(_12916_),
    .B(_08297_),
    .Y(_08464_));
 sky130_fd_sc_hd__nor2_2 _20799_ (.A(_12912_),
    .B(_08283_),
    .Y(_08465_));
 sky130_fd_sc_hd__a221oi_1 _20800_ (.A1(_08283_),
    .A2(_08310_),
    .B1(_08464_),
    .B2(_08465_),
    .C1(net295),
    .Y(_08466_));
 sky130_fd_sc_hd__a21oi_1 _20801_ (.A1(_12911_),
    .A2(_08284_),
    .B1(_12912_),
    .Y(_08467_));
 sky130_fd_sc_hd__nor2_1 _20802_ (.A(_12911_),
    .B(_08361_),
    .Y(_08468_));
 sky130_fd_sc_hd__nor3_1 _20803_ (.A(_08266_),
    .B(_08467_),
    .C(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__nor2_1 _20804_ (.A(_08466_),
    .B(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__nor2_1 _20805_ (.A(_08337_),
    .B(_08470_),
    .Y(_00983_));
 sky130_fd_sc_hd__a22oi_1 _20806_ (.A1(_12918_),
    .A2(_08360_),
    .B1(_08428_),
    .B2(_08359_),
    .Y(_08471_));
 sky130_fd_sc_hd__nand2_1 _20807_ (.A(net333),
    .B(_08333_),
    .Y(_08472_));
 sky130_fd_sc_hd__o211ai_1 _20808_ (.A1(net333),
    .A2(_08331_),
    .B1(_08472_),
    .C1(_08313_),
    .Y(_08473_));
 sky130_fd_sc_hd__inv_1 _20809_ (.A(_08455_),
    .Y(_08474_));
 sky130_fd_sc_hd__nand2_1 _20810_ (.A(_10373_),
    .B(_08428_),
    .Y(_08475_));
 sky130_fd_sc_hd__a21oi_1 _20811_ (.A1(_08340_),
    .A2(_08475_),
    .B1(net332),
    .Y(_08476_));
 sky130_fd_sc_hd__o21ai_0 _20812_ (.A1(_08474_),
    .A2(_08476_),
    .B1(net324),
    .Y(_08477_));
 sky130_fd_sc_hd__o2111ai_1 _20813_ (.A1(_08266_),
    .A2(_08471_),
    .B1(_08473_),
    .C1(_08477_),
    .D1(_08441_),
    .Y(_08478_));
 sky130_fd_sc_hd__a21o_4 _20814_ (.A1(_08350_),
    .A2(_08478_),
    .B1(net540),
    .X(_00984_));
 sky130_fd_sc_hd__o21ai_0 _20815_ (.A1(_12911_),
    .A2(_08405_),
    .B1(_08283_),
    .Y(_08479_));
 sky130_fd_sc_hd__o21ai_0 _20816_ (.A1(_08283_),
    .A2(_08343_),
    .B1(_12916_),
    .Y(_08480_));
 sky130_fd_sc_hd__a31oi_1 _20817_ (.A1(_08444_),
    .A2(_08479_),
    .A3(_08480_),
    .B1(_08337_),
    .Y(_00985_));
 sky130_fd_sc_hd__nor2_1 _20818_ (.A(_08266_),
    .B(_08323_),
    .Y(_08481_));
 sky130_fd_sc_hd__a21oi_1 _20819_ (.A1(_12916_),
    .A2(_08266_),
    .B1(_08481_),
    .Y(_08482_));
 sky130_fd_sc_hd__a22oi_1 _20820_ (.A1(_12911_),
    .A2(_08297_),
    .B1(_08343_),
    .B2(_12918_),
    .Y(_08483_));
 sky130_fd_sc_hd__o21ai_0 _20821_ (.A1(_08332_),
    .A2(_08294_),
    .B1(_12912_),
    .Y(_08484_));
 sky130_fd_sc_hd__o221ai_2 _20822_ (.A1(_08304_),
    .A2(_08482_),
    .B1(_08483_),
    .B2(_10348_),
    .C1(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__nor3_1 _20823_ (.A(_08370_),
    .B(_08369_),
    .C(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__o21bai_1 _20824_ (.A1(_08320_),
    .A2(_08486_),
    .B1_N(net540),
    .Y(_00986_));
 sky130_fd_sc_hd__o21ai_0 _20825_ (.A1(_08297_),
    .A2(_08330_),
    .B1(_08283_),
    .Y(_08487_));
 sky130_fd_sc_hd__nand2_1 _20826_ (.A(_08378_),
    .B(_08465_),
    .Y(_08488_));
 sky130_fd_sc_hd__o21ai_1 _20827_ (.A1(net330),
    .A2(_08308_),
    .B1(_08362_),
    .Y(_08489_));
 sky130_fd_sc_hd__a32oi_2 _20828_ (.A1(net295),
    .A2(_08487_),
    .A3(_08488_),
    .B1(_08489_),
    .B2(_12911_),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_2 _20829_ (.A(_08377_),
    .B(_08394_),
    .Y(_08491_));
 sky130_fd_sc_hd__nand3_1 _20830_ (.A(_12911_),
    .B(net325),
    .C(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__a31oi_2 _20831_ (.A1(_08473_),
    .A2(_08490_),
    .A3(_08492_),
    .B1(_08337_),
    .Y(_00987_));
 sky130_fd_sc_hd__a22oi_1 _20832_ (.A1(_12918_),
    .A2(_08332_),
    .B1(_08425_),
    .B2(_12912_),
    .Y(_08493_));
 sky130_fd_sc_hd__nor2_1 _20833_ (.A(_08283_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__nand2_1 _20834_ (.A(_12911_),
    .B(_08343_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand2_1 _20835_ (.A(_12916_),
    .B(_08315_),
    .Y(_08496_));
 sky130_fd_sc_hd__a21oi_1 _20836_ (.A1(_08495_),
    .A2(_08496_),
    .B1(net333),
    .Y(_08497_));
 sky130_fd_sc_hd__a211oi_1 _20837_ (.A1(_08313_),
    .A2(_08353_),
    .B1(_08494_),
    .C1(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__a21oi_1 _20838_ (.A1(_08404_),
    .A2(_08498_),
    .B1(_08337_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _20839_ (.A(_12911_),
    .B(_08361_),
    .Y(_08499_));
 sky130_fd_sc_hd__o21ai_0 _20840_ (.A1(_08333_),
    .A2(_08284_),
    .B1(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2_1 _20841_ (.A(_08266_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__a21oi_1 _20842_ (.A1(_12918_),
    .A2(_08315_),
    .B1(_12916_),
    .Y(_08502_));
 sky130_fd_sc_hd__nor2_1 _20843_ (.A(_08325_),
    .B(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__a21oi_1 _20844_ (.A1(_08313_),
    .A2(_08450_),
    .B1(_08355_),
    .Y(_08504_));
 sky130_fd_sc_hd__o21ai_0 _20845_ (.A1(_12912_),
    .A2(_08503_),
    .B1(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__a21oi_1 _20846_ (.A1(_08501_),
    .A2(_08505_),
    .B1(_08337_),
    .Y(_00989_));
 sky130_fd_sc_hd__nor2_1 _20847_ (.A(_12918_),
    .B(_08297_),
    .Y(_08506_));
 sky130_fd_sc_hd__a21oi_1 _20848_ (.A1(_08297_),
    .A2(_08449_),
    .B1(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__o21ai_0 _20849_ (.A1(net322),
    .A2(_08409_),
    .B1(net331),
    .Y(_08508_));
 sky130_fd_sc_hd__o211ai_1 _20850_ (.A1(_12916_),
    .A2(_08507_),
    .B1(_08508_),
    .C1(net295),
    .Y(_08509_));
 sky130_fd_sc_hd__a21oi_1 _20851_ (.A1(_12916_),
    .A2(net322),
    .B1(_12911_),
    .Y(_08510_));
 sky130_fd_sc_hd__or3_1 _20852_ (.A(net295),
    .B(_08359_),
    .C(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__a31oi_2 _20853_ (.A1(_08307_),
    .A2(_08509_),
    .A3(_08511_),
    .B1(_08337_),
    .Y(_00990_));
 sky130_fd_sc_hd__a222oi_1 _20854_ (.A1(_12912_),
    .A2(_08301_),
    .B1(_08366_),
    .B2(_12916_),
    .C1(_08491_),
    .C2(_12911_),
    .Y(_08512_));
 sky130_fd_sc_hd__nor2_1 _20855_ (.A(_08297_),
    .B(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__a21oi_1 _20856_ (.A1(_12916_),
    .A2(_08299_),
    .B1(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__a31oi_1 _20857_ (.A1(_08404_),
    .A2(_08490_),
    .A3(_08514_),
    .B1(_08337_),
    .Y(_00991_));
 sky130_fd_sc_hd__o21ai_0 _20858_ (.A1(net332),
    .A2(_10373_),
    .B1(_12916_),
    .Y(_08515_));
 sky130_fd_sc_hd__a21oi_1 _20859_ (.A1(_08397_),
    .A2(_08515_),
    .B1(_08297_),
    .Y(_08516_));
 sky130_fd_sc_hd__a21oi_1 _20860_ (.A1(_12912_),
    .A2(_08302_),
    .B1(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__o211ai_1 _20861_ (.A1(_08378_),
    .A2(_08491_),
    .B1(_08517_),
    .C1(_08371_),
    .Y(_08518_));
 sky130_fd_sc_hd__a21o_4 _20862_ (.A1(_08350_),
    .A2(_08518_),
    .B1(net540),
    .X(_00992_));
 sky130_fd_sc_hd__nor2_1 _20863_ (.A(_12911_),
    .B(_08266_),
    .Y(_08519_));
 sky130_fd_sc_hd__nor2_1 _20864_ (.A(net323),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__o22a_1 _20865_ (.A1(_12918_),
    .A2(_08298_),
    .B1(_08520_),
    .B2(_12912_),
    .X(_08521_));
 sky130_fd_sc_hd__o211ai_1 _20866_ (.A1(_12916_),
    .A2(_08521_),
    .B1(_08308_),
    .C1(net330),
    .Y(_08522_));
 sky130_fd_sc_hd__o22ai_1 _20867_ (.A1(_12911_),
    .A2(net331),
    .B1(_08377_),
    .B2(_12918_),
    .Y(_08523_));
 sky130_fd_sc_hd__a21oi_1 _20868_ (.A1(net323),
    .A2(_08523_),
    .B1(_08367_),
    .Y(_08524_));
 sky130_fd_sc_hd__o21ai_0 _20869_ (.A1(_12918_),
    .A2(_08266_),
    .B1(net323),
    .Y(_08525_));
 sky130_fd_sc_hd__nor2_1 _20870_ (.A(_12911_),
    .B(_08283_),
    .Y(_08526_));
 sky130_fd_sc_hd__nand2_1 _20871_ (.A(_08525_),
    .B(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__o21ai_0 _20872_ (.A1(net295),
    .A2(_08412_),
    .B1(_08297_),
    .Y(_08528_));
 sky130_fd_sc_hd__o211ai_1 _20873_ (.A1(_12912_),
    .A2(_08524_),
    .B1(_08527_),
    .C1(_08528_),
    .Y(_08529_));
 sky130_fd_sc_hd__a21oi_1 _20874_ (.A1(_08522_),
    .A2(_08529_),
    .B1(_08337_),
    .Y(_00993_));
 sky130_fd_sc_hd__nand2_1 _20875_ (.A(_12916_),
    .B(_08266_),
    .Y(_08530_));
 sky130_fd_sc_hd__and2_0 _20876_ (.A(_12912_),
    .B(_10373_),
    .X(_08531_));
 sky130_fd_sc_hd__o21ai_0 _20877_ (.A1(_12911_),
    .A2(_08531_),
    .B1(_10352_),
    .Y(_08532_));
 sky130_fd_sc_hd__a21oi_1 _20878_ (.A1(_08530_),
    .A2(_08532_),
    .B1(net333),
    .Y(_08533_));
 sky130_fd_sc_hd__nor2_1 _20879_ (.A(_10373_),
    .B(_08323_),
    .Y(_08534_));
 sky130_fd_sc_hd__a21oi_1 _20880_ (.A1(_12916_),
    .A2(_10373_),
    .B1(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__nand2_1 _20881_ (.A(_12912_),
    .B(_08299_),
    .Y(_08536_));
 sky130_fd_sc_hd__o21ai_0 _20882_ (.A1(_08304_),
    .A2(_08535_),
    .B1(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__nor2_1 _20883_ (.A(net333),
    .B(_08329_),
    .Y(_08538_));
 sky130_fd_sc_hd__o21ai_1 _20884_ (.A1(_08400_),
    .A2(_08538_),
    .B1(_08387_),
    .Y(_08539_));
 sky130_fd_sc_hd__nor4b_1 _20885_ (.A(_08341_),
    .B(_08533_),
    .C(_08537_),
    .D_N(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__o21bai_1 _20886_ (.A1(_08320_),
    .A2(_08540_),
    .B1_N(net540),
    .Y(_00994_));
 sky130_fd_sc_hd__nand2_1 _20887_ (.A(_08294_),
    .B(_08436_),
    .Y(_08541_));
 sky130_fd_sc_hd__nand2_2 _20888_ (.A(_08336_),
    .B(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__nor2_1 _20889_ (.A(_08360_),
    .B(_08432_),
    .Y(_08543_));
 sky130_fd_sc_hd__nor2_1 _20890_ (.A(_12911_),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__nor3_1 _20891_ (.A(_12916_),
    .B(_10352_),
    .C(net333),
    .Y(_08545_));
 sky130_fd_sc_hd__nor3_1 _20892_ (.A(_08266_),
    .B(_08544_),
    .C(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__o22ai_1 _20893_ (.A1(_08378_),
    .A2(_08374_),
    .B1(_08530_),
    .B2(_08297_),
    .Y(_08547_));
 sky130_fd_sc_hd__nor4_1 _20894_ (.A(_08537_),
    .B(_08542_),
    .C(_08546_),
    .D(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__o21bai_1 _20895_ (.A1(_08320_),
    .A2(_08548_),
    .B1_N(net540),
    .Y(_00995_));
 sky130_fd_sc_hd__o21ai_0 _20896_ (.A1(_08283_),
    .A2(_08475_),
    .B1(_08515_),
    .Y(_08549_));
 sky130_fd_sc_hd__a22oi_1 _20897_ (.A1(_08360_),
    .A2(_08481_),
    .B1(_08549_),
    .B2(_08297_),
    .Y(_08550_));
 sky130_fd_sc_hd__a21oi_1 _20898_ (.A1(_08514_),
    .A2(_08550_),
    .B1(_08337_),
    .Y(_00996_));
 sky130_fd_sc_hd__o21ai_0 _20899_ (.A1(_08531_),
    .A2(_08534_),
    .B1(_08294_),
    .Y(_08551_));
 sky130_fd_sc_hd__nor2_1 _20900_ (.A(_12916_),
    .B(_08377_),
    .Y(_08552_));
 sky130_fd_sc_hd__a21oi_1 _20901_ (.A1(_12916_),
    .A2(_08301_),
    .B1(_12911_),
    .Y(_08553_));
 sky130_fd_sc_hd__or3_1 _20902_ (.A(_08297_),
    .B(_08552_),
    .C(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__a41oi_1 _20903_ (.A1(_08473_),
    .A2(_08539_),
    .A3(_08551_),
    .A4(_08554_),
    .B1(_08337_),
    .Y(_00997_));
 sky130_fd_sc_hd__a21oi_1 _20904_ (.A1(_12916_),
    .A2(net331),
    .B1(net322),
    .Y(_08555_));
 sky130_fd_sc_hd__a21oi_1 _20905_ (.A1(net331),
    .A2(_08506_),
    .B1(_08449_),
    .Y(_08556_));
 sky130_fd_sc_hd__nor2_1 _20906_ (.A(_12912_),
    .B(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__a21oi_1 _20907_ (.A1(_12912_),
    .A2(_08284_),
    .B1(_12911_),
    .Y(_08558_));
 sky130_fd_sc_hd__nor2_1 _20908_ (.A(_08465_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__o221ai_1 _20909_ (.A1(net322),
    .A2(_08325_),
    .B1(_08559_),
    .B2(_12918_),
    .C1(_08308_),
    .Y(_08560_));
 sky130_fd_sc_hd__o311ai_2 _20910_ (.A1(net295),
    .A2(_08555_),
    .A3(_08557_),
    .B1(_08448_),
    .C1(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__o21ai_0 _20911_ (.A1(_08341_),
    .A2(_08561_),
    .B1(_08350_),
    .Y(_08562_));
 sky130_fd_sc_hd__nand2b_1 _20912_ (.A_N(net540),
    .B(_08562_),
    .Y(_00998_));
 sky130_fd_sc_hd__a21oi_1 _20913_ (.A1(_12916_),
    .A2(_08343_),
    .B1(_12911_),
    .Y(_08563_));
 sky130_fd_sc_hd__a22oi_1 _20914_ (.A1(_12912_),
    .A2(_08343_),
    .B1(_08418_),
    .B2(_12911_),
    .Y(_08564_));
 sky130_fd_sc_hd__o21ai_0 _20915_ (.A1(net332),
    .A2(_08563_),
    .B1(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__nor4b_1 _20916_ (.A(_08462_),
    .B(_08542_),
    .C(_08565_),
    .D_N(_08457_),
    .Y(_08566_));
 sky130_fd_sc_hd__o21bai_1 _20917_ (.A1(_08320_),
    .A2(_08566_),
    .B1_N(net540),
    .Y(_00999_));
 sky130_fd_sc_hd__a22oi_1 _20918_ (.A1(_08353_),
    .A2(_08387_),
    .B1(_08425_),
    .B2(_08538_),
    .Y(_08567_));
 sky130_fd_sc_hd__nand2_2 _20919_ (.A(_12916_),
    .B(_08380_),
    .Y(_08568_));
 sky130_fd_sc_hd__nand3_1 _20920_ (.A(_08420_),
    .B(_08567_),
    .C(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__nor3_1 _20921_ (.A(_08494_),
    .B(_08542_),
    .C(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__o21bai_1 _20922_ (.A1(_08320_),
    .A2(_08570_),
    .B1_N(net540),
    .Y(_01000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_948 ();
 sky130_fd_sc_hd__nor2_4 _20925_ (.A(_12902_),
    .B(_12906_),
    .Y(_08573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_946 ();
 sky130_fd_sc_hd__nor2_4 _20928_ (.A(_12901_),
    .B(_12904_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand2_8 _20929_ (.A(_08573_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand2_8 _20930_ (.A(_08322_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_944 ();
 sky130_fd_sc_hd__or2_4 _20933_ (.A(_12902_),
    .B(_12906_),
    .X(_08581_));
 sky130_fd_sc_hd__nor3_4 _20934_ (.A(_12901_),
    .B(_12904_),
    .C(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_940 ();
 sky130_fd_sc_hd__o21ai_0 _20939_ (.A1(_12901_),
    .A2(_12906_),
    .B1(net339),
    .Y(_08587_));
 sky130_fd_sc_hd__o31ai_1 _20940_ (.A1(net339),
    .A2(net298),
    .A3(_08582_),
    .B1(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__nor2_4 _20941_ (.A(_12901_),
    .B(_12902_),
    .Y(_08589_));
 sky130_fd_sc_hd__nor2_2 _20942_ (.A(net346),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__xnor2_4 _20943_ (.A(\count_hash2[3] ),
    .B(_12908_),
    .Y(_08591_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_939 ();
 sky130_fd_sc_hd__nor2_4 _20945_ (.A(_12904_),
    .B(_12906_),
    .Y(_08593_));
 sky130_fd_sc_hd__nor2_1 _20946_ (.A(net539),
    .B(_08593_),
    .Y(_08594_));
 sky130_fd_sc_hd__o21ai_4 _20947_ (.A1(_08590_),
    .A2(_08594_),
    .B1(net300),
    .Y(_08595_));
 sky130_fd_sc_hd__nand2_4 _20948_ (.A(net339),
    .B(net539),
    .Y(_08596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_937 ();
 sky130_fd_sc_hd__xor2_4 _20951_ (.A(\count_hash2[5] ),
    .B(_09866_),
    .X(_08599_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_935 ();
 sky130_fd_sc_hd__inv_6 _20954_ (.A(_12902_),
    .Y(_08602_));
 sky130_fd_sc_hd__nand2_1 _20955_ (.A(_08602_),
    .B(_08576_),
    .Y(_08603_));
 sky130_fd_sc_hd__a21oi_1 _20956_ (.A1(_12906_),
    .A2(_08599_),
    .B1(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__o22ai_1 _20957_ (.A1(net339),
    .A2(_08595_),
    .B1(_08596_),
    .B2(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__a21oi_2 _20958_ (.A1(net345),
    .A2(_08588_),
    .B1(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__o21bai_4 _20959_ (.A1(_08578_),
    .A2(_08606_),
    .B1_N(net357),
    .Y(_01001_));
 sky130_fd_sc_hd__xnor2_4 _20960_ (.A(\count_hash2[4] ),
    .B(_09856_),
    .Y(_08607_));
 sky130_fd_sc_hd__nand2_8 _20961_ (.A(_08607_),
    .B(net300),
    .Y(_08608_));
 sky130_fd_sc_hd__nor2_4 _20962_ (.A(net347),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_934 ();
 sky130_fd_sc_hd__nand2_4 _20964_ (.A(net347),
    .B(_08599_),
    .Y(_08611_));
 sky130_fd_sc_hd__nor2_2 _20965_ (.A(_08607_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__o21ai_0 _20966_ (.A1(_08609_),
    .A2(_08612_),
    .B1(_12901_),
    .Y(_08613_));
 sky130_fd_sc_hd__nand2_2 _20967_ (.A(_08591_),
    .B(_08599_),
    .Y(_08614_));
 sky130_fd_sc_hd__o21ai_0 _20968_ (.A1(_08573_),
    .A2(_08614_),
    .B1(_08595_),
    .Y(_08615_));
 sky130_fd_sc_hd__a21oi_1 _20969_ (.A1(net339),
    .A2(_08615_),
    .B1(_08582_),
    .Y(_08616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_933 ();
 sky130_fd_sc_hd__nor2_4 _20971_ (.A(net539),
    .B(_08599_),
    .Y(_08618_));
 sky130_fd_sc_hd__nor2_2 _20972_ (.A(_12906_),
    .B(_08614_),
    .Y(_08619_));
 sky130_fd_sc_hd__nor2_1 _20973_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_932 ();
 sky130_fd_sc_hd__nor2_1 _20975_ (.A(_12901_),
    .B(_08611_),
    .Y(_08622_));
 sky130_fd_sc_hd__a31oi_1 _20976_ (.A1(_08602_),
    .A2(_08591_),
    .A3(net298),
    .B1(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_931 ();
 sky130_fd_sc_hd__o221ai_1 _20978_ (.A1(_12904_),
    .A2(_08620_),
    .B1(_08623_),
    .B2(_12906_),
    .C1(_08607_),
    .Y(_08625_));
 sky130_fd_sc_hd__a31oi_1 _20979_ (.A1(_08613_),
    .A2(_08616_),
    .A3(_08625_),
    .B1(_08320_),
    .Y(_08626_));
 sky130_fd_sc_hd__or2_4 _20980_ (.A(net540),
    .B(_08626_),
    .X(_01002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_929 ();
 sky130_fd_sc_hd__nand2_1 _20983_ (.A(net539),
    .B(_08593_),
    .Y(_08629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_928 ();
 sky130_fd_sc_hd__nor2_4 _20985_ (.A(_12902_),
    .B(_12904_),
    .Y(_08631_));
 sky130_fd_sc_hd__nand2_1 _20986_ (.A(net347),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__nor2_4 _20987_ (.A(net339),
    .B(_08599_),
    .Y(_08633_));
 sky130_fd_sc_hd__o211ai_1 _20988_ (.A1(_12901_),
    .A2(_08629_),
    .B1(_08632_),
    .C1(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_927 ();
 sky130_fd_sc_hd__nand2_1 _20990_ (.A(_12902_),
    .B(_08607_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_1 _20991_ (.A(_12906_),
    .B(_09857_),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_1 _20992_ (.A(_08636_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__nor2_4 _20993_ (.A(net539),
    .B(net300),
    .Y(_08639_));
 sky130_fd_sc_hd__o21ai_1 _20994_ (.A1(_12901_),
    .A2(_08638_),
    .B1(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_924 ();
 sky130_fd_sc_hd__a21oi_1 _20998_ (.A1(_12904_),
    .A2(net300),
    .B1(_12901_),
    .Y(_08644_));
 sky130_fd_sc_hd__o21ai_0 _20999_ (.A1(_08607_),
    .A2(_08644_),
    .B1(_08602_),
    .Y(_08645_));
 sky130_fd_sc_hd__nand2_1 _21000_ (.A(net539),
    .B(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__nand2_8 _21001_ (.A(_08607_),
    .B(net539),
    .Y(_08647_));
 sky130_fd_sc_hd__nand2_2 _21002_ (.A(_09857_),
    .B(net346),
    .Y(_08648_));
 sky130_fd_sc_hd__nor2_2 _21003_ (.A(net346),
    .B(_08593_),
    .Y(_08649_));
 sky130_fd_sc_hd__a32oi_1 _21004_ (.A1(_12901_),
    .A2(_08647_),
    .A3(_08648_),
    .B1(_08649_),
    .B2(_09857_),
    .Y(_08650_));
 sky130_fd_sc_hd__nand2_2 _21005_ (.A(_09857_),
    .B(net300),
    .Y(_08651_));
 sky130_fd_sc_hd__nor2_4 _21006_ (.A(_09857_),
    .B(net300),
    .Y(_08652_));
 sky130_fd_sc_hd__nand2_1 _21007_ (.A(net539),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__o21ai_0 _21008_ (.A1(net539),
    .A2(_08651_),
    .B1(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__nand2_2 _21009_ (.A(net347),
    .B(net300),
    .Y(_08655_));
 sky130_fd_sc_hd__nand2_4 _21010_ (.A(_12904_),
    .B(_09857_),
    .Y(_08656_));
 sky130_fd_sc_hd__o22ai_1 _21011_ (.A1(_08655_),
    .A2(_08656_),
    .B1(_08653_),
    .B2(_08573_),
    .Y(_08657_));
 sky130_fd_sc_hd__a21oi_2 _21012_ (.A1(_12901_),
    .A2(_08654_),
    .B1(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand2_4 _21013_ (.A(_12906_),
    .B(net345),
    .Y(_08659_));
 sky130_fd_sc_hd__nor3_2 _21014_ (.A(_12901_),
    .B(_12904_),
    .C(_12906_),
    .Y(_08660_));
 sky130_fd_sc_hd__a21oi_1 _21015_ (.A1(net300),
    .A2(_08659_),
    .B1(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__nor3_1 _21016_ (.A(_12902_),
    .B(_08607_),
    .C(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__nor2_4 _21017_ (.A(net347),
    .B(net300),
    .Y(_08663_));
 sky130_fd_sc_hd__a221oi_1 _21018_ (.A1(_12904_),
    .A2(_08663_),
    .B1(_08618_),
    .B2(_12906_),
    .C1(_09857_),
    .Y(_08664_));
 sky130_fd_sc_hd__nor2_1 _21019_ (.A(_08662_),
    .B(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__a21oi_1 _21020_ (.A1(_08577_),
    .A2(_08639_),
    .B1(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__o211ai_1 _21021_ (.A1(_08599_),
    .A2(_08650_),
    .B1(_08658_),
    .C1(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__a41oi_2 _21022_ (.A1(_08634_),
    .A2(_08640_),
    .A3(_08646_),
    .A4(_08667_),
    .B1(net292),
    .Y(_01003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_923 ();
 sky130_fd_sc_hd__a22oi_1 _21024_ (.A1(net539),
    .A2(_08576_),
    .B1(_08618_),
    .B2(_08607_),
    .Y(_08669_));
 sky130_fd_sc_hd__nand2_4 _21025_ (.A(net339),
    .B(_08599_),
    .Y(_08670_));
 sky130_fd_sc_hd__o21ai_0 _21026_ (.A1(net345),
    .A2(_08633_),
    .B1(_12901_),
    .Y(_08671_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_922 ();
 sky130_fd_sc_hd__nor2_4 _21028_ (.A(net339),
    .B(net539),
    .Y(_08673_));
 sky130_fd_sc_hd__o21ai_0 _21029_ (.A1(_12904_),
    .A2(net298),
    .B1(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand3_1 _21030_ (.A(_08670_),
    .B(_08671_),
    .C(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__o21ai_0 _21031_ (.A1(_12902_),
    .A2(_08669_),
    .B1(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__nor2_1 _21032_ (.A(_08578_),
    .B(_08676_),
    .Y(_01004_));
 sky130_fd_sc_hd__a21oi_2 _21033_ (.A1(_08633_),
    .A2(_08649_),
    .B1(_08582_),
    .Y(_08677_));
 sky130_fd_sc_hd__nand2_1 _21034_ (.A(_08589_),
    .B(_08656_),
    .Y(_08678_));
 sky130_fd_sc_hd__nand2_2 _21035_ (.A(_08639_),
    .B(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__o21ai_0 _21036_ (.A1(_08602_),
    .A2(_08673_),
    .B1(_08637_),
    .Y(_08680_));
 sky130_fd_sc_hd__or3_4 _21037_ (.A(_12902_),
    .B(_12904_),
    .C(_12906_),
    .X(_08681_));
 sky130_fd_sc_hd__a22o_1 _21038_ (.A1(_12901_),
    .A2(net539),
    .B1(_08618_),
    .B2(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__a22oi_1 _21039_ (.A1(net298),
    .A2(_08680_),
    .B1(_08682_),
    .B2(_08607_),
    .Y(_08683_));
 sky130_fd_sc_hd__a31oi_2 _21040_ (.A1(_08677_),
    .A2(_08679_),
    .A3(_08683_),
    .B1(net292),
    .Y(_01005_));
 sky130_fd_sc_hd__nand3_2 _21041_ (.A(net298),
    .B(_08673_),
    .C(_08681_),
    .Y(_08684_));
 sky130_fd_sc_hd__nand2_4 _21042_ (.A(_08647_),
    .B(_08648_),
    .Y(_08685_));
 sky130_fd_sc_hd__nor2_2 _21043_ (.A(_12901_),
    .B(_08591_),
    .Y(_08686_));
 sky130_fd_sc_hd__a21oi_1 _21044_ (.A1(_12901_),
    .A2(_08647_),
    .B1(_12902_),
    .Y(_08687_));
 sky130_fd_sc_hd__a221oi_1 _21045_ (.A1(_08591_),
    .A2(_08652_),
    .B1(_08686_),
    .B2(_08670_),
    .C1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__o22ai_1 _21046_ (.A1(_08599_),
    .A2(_08685_),
    .B1(_08688_),
    .B2(_12906_),
    .Y(_08689_));
 sky130_fd_sc_hd__a21oi_1 _21047_ (.A1(_08684_),
    .A2(_08689_),
    .B1(_08578_),
    .Y(_08690_));
 sky130_fd_sc_hd__or2_0 _21048_ (.A(net357),
    .B(_08690_),
    .X(_01006_));
 sky130_fd_sc_hd__nand2_1 _21049_ (.A(net539),
    .B(_08603_),
    .Y(_08691_));
 sky130_fd_sc_hd__nand2_8 _21050_ (.A(_08607_),
    .B(_08599_),
    .Y(_08692_));
 sky130_fd_sc_hd__a21oi_1 _21051_ (.A1(_08659_),
    .A2(_08691_),
    .B1(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__nand2_2 _21052_ (.A(_12904_),
    .B(_08599_),
    .Y(_08694_));
 sky130_fd_sc_hd__nand2_1 _21053_ (.A(_12902_),
    .B(_09857_),
    .Y(_08695_));
 sky130_fd_sc_hd__nor2_4 _21054_ (.A(_08607_),
    .B(_08599_),
    .Y(_08696_));
 sky130_fd_sc_hd__nor2_2 _21055_ (.A(_08652_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__a221oi_1 _21056_ (.A1(_12904_),
    .A2(_08633_),
    .B1(_08697_),
    .B2(_12901_),
    .C1(net347),
    .Y(_08698_));
 sky130_fd_sc_hd__a31oi_1 _21057_ (.A1(net345),
    .A2(_08694_),
    .A3(_08695_),
    .B1(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__nor2_1 _21058_ (.A(_08693_),
    .B(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__nor2_1 _21059_ (.A(_08578_),
    .B(_08700_),
    .Y(_01007_));
 sky130_fd_sc_hd__nor2_2 _21060_ (.A(_08607_),
    .B(net539),
    .Y(_08701_));
 sky130_fd_sc_hd__a22o_1 _21061_ (.A1(_12906_),
    .A2(_08701_),
    .B1(_08685_),
    .B2(_12902_),
    .X(_08702_));
 sky130_fd_sc_hd__nand2_1 _21062_ (.A(_08599_),
    .B(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__o22ai_1 _21063_ (.A1(_08591_),
    .A2(_08608_),
    .B1(_08614_),
    .B2(_08607_),
    .Y(_08704_));
 sky130_fd_sc_hd__nor2_2 _21064_ (.A(_08602_),
    .B(net539),
    .Y(_08705_));
 sky130_fd_sc_hd__nor3_1 _21065_ (.A(net298),
    .B(_08576_),
    .C(_08596_),
    .Y(_08706_));
 sky130_fd_sc_hd__a221oi_2 _21066_ (.A1(_12906_),
    .A2(_08704_),
    .B1(_08705_),
    .B2(_08633_),
    .C1(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__a21oi_1 _21067_ (.A1(_12901_),
    .A2(_08607_),
    .B1(net539),
    .Y(_08708_));
 sky130_fd_sc_hd__nand2_1 _21068_ (.A(_08656_),
    .B(_08708_),
    .Y(_08709_));
 sky130_fd_sc_hd__a21oi_1 _21069_ (.A1(_08608_),
    .A2(_08681_),
    .B1(_12901_),
    .Y(_08710_));
 sky130_fd_sc_hd__a21oi_1 _21070_ (.A1(_12904_),
    .A2(net298),
    .B1(_08607_),
    .Y(_08711_));
 sky130_fd_sc_hd__nor3_1 _21071_ (.A(net539),
    .B(_08710_),
    .C(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__a31oi_1 _21072_ (.A1(_12906_),
    .A2(net298),
    .A3(_08709_),
    .B1(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__a31oi_1 _21073_ (.A1(_08703_),
    .A2(_08707_),
    .A3(_08713_),
    .B1(_08578_),
    .Y(_08714_));
 sky130_fd_sc_hd__or2_0 _21074_ (.A(net357),
    .B(_08714_),
    .X(_01008_));
 sky130_fd_sc_hd__a21oi_1 _21075_ (.A1(_12906_),
    .A2(_08608_),
    .B1(_12902_),
    .Y(_08715_));
 sky130_fd_sc_hd__nand2_2 _21076_ (.A(_12904_),
    .B(net347),
    .Y(_08716_));
 sky130_fd_sc_hd__mux2i_1 _21077_ (.A0(_12901_),
    .A1(_12906_),
    .S(_08591_),
    .Y(_08717_));
 sky130_fd_sc_hd__o22ai_1 _21078_ (.A1(_08670_),
    .A2(_08716_),
    .B1(_08717_),
    .B2(_08608_),
    .Y(_08718_));
 sky130_fd_sc_hd__nor2_1 _21079_ (.A(_08582_),
    .B(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__a21oi_1 _21080_ (.A1(_08602_),
    .A2(net339),
    .B1(_08591_),
    .Y(_08720_));
 sky130_fd_sc_hd__nand2_1 _21081_ (.A(net298),
    .B(_08596_),
    .Y(_08721_));
 sky130_fd_sc_hd__o311ai_0 _21082_ (.A1(_12906_),
    .A2(net298),
    .A3(_08720_),
    .B1(_08721_),
    .C1(_12904_),
    .Y(_08722_));
 sky130_fd_sc_hd__o311ai_2 _21083_ (.A1(_08619_),
    .A2(_08673_),
    .A3(_08715_),
    .B1(_08719_),
    .C1(_08722_),
    .Y(_08723_));
 sky130_fd_sc_hd__a21o_1 _21084_ (.A1(_08350_),
    .A2(_08723_),
    .B1(net357),
    .X(_01009_));
 sky130_fd_sc_hd__nor2_1 _21085_ (.A(_12901_),
    .B(_08581_),
    .Y(_08724_));
 sky130_fd_sc_hd__o22ai_1 _21086_ (.A1(_08573_),
    .A2(_08608_),
    .B1(_08670_),
    .B2(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__a21oi_1 _21087_ (.A1(_12906_),
    .A2(_08607_),
    .B1(_12901_),
    .Y(_08726_));
 sky130_fd_sc_hd__nor3_1 _21088_ (.A(_12904_),
    .B(net539),
    .C(_08692_),
    .Y(_08727_));
 sky130_fd_sc_hd__a221oi_1 _21089_ (.A1(net539),
    .A2(_08692_),
    .B1(_08694_),
    .B2(_08726_),
    .C1(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21oi_1 _21090_ (.A1(_08591_),
    .A2(_08725_),
    .B1(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__o21bai_1 _21091_ (.A1(_08578_),
    .A2(_08729_),
    .B1_N(net357),
    .Y(_01010_));
 sky130_fd_sc_hd__nor2_1 _21092_ (.A(_12902_),
    .B(net298),
    .Y(_08730_));
 sky130_fd_sc_hd__a211oi_1 _21093_ (.A1(net298),
    .A2(_08660_),
    .B1(_08596_),
    .C1(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__nor2_2 _21094_ (.A(_08582_),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__nor2_1 _21095_ (.A(_08631_),
    .B(_08647_),
    .Y(_08733_));
 sky130_fd_sc_hd__nor2_1 _21096_ (.A(_08573_),
    .B(_08648_),
    .Y(_08734_));
 sky130_fd_sc_hd__o21ai_1 _21097_ (.A1(_08733_),
    .A2(_08734_),
    .B1(net300),
    .Y(_08735_));
 sky130_fd_sc_hd__a41oi_2 _21098_ (.A1(_08658_),
    .A2(_08679_),
    .A3(_08732_),
    .A4(_08735_),
    .B1(net292),
    .Y(_01011_));
 sky130_fd_sc_hd__a21oi_2 _21099_ (.A1(_08591_),
    .A2(_08581_),
    .B1(_12904_),
    .Y(_08736_));
 sky130_fd_sc_hd__o21ai_0 _21100_ (.A1(_08692_),
    .A2(_08736_),
    .B1(_08684_),
    .Y(_08737_));
 sky130_fd_sc_hd__a21oi_1 _21101_ (.A1(_08636_),
    .A2(_08656_),
    .B1(net300),
    .Y(_08738_));
 sky130_fd_sc_hd__a21oi_1 _21102_ (.A1(_12901_),
    .A2(_08608_),
    .B1(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__o21ai_0 _21103_ (.A1(net346),
    .A2(_08576_),
    .B1(_08659_),
    .Y(_08740_));
 sky130_fd_sc_hd__a21oi_1 _21104_ (.A1(_09857_),
    .A2(_08740_),
    .B1(_08733_),
    .Y(_08741_));
 sky130_fd_sc_hd__o22ai_2 _21105_ (.A1(net539),
    .A2(_08739_),
    .B1(_08741_),
    .B2(_08599_),
    .Y(_08742_));
 sky130_fd_sc_hd__nor2_1 _21106_ (.A(_08737_),
    .B(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__nor2_2 _21107_ (.A(_08578_),
    .B(_08743_),
    .Y(_01012_));
 sky130_fd_sc_hd__o21ai_0 _21108_ (.A1(net347),
    .A2(_08651_),
    .B1(_08692_),
    .Y(_08744_));
 sky130_fd_sc_hd__o21ai_0 _21109_ (.A1(net347),
    .A2(_08577_),
    .B1(_08632_),
    .Y(_08745_));
 sky130_fd_sc_hd__o21ai_0 _21110_ (.A1(net300),
    .A2(_08745_),
    .B1(_08595_),
    .Y(_08746_));
 sky130_fd_sc_hd__nand2_4 _21111_ (.A(net539),
    .B(net300),
    .Y(_08747_));
 sky130_fd_sc_hd__nand3_1 _21112_ (.A(net539),
    .B(net300),
    .C(_08593_),
    .Y(_08748_));
 sky130_fd_sc_hd__a21oi_1 _21113_ (.A1(_08611_),
    .A2(_08748_),
    .B1(_12901_),
    .Y(_08749_));
 sky130_fd_sc_hd__a311oi_1 _21114_ (.A1(_08747_),
    .A2(_08611_),
    .A3(_08631_),
    .B1(_08749_),
    .C1(_09857_),
    .Y(_08750_));
 sky130_fd_sc_hd__a221oi_1 _21115_ (.A1(_12906_),
    .A2(_08744_),
    .B1(_08746_),
    .B2(_09857_),
    .C1(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__o21bai_1 _21116_ (.A1(_08578_),
    .A2(_08751_),
    .B1_N(net540),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _21117_ (.A(_12906_),
    .B(_08599_),
    .Y(_08752_));
 sky130_fd_sc_hd__nand2_1 _21118_ (.A(_12902_),
    .B(net298),
    .Y(_08753_));
 sky130_fd_sc_hd__a31oi_1 _21119_ (.A1(_08576_),
    .A2(_08752_),
    .A3(_08753_),
    .B1(_08596_),
    .Y(_08754_));
 sky130_fd_sc_hd__a21oi_1 _21120_ (.A1(_08573_),
    .A2(_08694_),
    .B1(net339),
    .Y(_08755_));
 sky130_fd_sc_hd__a21oi_1 _21121_ (.A1(_12901_),
    .A2(_08685_),
    .B1(_08705_),
    .Y(_08756_));
 sky130_fd_sc_hd__nor2_1 _21122_ (.A(_08599_),
    .B(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__nor3_1 _21123_ (.A(_08754_),
    .B(_08755_),
    .C(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__o21bai_1 _21124_ (.A1(_08578_),
    .A2(_08758_),
    .B1_N(net357),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _21125_ (.A(_08589_),
    .B(_08618_),
    .Y(_08759_));
 sky130_fd_sc_hd__o21ai_0 _21126_ (.A1(_12904_),
    .A2(net298),
    .B1(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__a21oi_1 _21127_ (.A1(_12901_),
    .A2(net345),
    .B1(_12902_),
    .Y(_08761_));
 sky130_fd_sc_hd__nor2_1 _21128_ (.A(_08609_),
    .B(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__a21oi_1 _21129_ (.A1(_08652_),
    .A2(_08686_),
    .B1(_08578_),
    .Y(_08763_));
 sky130_fd_sc_hd__o21ai_0 _21130_ (.A1(_12904_),
    .A2(_08762_),
    .B1(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__a21oi_1 _21131_ (.A1(net339),
    .A2(_08760_),
    .B1(_08764_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand3_1 _21132_ (.A(_12906_),
    .B(_08607_),
    .C(_08591_),
    .Y(_08765_));
 sky130_fd_sc_hd__nand2_4 _21133_ (.A(_08607_),
    .B(net347),
    .Y(_08766_));
 sky130_fd_sc_hd__o22ai_1 _21134_ (.A1(_12904_),
    .A2(net347),
    .B1(_08766_),
    .B2(_12906_),
    .Y(_08767_));
 sky130_fd_sc_hd__nor2_1 _21135_ (.A(_12901_),
    .B(_08599_),
    .Y(_08768_));
 sky130_fd_sc_hd__a32oi_1 _21136_ (.A1(_08608_),
    .A2(_08716_),
    .A3(_08765_),
    .B1(_08767_),
    .B2(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__nor3_1 _21137_ (.A(_08582_),
    .B(_08706_),
    .C(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__a21oi_1 _21138_ (.A1(_08703_),
    .A2(_08770_),
    .B1(net292),
    .Y(_01016_));
 sky130_fd_sc_hd__a21oi_1 _21139_ (.A1(_12904_),
    .A2(net339),
    .B1(_12906_),
    .Y(_08771_));
 sky130_fd_sc_hd__nand2_1 _21140_ (.A(_12904_),
    .B(_08673_),
    .Y(_08772_));
 sky130_fd_sc_hd__o221ai_1 _21141_ (.A1(_08607_),
    .A2(_08589_),
    .B1(_08771_),
    .B2(net347),
    .C1(_08772_),
    .Y(_08773_));
 sky130_fd_sc_hd__o21ai_0 _21142_ (.A1(_08591_),
    .A2(_08692_),
    .B1(_08651_),
    .Y(_08774_));
 sky130_fd_sc_hd__a22oi_1 _21143_ (.A1(_08599_),
    .A2(_08773_),
    .B1(_08774_),
    .B2(_12901_),
    .Y(_08775_));
 sky130_fd_sc_hd__o21bai_1 _21144_ (.A1(_08578_),
    .A2(_08775_),
    .B1_N(net540),
    .Y(_01017_));
 sky130_fd_sc_hd__nor2_2 _21145_ (.A(net339),
    .B(net347),
    .Y(_08776_));
 sky130_fd_sc_hd__nor2_2 _21146_ (.A(_08607_),
    .B(net298),
    .Y(_08777_));
 sky130_fd_sc_hd__nor2_1 _21147_ (.A(_08591_),
    .B(_08633_),
    .Y(_08778_));
 sky130_fd_sc_hd__nor2_1 _21148_ (.A(_12904_),
    .B(_08607_),
    .Y(_08779_));
 sky130_fd_sc_hd__o21ai_0 _21149_ (.A1(_08599_),
    .A2(_08779_),
    .B1(_08686_),
    .Y(_08780_));
 sky130_fd_sc_hd__o21ai_0 _21150_ (.A1(_12902_),
    .A2(_08778_),
    .B1(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__o21ai_0 _21151_ (.A1(_08612_),
    .A2(_08776_),
    .B1(_12906_),
    .Y(_08782_));
 sky130_fd_sc_hd__o311ai_0 _21152_ (.A1(_08609_),
    .A2(_08777_),
    .A3(_08781_),
    .B1(_08782_),
    .C1(_08732_),
    .Y(_08783_));
 sky130_fd_sc_hd__a21oi_1 _21153_ (.A1(_12904_),
    .A2(_08776_),
    .B1(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__nor2_1 _21154_ (.A(net292),
    .B(_08784_),
    .Y(_01018_));
 sky130_fd_sc_hd__nor2_1 _21155_ (.A(_08631_),
    .B(_08766_),
    .Y(_08785_));
 sky130_fd_sc_hd__a21oi_1 _21156_ (.A1(net300),
    .A2(_08649_),
    .B1(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__o21ai_0 _21157_ (.A1(_08633_),
    .A2(_08639_),
    .B1(_12901_),
    .Y(_08787_));
 sky130_fd_sc_hd__a31oi_1 _21158_ (.A1(_08658_),
    .A2(_08786_),
    .A3(_08787_),
    .B1(_08578_),
    .Y(_01019_));
 sky130_fd_sc_hd__a22oi_1 _21159_ (.A1(_12904_),
    .A2(_08633_),
    .B1(_08697_),
    .B2(_12902_),
    .Y(_08788_));
 sky130_fd_sc_hd__o21ai_0 _21160_ (.A1(net347),
    .A2(_08670_),
    .B1(_08766_),
    .Y(_08789_));
 sky130_fd_sc_hd__a22oi_1 _21161_ (.A1(_12906_),
    .A2(_08652_),
    .B1(_08789_),
    .B2(_12901_),
    .Y(_08790_));
 sky130_fd_sc_hd__o21ai_0 _21162_ (.A1(net347),
    .A2(_08788_),
    .B1(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__a221oi_1 _21163_ (.A1(_12906_),
    .A2(net298),
    .B1(_08663_),
    .B2(_12904_),
    .C1(_08791_),
    .Y(_08792_));
 sky130_fd_sc_hd__nor2_1 _21164_ (.A(_08578_),
    .B(_08792_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_1 _21165_ (.A(_08651_),
    .B(_08653_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand2_2 _21166_ (.A(_08747_),
    .B(_08611_),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_1 _21167_ (.A(_12906_),
    .B(_08697_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand2_1 _21168_ (.A(_12901_),
    .B(_08794_),
    .Y(_08796_));
 sky130_fd_sc_hd__nor3_1 _21169_ (.A(net300),
    .B(_08631_),
    .C(_08766_),
    .Y(_08797_));
 sky130_fd_sc_hd__a31oi_1 _21170_ (.A1(_12904_),
    .A2(net539),
    .A3(_08696_),
    .B1(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__o2111ai_1 _21171_ (.A1(_08656_),
    .A2(_08794_),
    .B1(_08795_),
    .C1(_08796_),
    .D1(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__a21oi_1 _21172_ (.A1(_12902_),
    .A2(_08793_),
    .B1(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__o21bai_1 _21173_ (.A1(_08578_),
    .A2(_08800_),
    .B1_N(net540),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _21174_ (.A(_12901_),
    .B(_08652_),
    .Y(_08801_));
 sky130_fd_sc_hd__o21ai_0 _21175_ (.A1(_08652_),
    .A2(_08696_),
    .B1(_12906_),
    .Y(_08802_));
 sky130_fd_sc_hd__a21o_1 _21176_ (.A1(_08801_),
    .A2(_08802_),
    .B1(_08591_),
    .X(_08803_));
 sky130_fd_sc_hd__o21ai_0 _21177_ (.A1(_12901_),
    .A2(_08581_),
    .B1(_08663_),
    .Y(_08804_));
 sky130_fd_sc_hd__o22ai_1 _21178_ (.A1(_08589_),
    .A2(_08647_),
    .B1(_08685_),
    .B2(_08593_),
    .Y(_08805_));
 sky130_fd_sc_hd__nand2_1 _21179_ (.A(net298),
    .B(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__a31oi_1 _21180_ (.A1(_08803_),
    .A2(_08804_),
    .A3(_08806_),
    .B1(_08578_),
    .Y(_08807_));
 sky130_fd_sc_hd__or2_0 _21181_ (.A(net540),
    .B(_08807_),
    .X(_01022_));
 sky130_fd_sc_hd__a21oi_1 _21182_ (.A1(_12901_),
    .A2(_08591_),
    .B1(_09857_),
    .Y(_08808_));
 sky130_fd_sc_hd__o21ai_0 _21183_ (.A1(_08582_),
    .A2(_08611_),
    .B1(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__a31oi_2 _21184_ (.A1(_12906_),
    .A2(_08747_),
    .A3(_08611_),
    .B1(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__a22oi_1 _21185_ (.A1(_12901_),
    .A2(_08663_),
    .B1(_08655_),
    .B2(_12902_),
    .Y(_08811_));
 sky130_fd_sc_hd__nand3_1 _21186_ (.A(_09857_),
    .B(_08716_),
    .C(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__nor3b_4 _21187_ (.A(_08810_),
    .B(_08578_),
    .C_N(_08812_),
    .Y(_01023_));
 sky130_fd_sc_hd__nand2_1 _21188_ (.A(_12904_),
    .B(_08766_),
    .Y(_08813_));
 sky130_fd_sc_hd__a22oi_1 _21189_ (.A1(_12902_),
    .A2(_08776_),
    .B1(_08701_),
    .B2(_12901_),
    .Y(_08814_));
 sky130_fd_sc_hd__a21oi_1 _21190_ (.A1(_08813_),
    .A2(_08814_),
    .B1(_08599_),
    .Y(_08815_));
 sky130_fd_sc_hd__nand2_1 _21191_ (.A(_12902_),
    .B(_08639_),
    .Y(_08816_));
 sky130_fd_sc_hd__a21oi_1 _21192_ (.A1(_08796_),
    .A2(_08816_),
    .B1(_08607_),
    .Y(_08817_));
 sky130_fd_sc_hd__nor2_1 _21193_ (.A(_08815_),
    .B(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__o2111ai_1 _21194_ (.A1(_08692_),
    .A2(_08736_),
    .B1(_08818_),
    .C1(_08707_),
    .D1(_08577_),
    .Y(_08819_));
 sky130_fd_sc_hd__a21o_1 _21195_ (.A1(_08350_),
    .A2(_08819_),
    .B1(net540),
    .X(_01024_));
 sky130_fd_sc_hd__a21oi_1 _21196_ (.A1(_12902_),
    .A2(net298),
    .B1(_12904_),
    .Y(_08820_));
 sky130_fd_sc_hd__a21oi_1 _21197_ (.A1(_12906_),
    .A2(_08663_),
    .B1(_09857_),
    .Y(_08821_));
 sky130_fd_sc_hd__o21ai_0 _21198_ (.A1(_08591_),
    .A2(_08820_),
    .B1(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__a32oi_1 _21199_ (.A1(_12901_),
    .A2(net347),
    .A3(net298),
    .B1(_08812_),
    .B2(_08822_),
    .Y(_08823_));
 sky130_fd_sc_hd__a21oi_1 _21200_ (.A1(_08803_),
    .A2(_08823_),
    .B1(_08578_),
    .Y(_01025_));
 sky130_fd_sc_hd__a21oi_1 _21201_ (.A1(_12901_),
    .A2(net345),
    .B1(_12904_),
    .Y(_08824_));
 sky130_fd_sc_hd__nor2_1 _21202_ (.A(_08701_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__o211ai_1 _21203_ (.A1(_12906_),
    .A2(_08825_),
    .B1(_08647_),
    .C1(net298),
    .Y(_08826_));
 sky130_fd_sc_hd__nor2_1 _21204_ (.A(_12906_),
    .B(_08766_),
    .Y(_08827_));
 sky130_fd_sc_hd__a21oi_1 _21205_ (.A1(_08607_),
    .A2(_08603_),
    .B1(net345),
    .Y(_08828_));
 sky130_fd_sc_hd__or4_1 _21206_ (.A(net298),
    .B(_08827_),
    .C(_08779_),
    .D(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__a31oi_1 _21207_ (.A1(_08677_),
    .A2(_08826_),
    .A3(_08829_),
    .B1(net292),
    .Y(_01026_));
 sky130_fd_sc_hd__a21oi_1 _21208_ (.A1(_12901_),
    .A2(net298),
    .B1(_12902_),
    .Y(_08830_));
 sky130_fd_sc_hd__nor2_1 _21209_ (.A(net339),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__a21oi_1 _21210_ (.A1(_12906_),
    .A2(_08777_),
    .B1(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__a22oi_1 _21211_ (.A1(_12904_),
    .A2(_08777_),
    .B1(_08692_),
    .B2(_08705_),
    .Y(_08833_));
 sky130_fd_sc_hd__o211ai_1 _21212_ (.A1(net345),
    .A2(_08832_),
    .B1(_08833_),
    .C1(_08732_),
    .Y(_08834_));
 sky130_fd_sc_hd__a21o_4 _21213_ (.A1(_08350_),
    .A2(_08834_),
    .B1(net357),
    .X(_01027_));
 sky130_fd_sc_hd__a21oi_1 _21214_ (.A1(_12901_),
    .A2(net339),
    .B1(_12904_),
    .Y(_08835_));
 sky130_fd_sc_hd__nand2_1 _21215_ (.A(_12906_),
    .B(_08673_),
    .Y(_08836_));
 sky130_fd_sc_hd__o21ai_0 _21216_ (.A1(net345),
    .A2(_08835_),
    .B1(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__a21oi_1 _21217_ (.A1(_12906_),
    .A2(_08607_),
    .B1(_12904_),
    .Y(_08838_));
 sky130_fd_sc_hd__o21ai_0 _21218_ (.A1(_08652_),
    .A2(_08838_),
    .B1(_08602_),
    .Y(_08839_));
 sky130_fd_sc_hd__a21oi_1 _21219_ (.A1(_08602_),
    .A2(_08607_),
    .B1(net346),
    .Y(_08840_));
 sky130_fd_sc_hd__o221ai_1 _21220_ (.A1(_08607_),
    .A2(_08629_),
    .B1(_08840_),
    .B2(_12901_),
    .C1(_08766_),
    .Y(_08841_));
 sky130_fd_sc_hd__nor2_1 _21221_ (.A(_08599_),
    .B(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__a221oi_1 _21222_ (.A1(_08599_),
    .A2(_08837_),
    .B1(_08839_),
    .B2(net345),
    .C1(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__nor2_2 _21223_ (.A(_08578_),
    .B(_08843_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand2_1 _21224_ (.A(_12904_),
    .B(_08692_),
    .Y(_08844_));
 sky130_fd_sc_hd__a311o_1 _21225_ (.A1(_08602_),
    .A2(_08801_),
    .A3(_08844_),
    .B1(net347),
    .C1(_08696_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _21226_ (.A(net298),
    .B(_08576_),
    .Y(_08846_));
 sky130_fd_sc_hd__a2bb2oi_1 _21227_ (.A1_N(_12906_),
    .A2_N(_08846_),
    .B1(_08777_),
    .B2(_08576_),
    .Y(_08847_));
 sky130_fd_sc_hd__o21ai_0 _21228_ (.A1(_12902_),
    .A2(_08847_),
    .B1(_08778_),
    .Y(_08848_));
 sky130_fd_sc_hd__a31oi_1 _21229_ (.A1(_08684_),
    .A2(_08845_),
    .A3(_08848_),
    .B1(_08578_),
    .Y(_01029_));
 sky130_fd_sc_hd__a21oi_1 _21230_ (.A1(net539),
    .A2(net300),
    .B1(_08593_),
    .Y(_08849_));
 sky130_fd_sc_hd__o22ai_1 _21231_ (.A1(_12904_),
    .A2(_08655_),
    .B1(_08849_),
    .B2(_12901_),
    .Y(_08850_));
 sky130_fd_sc_hd__a21oi_1 _21232_ (.A1(_08602_),
    .A2(_08850_),
    .B1(_08622_),
    .Y(_08851_));
 sky130_fd_sc_hd__nor2_1 _21233_ (.A(net298),
    .B(_08736_),
    .Y(_08852_));
 sky130_fd_sc_hd__a21oi_1 _21234_ (.A1(_12901_),
    .A2(_08747_),
    .B1(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__a21oi_1 _21235_ (.A1(_12904_),
    .A2(net339),
    .B1(_12902_),
    .Y(_08854_));
 sky130_fd_sc_hd__o221ai_1 _21236_ (.A1(_08607_),
    .A2(_08853_),
    .B1(_08854_),
    .B2(_08747_),
    .C1(_08577_),
    .Y(_08855_));
 sky130_fd_sc_hd__a21oi_1 _21237_ (.A1(_08607_),
    .A2(_08851_),
    .B1(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__o21bai_1 _21238_ (.A1(_08320_),
    .A2(_08856_),
    .B1_N(net540),
    .Y(_01030_));
 sky130_fd_sc_hd__o21ai_0 _21239_ (.A1(_08609_),
    .A2(_08639_),
    .B1(_12902_),
    .Y(_08857_));
 sky130_fd_sc_hd__nand3_1 _21240_ (.A(_12904_),
    .B(_08599_),
    .C(_08647_),
    .Y(_08858_));
 sky130_fd_sc_hd__a21oi_1 _21241_ (.A1(_08681_),
    .A2(_08858_),
    .B1(_12901_),
    .Y(_08859_));
 sky130_fd_sc_hd__a21oi_1 _21242_ (.A1(_12901_),
    .A2(_08608_),
    .B1(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__xnor2_1 _21243_ (.A(_09857_),
    .B(_08794_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand2_1 _21244_ (.A(_12906_),
    .B(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__a31oi_2 _21245_ (.A1(_08857_),
    .A2(_08860_),
    .A3(_08862_),
    .B1(net292),
    .Y(_01031_));
 sky130_fd_sc_hd__nor2_1 _21246_ (.A(_08659_),
    .B(_08652_),
    .Y(_08863_));
 sky130_fd_sc_hd__a2111oi_0 _21247_ (.A1(_12904_),
    .A2(_08696_),
    .B1(_08791_),
    .C1(_08863_),
    .D1(_08582_),
    .Y(_08864_));
 sky130_fd_sc_hd__nor2_1 _21248_ (.A(net292),
    .B(_08864_),
    .Y(_01032_));
 sky130_fd_sc_hd__nor2_1 _21249_ (.A(net540),
    .B(_08258_),
    .Y(_01033_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_921 ();
 sky130_fd_sc_hd__nand2_8 _21251_ (.A(_09745_),
    .B(_04784_),
    .Y(_08866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_920 ();
 sky130_fd_sc_hd__nor2_1 _21253_ (.A(_04790_),
    .B(_08866_),
    .Y(_01034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_919 ();
 sky130_fd_sc_hd__nor2_1 _21255_ (.A(_04871_),
    .B(_08866_),
    .Y(_01035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_918 ();
 sky130_fd_sc_hd__nor2_1 _21257_ (.A(_04883_),
    .B(_08866_),
    .Y(_01036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_917 ();
 sky130_fd_sc_hd__nor2_1 _21259_ (.A(_04892_),
    .B(_08866_),
    .Y(_01037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_916 ();
 sky130_fd_sc_hd__nor2_1 _21261_ (.A(_04899_),
    .B(_08866_),
    .Y(_01038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_915 ();
 sky130_fd_sc_hd__nor2_1 _21263_ (.A(_04906_),
    .B(_08866_),
    .Y(_01039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_914 ();
 sky130_fd_sc_hd__nor2_1 _21265_ (.A(_04913_),
    .B(_08866_),
    .Y(_01040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_913 ();
 sky130_fd_sc_hd__nor2_1 _21267_ (.A(_04923_),
    .B(_08866_),
    .Y(_01041_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_912 ();
 sky130_fd_sc_hd__nor2_1 _21269_ (.A(_04932_),
    .B(_08866_),
    .Y(_01042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_911 ();
 sky130_fd_sc_hd__nor2_1 _21271_ (.A(_04939_),
    .B(_08866_),
    .Y(_01043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_909 ();
 sky130_fd_sc_hd__nor2_1 _21274_ (.A(_04951_),
    .B(_08866_),
    .Y(_01044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_908 ();
 sky130_fd_sc_hd__nor2_1 _21276_ (.A(_04794_),
    .B(_08866_),
    .Y(_01045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_907 ();
 sky130_fd_sc_hd__nor2_1 _21278_ (.A(_04960_),
    .B(_08866_),
    .Y(_01046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_906 ();
 sky130_fd_sc_hd__nor2_1 _21280_ (.A(_04974_),
    .B(_08866_),
    .Y(_01047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_905 ();
 sky130_fd_sc_hd__nor2_1 _21282_ (.A(_04984_),
    .B(_08866_),
    .Y(_01048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_904 ();
 sky130_fd_sc_hd__nor2_1 _21284_ (.A(_04990_),
    .B(_08866_),
    .Y(_01049_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_903 ();
 sky130_fd_sc_hd__nor2_1 _21286_ (.A(_05000_),
    .B(_08866_),
    .Y(_01050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_902 ();
 sky130_fd_sc_hd__nor2_1 _21288_ (.A(_05011_),
    .B(_08866_),
    .Y(_01051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_901 ();
 sky130_fd_sc_hd__nor2_1 _21290_ (.A(_05020_),
    .B(_08866_),
    .Y(_01052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_900 ();
 sky130_fd_sc_hd__nor2_1 _21292_ (.A(_05029_),
    .B(_08866_),
    .Y(_01053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_898 ();
 sky130_fd_sc_hd__nor2_1 _21295_ (.A(_05035_),
    .B(_08866_),
    .Y(_01054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_897 ();
 sky130_fd_sc_hd__nor2_1 _21297_ (.A(net1143),
    .B(_08866_),
    .Y(_01055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_896 ();
 sky130_fd_sc_hd__nor2_1 _21299_ (.A(_04801_),
    .B(_08866_),
    .Y(_01056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_895 ();
 sky130_fd_sc_hd__nor2_1 _21301_ (.A(_05060_),
    .B(_08866_),
    .Y(_01057_));
 sky130_fd_sc_hd__o21bai_1 _21302_ (.A1(_05107_),
    .A2(_05109_),
    .B1_N(_13104_),
    .Y(_08893_));
 sky130_fd_sc_hd__xnor2_1 _21303_ (.A(_05103_),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__mux2i_4 _21304_ (.A0(\w[62][31] ),
    .A1(_08894_),
    .S(net348),
    .Y(_08895_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_894 ();
 sky130_fd_sc_hd__nor2_1 _21306_ (.A(_08866_),
    .B(_08895_),
    .Y(_01058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_893 ();
 sky130_fd_sc_hd__nor2_1 _21308_ (.A(_04808_),
    .B(_08866_),
    .Y(_01059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_892 ();
 sky130_fd_sc_hd__nor2_1 _21310_ (.A(_04817_),
    .B(_08866_),
    .Y(_01060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_891 ();
 sky130_fd_sc_hd__nor2_1 _21312_ (.A(_04826_),
    .B(_08866_),
    .Y(_01061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_890 ();
 sky130_fd_sc_hd__nor2_1 _21314_ (.A(_04834_),
    .B(_08866_),
    .Y(_01062_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_889 ();
 sky130_fd_sc_hd__nor2_1 _21316_ (.A(_04843_),
    .B(_08866_),
    .Y(_01063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_888 ();
 sky130_fd_sc_hd__nor2_1 _21318_ (.A(_04852_),
    .B(_08866_),
    .Y(_01064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_887 ();
 sky130_fd_sc_hd__nor2_1 _21320_ (.A(_04860_),
    .B(_08866_),
    .Y(_01065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_886 ();
 sky130_fd_sc_hd__nand2_8 _21322_ (.A(_09794_),
    .B(_05115_),
    .Y(_08905_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_885 ();
 sky130_fd_sc_hd__nor2_1 _21324_ (.A(_05118_),
    .B(_08905_),
    .Y(_01066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_884 ();
 sky130_fd_sc_hd__nor2_1 _21326_ (.A(_05192_),
    .B(_08905_),
    .Y(_01067_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_883 ();
 sky130_fd_sc_hd__nor2_1 _21328_ (.A(_05204_),
    .B(_08905_),
    .Y(_01068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_882 ();
 sky130_fd_sc_hd__nor2_1 _21330_ (.A(_05214_),
    .B(_08905_),
    .Y(_01069_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_881 ();
 sky130_fd_sc_hd__nor2_1 _21332_ (.A(_05221_),
    .B(_08905_),
    .Y(_01070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_880 ();
 sky130_fd_sc_hd__nor2_1 _21334_ (.A(net1136),
    .B(_08905_),
    .Y(_01071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_879 ();
 sky130_fd_sc_hd__nor2_1 _21336_ (.A(_05238_),
    .B(_08905_),
    .Y(_01072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_878 ();
 sky130_fd_sc_hd__nor2_1 _21338_ (.A(net1135),
    .B(_08905_),
    .Y(_01073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_877 ();
 sky130_fd_sc_hd__nor2_1 _21340_ (.A(_05258_),
    .B(_08905_),
    .Y(_01074_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_876 ();
 sky130_fd_sc_hd__nor2_1 _21342_ (.A(_05267_),
    .B(_08905_),
    .Y(_01075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_874 ();
 sky130_fd_sc_hd__nor2_1 _21345_ (.A(_05280_),
    .B(_08905_),
    .Y(_01076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_873 ();
 sky130_fd_sc_hd__nor2_1 _21347_ (.A(_05122_),
    .B(_08905_),
    .Y(_01077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_872 ();
 sky130_fd_sc_hd__nor2_1 _21349_ (.A(_05291_),
    .B(_08905_),
    .Y(_01078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_871 ();
 sky130_fd_sc_hd__nor2_1 _21351_ (.A(_05301_),
    .B(_08905_),
    .Y(_01079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_870 ();
 sky130_fd_sc_hd__nor2_1 _21353_ (.A(_05309_),
    .B(_08905_),
    .Y(_01080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_869 ();
 sky130_fd_sc_hd__nor2_1 _21355_ (.A(_05320_),
    .B(_08905_),
    .Y(_01081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_868 ();
 sky130_fd_sc_hd__nor2_1 _21357_ (.A(net1137),
    .B(_08905_),
    .Y(_01082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_867 ();
 sky130_fd_sc_hd__nor2_1 _21359_ (.A(_05339_),
    .B(_08905_),
    .Y(_01083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_866 ();
 sky130_fd_sc_hd__nor2_1 _21361_ (.A(_05347_),
    .B(_08905_),
    .Y(_01084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_865 ();
 sky130_fd_sc_hd__nor2_1 _21363_ (.A(net538),
    .B(_08905_),
    .Y(_01085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_863 ();
 sky130_fd_sc_hd__nor2_1 _21366_ (.A(net1142),
    .B(_08905_),
    .Y(_01086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_862 ();
 sky130_fd_sc_hd__nor2_1 _21368_ (.A(_05380_),
    .B(_08905_),
    .Y(_01087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_861 ();
 sky130_fd_sc_hd__nor2_1 _21370_ (.A(_05126_),
    .B(_08905_),
    .Y(_01088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_860 ();
 sky130_fd_sc_hd__nor2_1 _21372_ (.A(net1129),
    .B(_08905_),
    .Y(_01089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_859 ();
 sky130_fd_sc_hd__nor2_1 _21374_ (.A(net1042),
    .B(_08905_),
    .Y(_01090_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_858 ();
 sky130_fd_sc_hd__nor2_1 _21376_ (.A(_05132_),
    .B(_08905_),
    .Y(_01091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_857 ();
 sky130_fd_sc_hd__nor2_1 _21378_ (.A(_05140_),
    .B(_08905_),
    .Y(_01092_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_856 ();
 sky130_fd_sc_hd__nor2_1 _21380_ (.A(_05149_),
    .B(_08905_),
    .Y(_01093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_855 ();
 sky130_fd_sc_hd__nor2_1 _21382_ (.A(_05157_),
    .B(_08905_),
    .Y(_01094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_854 ();
 sky130_fd_sc_hd__nor2_1 _21384_ (.A(_05166_),
    .B(_08905_),
    .Y(_01095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_853 ();
 sky130_fd_sc_hd__nor2_1 _21386_ (.A(_05173_),
    .B(_08905_),
    .Y(_01096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_852 ();
 sky130_fd_sc_hd__nor2_1 _21388_ (.A(_05183_),
    .B(_08905_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_8 _21389_ (.A(_09745_),
    .B(_05433_),
    .Y(_08940_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_851 ();
 sky130_fd_sc_hd__nor2_1 _21391_ (.A(_04790_),
    .B(_08940_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_1 _21392_ (.A(_04871_),
    .B(_08940_),
    .Y(_01099_));
 sky130_fd_sc_hd__nor2_1 _21393_ (.A(_04883_),
    .B(_08940_),
    .Y(_01100_));
 sky130_fd_sc_hd__nor2_1 _21394_ (.A(_04892_),
    .B(_08940_),
    .Y(_01101_));
 sky130_fd_sc_hd__nor2_1 _21395_ (.A(_04899_),
    .B(_08940_),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_1 _21396_ (.A(_04906_),
    .B(_08940_),
    .Y(_01103_));
 sky130_fd_sc_hd__nor2_1 _21397_ (.A(_04913_),
    .B(_08940_),
    .Y(_01104_));
 sky130_fd_sc_hd__nor2_1 _21398_ (.A(_04923_),
    .B(_08940_),
    .Y(_01105_));
 sky130_fd_sc_hd__nor2_1 _21399_ (.A(_04932_),
    .B(_08940_),
    .Y(_01106_));
 sky130_fd_sc_hd__nor2_1 _21400_ (.A(_04939_),
    .B(_08940_),
    .Y(_01107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_850 ();
 sky130_fd_sc_hd__nor2_1 _21402_ (.A(_04951_),
    .B(_08940_),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _21403_ (.A(_04794_),
    .B(_08940_),
    .Y(_01109_));
 sky130_fd_sc_hd__nor2_1 _21404_ (.A(_04960_),
    .B(_08940_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2_1 _21405_ (.A(_04974_),
    .B(_08940_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_1 _21406_ (.A(_04984_),
    .B(_08940_),
    .Y(_01112_));
 sky130_fd_sc_hd__nor2_1 _21407_ (.A(_04990_),
    .B(_08940_),
    .Y(_01113_));
 sky130_fd_sc_hd__nor2_1 _21408_ (.A(net1139),
    .B(_08940_),
    .Y(_01114_));
 sky130_fd_sc_hd__nor2_1 _21409_ (.A(_05011_),
    .B(_08940_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _21410_ (.A(_05020_),
    .B(_08940_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor2_1 _21411_ (.A(_05029_),
    .B(_08940_),
    .Y(_01117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_849 ();
 sky130_fd_sc_hd__nor2_1 _21413_ (.A(_05035_),
    .B(_08940_),
    .Y(_01118_));
 sky130_fd_sc_hd__nor2_1 _21414_ (.A(_05044_),
    .B(_08940_),
    .Y(_01119_));
 sky130_fd_sc_hd__nor2_1 _21415_ (.A(_04801_),
    .B(_08940_),
    .Y(_01120_));
 sky130_fd_sc_hd__nor2_1 _21416_ (.A(_05060_),
    .B(_08940_),
    .Y(_01121_));
 sky130_fd_sc_hd__nor2_1 _21417_ (.A(_08895_),
    .B(_08940_),
    .Y(_01122_));
 sky130_fd_sc_hd__nor2_1 _21418_ (.A(_04808_),
    .B(_08940_),
    .Y(_01123_));
 sky130_fd_sc_hd__nor2_1 _21419_ (.A(_04817_),
    .B(_08940_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _21420_ (.A(_04826_),
    .B(_08940_),
    .Y(_01125_));
 sky130_fd_sc_hd__nor2_1 _21421_ (.A(_04834_),
    .B(_08940_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_1 _21422_ (.A(_04843_),
    .B(_08940_),
    .Y(_01127_));
 sky130_fd_sc_hd__nor2_1 _21423_ (.A(_04852_),
    .B(_08940_),
    .Y(_01128_));
 sky130_fd_sc_hd__nor2_1 _21424_ (.A(_04860_),
    .B(_08940_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_8 _21425_ (.A(_09794_),
    .B(_05474_),
    .Y(_08944_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_848 ();
 sky130_fd_sc_hd__nor2_1 _21427_ (.A(_05118_),
    .B(_08944_),
    .Y(_01130_));
 sky130_fd_sc_hd__nor2_1 _21428_ (.A(_05192_),
    .B(_08944_),
    .Y(_01131_));
 sky130_fd_sc_hd__nor2_1 _21429_ (.A(_05204_),
    .B(_08944_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_1 _21430_ (.A(_05214_),
    .B(_08944_),
    .Y(_01133_));
 sky130_fd_sc_hd__nor2_1 _21431_ (.A(_05221_),
    .B(_08944_),
    .Y(_01134_));
 sky130_fd_sc_hd__nor2_1 _21432_ (.A(net1136),
    .B(_08944_),
    .Y(_01135_));
 sky130_fd_sc_hd__nor2_1 _21433_ (.A(_05238_),
    .B(_08944_),
    .Y(_01136_));
 sky130_fd_sc_hd__nor2_1 _21434_ (.A(_05247_),
    .B(_08944_),
    .Y(_01137_));
 sky130_fd_sc_hd__nor2_1 _21435_ (.A(_05258_),
    .B(_08944_),
    .Y(_01138_));
 sky130_fd_sc_hd__nor2_1 _21436_ (.A(net1102),
    .B(_08944_),
    .Y(_01139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_847 ();
 sky130_fd_sc_hd__nor2_1 _21438_ (.A(_05280_),
    .B(_08944_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _21439_ (.A(_05122_),
    .B(_08944_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _21440_ (.A(_05291_),
    .B(_08944_),
    .Y(_01142_));
 sky130_fd_sc_hd__nor2_1 _21441_ (.A(_05301_),
    .B(_08944_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_1 _21442_ (.A(_05309_),
    .B(_08944_),
    .Y(_01144_));
 sky130_fd_sc_hd__nor2_1 _21443_ (.A(_05320_),
    .B(_08944_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _21444_ (.A(net1137),
    .B(_08944_),
    .Y(_01146_));
 sky130_fd_sc_hd__nor2_1 _21445_ (.A(_05339_),
    .B(_08944_),
    .Y(_01147_));
 sky130_fd_sc_hd__nor2_1 _21446_ (.A(_05347_),
    .B(_08944_),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_1 _21447_ (.A(net538),
    .B(_08944_),
    .Y(_01149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_846 ();
 sky130_fd_sc_hd__nor2_1 _21449_ (.A(net1101),
    .B(_08944_),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_1 _21450_ (.A(_05380_),
    .B(_08944_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _21451_ (.A(_05126_),
    .B(_08944_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor2_1 _21452_ (.A(net1129),
    .B(_08944_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor2_1 _21453_ (.A(net1042),
    .B(_08944_),
    .Y(_01154_));
 sky130_fd_sc_hd__nor2_1 _21454_ (.A(_05132_),
    .B(_08944_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _21455_ (.A(_05140_),
    .B(_08944_),
    .Y(_01156_));
 sky130_fd_sc_hd__nor2_1 _21456_ (.A(_05149_),
    .B(_08944_),
    .Y(_01157_));
 sky130_fd_sc_hd__nor2_1 _21457_ (.A(_05157_),
    .B(_08944_),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _21458_ (.A(_05166_),
    .B(_08944_),
    .Y(_01159_));
 sky130_fd_sc_hd__nor2_1 _21459_ (.A(_05173_),
    .B(_08944_),
    .Y(_01160_));
 sky130_fd_sc_hd__nor2_1 _21460_ (.A(_05183_),
    .B(_08944_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2_8 _21461_ (.A(_09745_),
    .B(_05516_),
    .Y(_08948_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_845 ();
 sky130_fd_sc_hd__nor2_1 _21463_ (.A(_04790_),
    .B(_08948_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_1 _21464_ (.A(_04871_),
    .B(_08948_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_1 _21465_ (.A(_04883_),
    .B(_08948_),
    .Y(_01164_));
 sky130_fd_sc_hd__nor2_1 _21466_ (.A(_04892_),
    .B(_08948_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _21467_ (.A(_04899_),
    .B(_08948_),
    .Y(_01166_));
 sky130_fd_sc_hd__nor2_1 _21468_ (.A(_04906_),
    .B(_08948_),
    .Y(_01167_));
 sky130_fd_sc_hd__nor2_1 _21469_ (.A(_04913_),
    .B(_08948_),
    .Y(_01168_));
 sky130_fd_sc_hd__nor2_1 _21470_ (.A(_04923_),
    .B(_08948_),
    .Y(_01169_));
 sky130_fd_sc_hd__nor2_1 _21471_ (.A(_04932_),
    .B(_08948_),
    .Y(_01170_));
 sky130_fd_sc_hd__nor2_1 _21472_ (.A(_04939_),
    .B(_08948_),
    .Y(_01171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_844 ();
 sky130_fd_sc_hd__nor2_1 _21474_ (.A(_04951_),
    .B(_08948_),
    .Y(_01172_));
 sky130_fd_sc_hd__nor2_1 _21475_ (.A(_04794_),
    .B(_08948_),
    .Y(_01173_));
 sky130_fd_sc_hd__nor2_1 _21476_ (.A(_04960_),
    .B(_08948_),
    .Y(_01174_));
 sky130_fd_sc_hd__nor2_1 _21477_ (.A(_04974_),
    .B(_08948_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor2_1 _21478_ (.A(_04984_),
    .B(_08948_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2_1 _21479_ (.A(_04990_),
    .B(_08948_),
    .Y(_01177_));
 sky130_fd_sc_hd__nor2_1 _21480_ (.A(_05000_),
    .B(_08948_),
    .Y(_01178_));
 sky130_fd_sc_hd__nor2_1 _21481_ (.A(_05011_),
    .B(_08948_),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_1 _21482_ (.A(_05020_),
    .B(_08948_),
    .Y(_01180_));
 sky130_fd_sc_hd__nor2_1 _21483_ (.A(_05029_),
    .B(_08948_),
    .Y(_01181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_843 ();
 sky130_fd_sc_hd__nor2_1 _21485_ (.A(net1138),
    .B(_08948_),
    .Y(_01182_));
 sky130_fd_sc_hd__nor2_1 _21486_ (.A(_05044_),
    .B(_08948_),
    .Y(_01183_));
 sky130_fd_sc_hd__nor2_1 _21487_ (.A(_04801_),
    .B(_08948_),
    .Y(_01184_));
 sky130_fd_sc_hd__nor2_1 _21488_ (.A(_05060_),
    .B(_08948_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_1 _21489_ (.A(_08895_),
    .B(_08948_),
    .Y(_01186_));
 sky130_fd_sc_hd__nor2_1 _21490_ (.A(_04808_),
    .B(_08948_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_1 _21491_ (.A(_04817_),
    .B(_08948_),
    .Y(_01188_));
 sky130_fd_sc_hd__nor2_1 _21492_ (.A(_04826_),
    .B(_08948_),
    .Y(_01189_));
 sky130_fd_sc_hd__nor2_1 _21493_ (.A(_04834_),
    .B(_08948_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _21494_ (.A(_04843_),
    .B(_08948_),
    .Y(_01191_));
 sky130_fd_sc_hd__nor2_1 _21495_ (.A(_04852_),
    .B(_08948_),
    .Y(_01192_));
 sky130_fd_sc_hd__nor2_1 _21496_ (.A(_04860_),
    .B(_08948_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_8 _21497_ (.A(_09794_),
    .B(_05557_),
    .Y(_08952_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_842 ();
 sky130_fd_sc_hd__nor2_1 _21499_ (.A(_05118_),
    .B(_08952_),
    .Y(_01194_));
 sky130_fd_sc_hd__nor2_1 _21500_ (.A(_05192_),
    .B(_08952_),
    .Y(_01195_));
 sky130_fd_sc_hd__nor2_1 _21501_ (.A(_05204_),
    .B(_08952_),
    .Y(_01196_));
 sky130_fd_sc_hd__nor2_1 _21502_ (.A(_05214_),
    .B(_08952_),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_1 _21503_ (.A(_05221_),
    .B(_08952_),
    .Y(_01198_));
 sky130_fd_sc_hd__nor2_1 _21504_ (.A(_05228_),
    .B(_08952_),
    .Y(_01199_));
 sky130_fd_sc_hd__nor2_1 _21505_ (.A(_05238_),
    .B(_08952_),
    .Y(_01200_));
 sky130_fd_sc_hd__nor2_1 _21506_ (.A(net1135),
    .B(_08952_),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _21507_ (.A(_05258_),
    .B(_08952_),
    .Y(_01202_));
 sky130_fd_sc_hd__nor2_1 _21508_ (.A(_05267_),
    .B(_08952_),
    .Y(_01203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_841 ();
 sky130_fd_sc_hd__nor2_1 _21510_ (.A(_05280_),
    .B(_08952_),
    .Y(_01204_));
 sky130_fd_sc_hd__nor2_1 _21511_ (.A(_05122_),
    .B(_08952_),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_1 _21512_ (.A(_05291_),
    .B(_08952_),
    .Y(_01206_));
 sky130_fd_sc_hd__nor2_1 _21513_ (.A(_05301_),
    .B(_08952_),
    .Y(_01207_));
 sky130_fd_sc_hd__nor2_1 _21514_ (.A(_05309_),
    .B(_08952_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _21515_ (.A(_05320_),
    .B(_08952_),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_1 _21516_ (.A(net1100),
    .B(_08952_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor2_1 _21517_ (.A(_05339_),
    .B(_08952_),
    .Y(_01211_));
 sky130_fd_sc_hd__nor2_1 _21518_ (.A(_05347_),
    .B(_08952_),
    .Y(_01212_));
 sky130_fd_sc_hd__nor2_1 _21519_ (.A(net538),
    .B(_08952_),
    .Y(_01213_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_840 ();
 sky130_fd_sc_hd__nor2_1 _21521_ (.A(net1101),
    .B(_08952_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_1 _21522_ (.A(_05380_),
    .B(_08952_),
    .Y(_01215_));
 sky130_fd_sc_hd__nor2_1 _21523_ (.A(_05126_),
    .B(_08952_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_1 _21524_ (.A(net1129),
    .B(_08952_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _21525_ (.A(net1042),
    .B(_08952_),
    .Y(_01218_));
 sky130_fd_sc_hd__nor2_1 _21526_ (.A(_05132_),
    .B(_08952_),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_1 _21527_ (.A(_05140_),
    .B(_08952_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor2_1 _21528_ (.A(_05149_),
    .B(_08952_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _21529_ (.A(_05157_),
    .B(_08952_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_1 _21530_ (.A(_05166_),
    .B(_08952_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_1 _21531_ (.A(_05173_),
    .B(_08952_),
    .Y(_01224_));
 sky130_fd_sc_hd__nor2_1 _21532_ (.A(_05183_),
    .B(_08952_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_8 _21533_ (.A(_09745_),
    .B(_05598_),
    .Y(_08956_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_839 ();
 sky130_fd_sc_hd__nor2_1 _21535_ (.A(_04790_),
    .B(_08956_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _21536_ (.A(_04871_),
    .B(_08956_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor2_1 _21537_ (.A(_04883_),
    .B(_08956_),
    .Y(_01228_));
 sky130_fd_sc_hd__nor2_1 _21538_ (.A(_04892_),
    .B(_08956_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_1 _21539_ (.A(_04899_),
    .B(_08956_),
    .Y(_01230_));
 sky130_fd_sc_hd__nor2_1 _21540_ (.A(_04906_),
    .B(_08956_),
    .Y(_01231_));
 sky130_fd_sc_hd__nor2_1 _21541_ (.A(_04913_),
    .B(_08956_),
    .Y(_01232_));
 sky130_fd_sc_hd__nor2_1 _21542_ (.A(_04923_),
    .B(_08956_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_1 _21543_ (.A(_04932_),
    .B(_08956_),
    .Y(_01234_));
 sky130_fd_sc_hd__nor2_1 _21544_ (.A(_04939_),
    .B(_08956_),
    .Y(_01235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_838 ();
 sky130_fd_sc_hd__nor2_1 _21546_ (.A(_04951_),
    .B(_08956_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_1 _21547_ (.A(_04794_),
    .B(_08956_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _21548_ (.A(_04960_),
    .B(_08956_),
    .Y(_01238_));
 sky130_fd_sc_hd__nor2_1 _21549_ (.A(_04974_),
    .B(_08956_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _21550_ (.A(_04984_),
    .B(_08956_),
    .Y(_01240_));
 sky130_fd_sc_hd__nor2_1 _21551_ (.A(_04990_),
    .B(_08956_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_1 _21552_ (.A(_05000_),
    .B(_08956_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_1 _21553_ (.A(_05011_),
    .B(_08956_),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _21554_ (.A(_05020_),
    .B(_08956_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _21555_ (.A(_05029_),
    .B(_08956_),
    .Y(_01245_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_837 ();
 sky130_fd_sc_hd__nor2_1 _21557_ (.A(net1138),
    .B(_08956_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _21558_ (.A(_05044_),
    .B(_08956_),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_1 _21559_ (.A(_04801_),
    .B(_08956_),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _21560_ (.A(_05060_),
    .B(_08956_),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_1 _21561_ (.A(_08895_),
    .B(_08956_),
    .Y(_01250_));
 sky130_fd_sc_hd__nor2_1 _21562_ (.A(_04808_),
    .B(_08956_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor2_1 _21563_ (.A(_04817_),
    .B(_08956_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _21564_ (.A(_04826_),
    .B(_08956_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor2_1 _21565_ (.A(_04834_),
    .B(_08956_),
    .Y(_01254_));
 sky130_fd_sc_hd__nor2_1 _21566_ (.A(_04843_),
    .B(_08956_),
    .Y(_01255_));
 sky130_fd_sc_hd__nor2_1 _21567_ (.A(_04852_),
    .B(_08956_),
    .Y(_01256_));
 sky130_fd_sc_hd__nor2_1 _21568_ (.A(_04860_),
    .B(_08956_),
    .Y(_01257_));
 sky130_fd_sc_hd__or3_4 _21569_ (.A(net1043),
    .B(_09793_),
    .C(_09803_),
    .X(_08960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_835 ();
 sky130_fd_sc_hd__nor2_1 _21572_ (.A(_05118_),
    .B(_08960_),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _21573_ (.A(_05192_),
    .B(_08960_),
    .Y(_01259_));
 sky130_fd_sc_hd__nor2_1 _21574_ (.A(_05204_),
    .B(_08960_),
    .Y(_01260_));
 sky130_fd_sc_hd__nor2_1 _21575_ (.A(_05214_),
    .B(_08960_),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_1 _21576_ (.A(_05221_),
    .B(_08960_),
    .Y(_01262_));
 sky130_fd_sc_hd__nor2_1 _21577_ (.A(_05228_),
    .B(_08960_),
    .Y(_01263_));
 sky130_fd_sc_hd__nor2_1 _21578_ (.A(_05238_),
    .B(_08960_),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_1 _21579_ (.A(net1135),
    .B(_08960_),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _21580_ (.A(_05258_),
    .B(_08960_),
    .Y(_01266_));
 sky130_fd_sc_hd__nor2_1 _21581_ (.A(_05267_),
    .B(_08960_),
    .Y(_01267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_834 ();
 sky130_fd_sc_hd__nor2_1 _21583_ (.A(_05280_),
    .B(_08960_),
    .Y(_01268_));
 sky130_fd_sc_hd__nor2_1 _21584_ (.A(_05122_),
    .B(_08960_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_1 _21585_ (.A(_05291_),
    .B(_08960_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _21586_ (.A(_05301_),
    .B(_08960_),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_1 _21587_ (.A(_05309_),
    .B(_08960_),
    .Y(_01272_));
 sky130_fd_sc_hd__nor2_1 _21588_ (.A(_05320_),
    .B(_08960_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor2_1 _21589_ (.A(net1137),
    .B(_08960_),
    .Y(_01274_));
 sky130_fd_sc_hd__nor2_1 _21590_ (.A(_05339_),
    .B(_08960_),
    .Y(_01275_));
 sky130_fd_sc_hd__nor2_1 _21591_ (.A(_05347_),
    .B(_08960_),
    .Y(_01276_));
 sky130_fd_sc_hd__nor2_1 _21592_ (.A(net538),
    .B(_08960_),
    .Y(_01277_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_833 ();
 sky130_fd_sc_hd__nor2_1 _21594_ (.A(net1142),
    .B(_08960_),
    .Y(_01278_));
 sky130_fd_sc_hd__nor2_1 _21595_ (.A(_05380_),
    .B(_08960_),
    .Y(_01279_));
 sky130_fd_sc_hd__nor2_1 _21596_ (.A(_05126_),
    .B(_08960_),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_1 _21597_ (.A(net1134),
    .B(_08960_),
    .Y(_01281_));
 sky130_fd_sc_hd__nor2_1 _21598_ (.A(net1042),
    .B(_08960_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor2_1 _21599_ (.A(_05132_),
    .B(_08960_),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_1 _21600_ (.A(_05140_),
    .B(_08960_),
    .Y(_01284_));
 sky130_fd_sc_hd__nor2_1 _21601_ (.A(_05149_),
    .B(_08960_),
    .Y(_01285_));
 sky130_fd_sc_hd__nor2_1 _21602_ (.A(_05157_),
    .B(_08960_),
    .Y(_01286_));
 sky130_fd_sc_hd__nor2_1 _21603_ (.A(_05166_),
    .B(_08960_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_1 _21604_ (.A(_05173_),
    .B(_08960_),
    .Y(_01288_));
 sky130_fd_sc_hd__nor2_1 _21605_ (.A(_05183_),
    .B(_08960_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_8 _21606_ (.A(_09751_),
    .B(_04784_),
    .Y(_08965_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_832 ();
 sky130_fd_sc_hd__nor2_1 _21608_ (.A(_04790_),
    .B(_08965_),
    .Y(_01290_));
 sky130_fd_sc_hd__nor2_1 _21609_ (.A(_04871_),
    .B(_08965_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_1 _21610_ (.A(_04883_),
    .B(_08965_),
    .Y(_01292_));
 sky130_fd_sc_hd__nor2_1 _21611_ (.A(_04892_),
    .B(_08965_),
    .Y(_01293_));
 sky130_fd_sc_hd__nor2_1 _21612_ (.A(_04899_),
    .B(_08965_),
    .Y(_01294_));
 sky130_fd_sc_hd__nor2_1 _21613_ (.A(_04906_),
    .B(_08965_),
    .Y(_01295_));
 sky130_fd_sc_hd__nor2_1 _21614_ (.A(_04913_),
    .B(_08965_),
    .Y(_01296_));
 sky130_fd_sc_hd__nor2_1 _21615_ (.A(_04923_),
    .B(_08965_),
    .Y(_01297_));
 sky130_fd_sc_hd__nor2_1 _21616_ (.A(_04932_),
    .B(_08965_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_1 _21617_ (.A(_04939_),
    .B(_08965_),
    .Y(_01299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_831 ();
 sky130_fd_sc_hd__nor2_1 _21619_ (.A(_04951_),
    .B(_08965_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _21620_ (.A(_04794_),
    .B(_08965_),
    .Y(_01301_));
 sky130_fd_sc_hd__nor2_1 _21621_ (.A(_04960_),
    .B(_08965_),
    .Y(_01302_));
 sky130_fd_sc_hd__nor2_1 _21622_ (.A(_04974_),
    .B(_08965_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_1 _21623_ (.A(_04984_),
    .B(_08965_),
    .Y(_01304_));
 sky130_fd_sc_hd__nor2_1 _21624_ (.A(_04990_),
    .B(_08965_),
    .Y(_01305_));
 sky130_fd_sc_hd__nor2_1 _21625_ (.A(net1139),
    .B(_08965_),
    .Y(_01306_));
 sky130_fd_sc_hd__nor2_1 _21626_ (.A(_05011_),
    .B(_08965_),
    .Y(_01307_));
 sky130_fd_sc_hd__nor2_1 _21627_ (.A(_05020_),
    .B(_08965_),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_1 _21628_ (.A(_05029_),
    .B(_08965_),
    .Y(_01309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_830 ();
 sky130_fd_sc_hd__nor2_1 _21630_ (.A(net1138),
    .B(_08965_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor2_1 _21631_ (.A(net1143),
    .B(_08965_),
    .Y(_01311_));
 sky130_fd_sc_hd__nor2_1 _21632_ (.A(_04801_),
    .B(_08965_),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _21633_ (.A(_05060_),
    .B(_08965_),
    .Y(_01313_));
 sky130_fd_sc_hd__nor2_1 _21634_ (.A(_08895_),
    .B(_08965_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_1 _21635_ (.A(_04808_),
    .B(_08965_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2_1 _21636_ (.A(_04817_),
    .B(_08965_),
    .Y(_01316_));
 sky130_fd_sc_hd__nor2_1 _21637_ (.A(_04826_),
    .B(_08965_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_1 _21638_ (.A(_04834_),
    .B(_08965_),
    .Y(_01318_));
 sky130_fd_sc_hd__nor2_1 _21639_ (.A(_04843_),
    .B(_08965_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_1 _21640_ (.A(_04852_),
    .B(_08965_),
    .Y(_01320_));
 sky130_fd_sc_hd__nor2_1 _21641_ (.A(_04860_),
    .B(_08965_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_8 _21642_ (.A(_09805_),
    .B(_05115_),
    .Y(_08969_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_829 ();
 sky130_fd_sc_hd__nor2_1 _21644_ (.A(_05118_),
    .B(_08969_),
    .Y(_01322_));
 sky130_fd_sc_hd__nor2_1 _21645_ (.A(_05192_),
    .B(_08969_),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2_1 _21646_ (.A(_05204_),
    .B(_08969_),
    .Y(_01324_));
 sky130_fd_sc_hd__nor2_1 _21647_ (.A(_05214_),
    .B(_08969_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_1 _21648_ (.A(_05221_),
    .B(_08969_),
    .Y(_01326_));
 sky130_fd_sc_hd__nor2_1 _21649_ (.A(net1136),
    .B(_08969_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_1 _21650_ (.A(_05238_),
    .B(_08969_),
    .Y(_01328_));
 sky130_fd_sc_hd__nor2_1 _21651_ (.A(net1135),
    .B(_08969_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _21652_ (.A(_05258_),
    .B(_08969_),
    .Y(_01330_));
 sky130_fd_sc_hd__nor2_1 _21653_ (.A(_05267_),
    .B(_08969_),
    .Y(_01331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_828 ();
 sky130_fd_sc_hd__nor2_1 _21655_ (.A(_05280_),
    .B(_08969_),
    .Y(_01332_));
 sky130_fd_sc_hd__nor2_1 _21656_ (.A(_05122_),
    .B(_08969_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2_1 _21657_ (.A(_05291_),
    .B(_08969_),
    .Y(_01334_));
 sky130_fd_sc_hd__nor2_1 _21658_ (.A(_05301_),
    .B(_08969_),
    .Y(_01335_));
 sky130_fd_sc_hd__nor2_1 _21659_ (.A(_05309_),
    .B(_08969_),
    .Y(_01336_));
 sky130_fd_sc_hd__nor2_1 _21660_ (.A(_05320_),
    .B(_08969_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2_1 _21661_ (.A(net1100),
    .B(_08969_),
    .Y(_01338_));
 sky130_fd_sc_hd__nor2_1 _21662_ (.A(_05339_),
    .B(_08969_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2_1 _21663_ (.A(_05347_),
    .B(_08969_),
    .Y(_01340_));
 sky130_fd_sc_hd__nor2_1 _21664_ (.A(net538),
    .B(_08969_),
    .Y(_01341_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_827 ();
 sky130_fd_sc_hd__nor2_1 _21666_ (.A(net1101),
    .B(_08969_),
    .Y(_01342_));
 sky130_fd_sc_hd__nor2_1 _21667_ (.A(_05380_),
    .B(_08969_),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_1 _21668_ (.A(_05126_),
    .B(_08969_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _21669_ (.A(net1129),
    .B(_08969_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _21670_ (.A(net1042),
    .B(_08969_),
    .Y(_01346_));
 sky130_fd_sc_hd__nor2_1 _21671_ (.A(_05132_),
    .B(_08969_),
    .Y(_01347_));
 sky130_fd_sc_hd__nor2_1 _21672_ (.A(_05140_),
    .B(_08969_),
    .Y(_01348_));
 sky130_fd_sc_hd__nor2_1 _21673_ (.A(_05149_),
    .B(_08969_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2_1 _21674_ (.A(_05157_),
    .B(_08969_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor2_1 _21675_ (.A(_05166_),
    .B(_08969_),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2_1 _21676_ (.A(_05173_),
    .B(_08969_),
    .Y(_01352_));
 sky130_fd_sc_hd__nor2_1 _21677_ (.A(_05183_),
    .B(_08969_),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_8 _21678_ (.A(_09751_),
    .B(_05433_),
    .Y(_08973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_826 ();
 sky130_fd_sc_hd__nor2_1 _21680_ (.A(_04790_),
    .B(_08973_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor2_1 _21681_ (.A(_04871_),
    .B(_08973_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2_1 _21682_ (.A(_04883_),
    .B(_08973_),
    .Y(_01356_));
 sky130_fd_sc_hd__nor2_1 _21683_ (.A(_04892_),
    .B(_08973_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_1 _21684_ (.A(_04899_),
    .B(_08973_),
    .Y(_01358_));
 sky130_fd_sc_hd__nor2_1 _21685_ (.A(_04906_),
    .B(_08973_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _21686_ (.A(_04913_),
    .B(_08973_),
    .Y(_01360_));
 sky130_fd_sc_hd__nor2_1 _21687_ (.A(_04923_),
    .B(_08973_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2_1 _21688_ (.A(_04932_),
    .B(_08973_),
    .Y(_01362_));
 sky130_fd_sc_hd__nor2_1 _21689_ (.A(_04939_),
    .B(_08973_),
    .Y(_01363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_825 ();
 sky130_fd_sc_hd__nor2_1 _21691_ (.A(_04951_),
    .B(_08973_),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_1 _21692_ (.A(_04794_),
    .B(_08973_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_1 _21693_ (.A(_04960_),
    .B(_08973_),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_1 _21694_ (.A(_04974_),
    .B(_08973_),
    .Y(_01367_));
 sky130_fd_sc_hd__nor2_1 _21695_ (.A(_04984_),
    .B(_08973_),
    .Y(_01368_));
 sky130_fd_sc_hd__nor2_1 _21696_ (.A(_04990_),
    .B(_08973_),
    .Y(_01369_));
 sky130_fd_sc_hd__nor2_1 _21697_ (.A(net1139),
    .B(_08973_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _21698_ (.A(_05011_),
    .B(_08973_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_1 _21699_ (.A(_05020_),
    .B(_08973_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_1 _21700_ (.A(_05029_),
    .B(_08973_),
    .Y(_01373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_824 ();
 sky130_fd_sc_hd__nor2_1 _21702_ (.A(_05035_),
    .B(_08973_),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_1 _21703_ (.A(_05044_),
    .B(_08973_),
    .Y(_01375_));
 sky130_fd_sc_hd__nor2_1 _21704_ (.A(_04801_),
    .B(_08973_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _21705_ (.A(_05060_),
    .B(_08973_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _21706_ (.A(_08895_),
    .B(_08973_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_1 _21707_ (.A(_04808_),
    .B(_08973_),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_1 _21708_ (.A(_04817_),
    .B(_08973_),
    .Y(_01380_));
 sky130_fd_sc_hd__nor2_1 _21709_ (.A(_04826_),
    .B(_08973_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _21710_ (.A(_04834_),
    .B(_08973_),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_1 _21711_ (.A(_04843_),
    .B(_08973_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _21712_ (.A(_04852_),
    .B(_08973_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_1 _21713_ (.A(_04860_),
    .B(_08973_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_8 _21714_ (.A(_09805_),
    .B(_05474_),
    .Y(_08977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_823 ();
 sky130_fd_sc_hd__nor2_1 _21716_ (.A(_05118_),
    .B(_08977_),
    .Y(_01386_));
 sky130_fd_sc_hd__nor2_1 _21717_ (.A(_05192_),
    .B(_08977_),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_1 _21718_ (.A(_05204_),
    .B(_08977_),
    .Y(_01388_));
 sky130_fd_sc_hd__nor2_1 _21719_ (.A(_05214_),
    .B(_08977_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _21720_ (.A(_05221_),
    .B(_08977_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_1 _21721_ (.A(_05228_),
    .B(_08977_),
    .Y(_01391_));
 sky130_fd_sc_hd__nor2_1 _21722_ (.A(_05238_),
    .B(_08977_),
    .Y(_01392_));
 sky130_fd_sc_hd__nor2_1 _21723_ (.A(net1135),
    .B(_08977_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _21724_ (.A(_05258_),
    .B(_08977_),
    .Y(_01394_));
 sky130_fd_sc_hd__nor2_1 _21725_ (.A(net1102),
    .B(_08977_),
    .Y(_01395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_822 ();
 sky130_fd_sc_hd__nor2_1 _21727_ (.A(_05280_),
    .B(_08977_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _21728_ (.A(_05122_),
    .B(_08977_),
    .Y(_01397_));
 sky130_fd_sc_hd__nor2_1 _21729_ (.A(_05291_),
    .B(_08977_),
    .Y(_01398_));
 sky130_fd_sc_hd__nor2_1 _21730_ (.A(_05301_),
    .B(_08977_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor2_1 _21731_ (.A(_05309_),
    .B(_08977_),
    .Y(_01400_));
 sky130_fd_sc_hd__nor2_1 _21732_ (.A(_05320_),
    .B(_08977_),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(net1137),
    .B(_08977_),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_1 _21734_ (.A(_05339_),
    .B(_08977_),
    .Y(_01403_));
 sky130_fd_sc_hd__nor2_1 _21735_ (.A(_05347_),
    .B(_08977_),
    .Y(_01404_));
 sky130_fd_sc_hd__nor2_1 _21736_ (.A(net538),
    .B(_08977_),
    .Y(_01405_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_821 ();
 sky130_fd_sc_hd__nor2_1 _21738_ (.A(net1142),
    .B(_08977_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _21739_ (.A(_05380_),
    .B(_08977_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _21740_ (.A(_05126_),
    .B(_08977_),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_1 _21741_ (.A(net1134),
    .B(_08977_),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_1 _21742_ (.A(net1042),
    .B(_08977_),
    .Y(_01410_));
 sky130_fd_sc_hd__nor2_1 _21743_ (.A(_05132_),
    .B(_08977_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor2_1 _21744_ (.A(_05140_),
    .B(_08977_),
    .Y(_01412_));
 sky130_fd_sc_hd__nor2_1 _21745_ (.A(_05149_),
    .B(_08977_),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_1 _21746_ (.A(_05157_),
    .B(_08977_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _21747_ (.A(_05166_),
    .B(_08977_),
    .Y(_01415_));
 sky130_fd_sc_hd__nor2_1 _21748_ (.A(_05173_),
    .B(_08977_),
    .Y(_01416_));
 sky130_fd_sc_hd__nor2_1 _21749_ (.A(_05183_),
    .B(_08977_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_8 _21750_ (.A(_09751_),
    .B(_05516_),
    .Y(_08981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_820 ();
 sky130_fd_sc_hd__nor2_1 _21752_ (.A(_04790_),
    .B(_08981_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _21753_ (.A(_04871_),
    .B(_08981_),
    .Y(_01419_));
 sky130_fd_sc_hd__nor2_1 _21754_ (.A(_04883_),
    .B(_08981_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_1 _21755_ (.A(_04892_),
    .B(_08981_),
    .Y(_01421_));
 sky130_fd_sc_hd__nor2_1 _21756_ (.A(_04899_),
    .B(_08981_),
    .Y(_01422_));
 sky130_fd_sc_hd__nor2_1 _21757_ (.A(_04906_),
    .B(_08981_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _21758_ (.A(_04913_),
    .B(_08981_),
    .Y(_01424_));
 sky130_fd_sc_hd__nor2_1 _21759_ (.A(_04923_),
    .B(_08981_),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_1 _21760_ (.A(_04932_),
    .B(_08981_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_1 _21761_ (.A(_04939_),
    .B(_08981_),
    .Y(_01427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_819 ();
 sky130_fd_sc_hd__nor2_1 _21763_ (.A(_04951_),
    .B(_08981_),
    .Y(_01428_));
 sky130_fd_sc_hd__nor2_1 _21764_ (.A(_04794_),
    .B(_08981_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _21765_ (.A(_04960_),
    .B(_08981_),
    .Y(_01430_));
 sky130_fd_sc_hd__nor2_1 _21766_ (.A(_04974_),
    .B(_08981_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_1 _21767_ (.A(_04984_),
    .B(_08981_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_1 _21768_ (.A(_04990_),
    .B(_08981_),
    .Y(_01433_));
 sky130_fd_sc_hd__nor2_1 _21769_ (.A(net1139),
    .B(_08981_),
    .Y(_01434_));
 sky130_fd_sc_hd__nor2_1 _21770_ (.A(_05011_),
    .B(_08981_),
    .Y(_01435_));
 sky130_fd_sc_hd__nor2_1 _21771_ (.A(_05020_),
    .B(_08981_),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_1 _21772_ (.A(_05029_),
    .B(_08981_),
    .Y(_01437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_818 ();
 sky130_fd_sc_hd__nor2_1 _21774_ (.A(_05035_),
    .B(_08981_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _21775_ (.A(net1143),
    .B(_08981_),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_1 _21776_ (.A(_04801_),
    .B(_08981_),
    .Y(_01440_));
 sky130_fd_sc_hd__nor2_1 _21777_ (.A(_05060_),
    .B(_08981_),
    .Y(_01441_));
 sky130_fd_sc_hd__nor2_1 _21778_ (.A(_08895_),
    .B(_08981_),
    .Y(_01442_));
 sky130_fd_sc_hd__nor2_1 _21779_ (.A(_04808_),
    .B(_08981_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2_1 _21780_ (.A(_04817_),
    .B(_08981_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _21781_ (.A(_04826_),
    .B(_08981_),
    .Y(_01445_));
 sky130_fd_sc_hd__nor2_1 _21782_ (.A(_04834_),
    .B(_08981_),
    .Y(_01446_));
 sky130_fd_sc_hd__nor2_1 _21783_ (.A(_04843_),
    .B(_08981_),
    .Y(_01447_));
 sky130_fd_sc_hd__nor2_1 _21784_ (.A(_04852_),
    .B(_08981_),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_1 _21785_ (.A(_04860_),
    .B(_08981_),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_8 _21786_ (.A(_09805_),
    .B(_05557_),
    .Y(_08985_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_817 ();
 sky130_fd_sc_hd__nor2_1 _21788_ (.A(_05118_),
    .B(_08985_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _21789_ (.A(_05192_),
    .B(_08985_),
    .Y(_01451_));
 sky130_fd_sc_hd__nor2_1 _21790_ (.A(_05204_),
    .B(_08985_),
    .Y(_01452_));
 sky130_fd_sc_hd__nor2_1 _21791_ (.A(_05214_),
    .B(_08985_),
    .Y(_01453_));
 sky130_fd_sc_hd__nor2_1 _21792_ (.A(_05221_),
    .B(_08985_),
    .Y(_01454_));
 sky130_fd_sc_hd__nor2_1 _21793_ (.A(_05228_),
    .B(_08985_),
    .Y(_01455_));
 sky130_fd_sc_hd__nor2_1 _21794_ (.A(_05238_),
    .B(_08985_),
    .Y(_01456_));
 sky130_fd_sc_hd__nor2_1 _21795_ (.A(net1135),
    .B(_08985_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor2_1 _21796_ (.A(_05258_),
    .B(_08985_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_1 _21797_ (.A(_05267_),
    .B(_08985_),
    .Y(_01459_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_816 ();
 sky130_fd_sc_hd__nor2_1 _21799_ (.A(_05280_),
    .B(_08985_),
    .Y(_01460_));
 sky130_fd_sc_hd__nor2_1 _21800_ (.A(_05122_),
    .B(_08985_),
    .Y(_01461_));
 sky130_fd_sc_hd__nor2_1 _21801_ (.A(_05291_),
    .B(_08985_),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_1 _21802_ (.A(_05301_),
    .B(_08985_),
    .Y(_01463_));
 sky130_fd_sc_hd__nor2_1 _21803_ (.A(_05309_),
    .B(_08985_),
    .Y(_01464_));
 sky130_fd_sc_hd__nor2_1 _21804_ (.A(_05320_),
    .B(_08985_),
    .Y(_01465_));
 sky130_fd_sc_hd__nor2_1 _21805_ (.A(net1137),
    .B(_08985_),
    .Y(_01466_));
 sky130_fd_sc_hd__nor2_1 _21806_ (.A(_05339_),
    .B(_08985_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _21807_ (.A(_05347_),
    .B(_08985_),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_1 _21808_ (.A(net538),
    .B(_08985_),
    .Y(_01469_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_815 ();
 sky130_fd_sc_hd__nor2_1 _21810_ (.A(net1142),
    .B(_08985_),
    .Y(_01470_));
 sky130_fd_sc_hd__nor2_1 _21811_ (.A(_05380_),
    .B(_08985_),
    .Y(_01471_));
 sky130_fd_sc_hd__nor2_1 _21812_ (.A(_05126_),
    .B(_08985_),
    .Y(_01472_));
 sky130_fd_sc_hd__nor2_1 _21813_ (.A(net1129),
    .B(_08985_),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_1 _21814_ (.A(net1042),
    .B(_08985_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor2_1 _21815_ (.A(_05132_),
    .B(_08985_),
    .Y(_01475_));
 sky130_fd_sc_hd__nor2_1 _21816_ (.A(_05140_),
    .B(_08985_),
    .Y(_01476_));
 sky130_fd_sc_hd__nor2_1 _21817_ (.A(_05149_),
    .B(_08985_),
    .Y(_01477_));
 sky130_fd_sc_hd__nor2_1 _21818_ (.A(_05157_),
    .B(_08985_),
    .Y(_01478_));
 sky130_fd_sc_hd__nor2_1 _21819_ (.A(_05166_),
    .B(_08985_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_1 _21820_ (.A(_05173_),
    .B(_08985_),
    .Y(_01480_));
 sky130_fd_sc_hd__nor2_1 _21821_ (.A(_05183_),
    .B(_08985_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand2_8 _21822_ (.A(_09751_),
    .B(_05598_),
    .Y(_08989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_814 ();
 sky130_fd_sc_hd__nor2_1 _21824_ (.A(_04790_),
    .B(_08989_),
    .Y(_01482_));
 sky130_fd_sc_hd__nor2_1 _21825_ (.A(_04871_),
    .B(_08989_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _21826_ (.A(_04883_),
    .B(_08989_),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_1 _21827_ (.A(_04892_),
    .B(_08989_),
    .Y(_01485_));
 sky130_fd_sc_hd__nor2_1 _21828_ (.A(_04899_),
    .B(_08989_),
    .Y(_01486_));
 sky130_fd_sc_hd__nor2_1 _21829_ (.A(_04906_),
    .B(_08989_),
    .Y(_01487_));
 sky130_fd_sc_hd__nor2_1 _21830_ (.A(_04913_),
    .B(_08989_),
    .Y(_01488_));
 sky130_fd_sc_hd__nor2_1 _21831_ (.A(_04923_),
    .B(_08989_),
    .Y(_01489_));
 sky130_fd_sc_hd__nor2_1 _21832_ (.A(_04932_),
    .B(_08989_),
    .Y(_01490_));
 sky130_fd_sc_hd__nor2_1 _21833_ (.A(_04939_),
    .B(_08989_),
    .Y(_01491_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_813 ();
 sky130_fd_sc_hd__nor2_1 _21835_ (.A(_04951_),
    .B(_08989_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_1 _21836_ (.A(_04794_),
    .B(_08989_),
    .Y(_01493_));
 sky130_fd_sc_hd__nor2_1 _21837_ (.A(_04960_),
    .B(_08989_),
    .Y(_01494_));
 sky130_fd_sc_hd__nor2_1 _21838_ (.A(_04974_),
    .B(_08989_),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_1 _21839_ (.A(_04984_),
    .B(_08989_),
    .Y(_01496_));
 sky130_fd_sc_hd__nor2_1 _21840_ (.A(_04990_),
    .B(_08989_),
    .Y(_01497_));
 sky130_fd_sc_hd__nor2_1 _21841_ (.A(_05000_),
    .B(_08989_),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_1 _21842_ (.A(_05011_),
    .B(_08989_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _21843_ (.A(_05020_),
    .B(_08989_),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_1 _21844_ (.A(_05029_),
    .B(_08989_),
    .Y(_01501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_812 ();
 sky130_fd_sc_hd__nor2_1 _21846_ (.A(_05035_),
    .B(_08989_),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _21847_ (.A(net1143),
    .B(_08989_),
    .Y(_01503_));
 sky130_fd_sc_hd__nor2_1 _21848_ (.A(_04801_),
    .B(_08989_),
    .Y(_01504_));
 sky130_fd_sc_hd__nor2_1 _21849_ (.A(_05060_),
    .B(_08989_),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_1 _21850_ (.A(_08895_),
    .B(_08989_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_1 _21851_ (.A(_04808_),
    .B(_08989_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_1 _21852_ (.A(_04817_),
    .B(_08989_),
    .Y(_01508_));
 sky130_fd_sc_hd__nor2_1 _21853_ (.A(_04826_),
    .B(_08989_),
    .Y(_01509_));
 sky130_fd_sc_hd__nor2_1 _21854_ (.A(_04834_),
    .B(_08989_),
    .Y(_01510_));
 sky130_fd_sc_hd__nor2_1 _21855_ (.A(_04843_),
    .B(_08989_),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_1 _21856_ (.A(_04852_),
    .B(_08989_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_1 _21857_ (.A(_04860_),
    .B(_08989_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_8 _21858_ (.A(_09805_),
    .B(_05951_),
    .Y(_08993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_811 ();
 sky130_fd_sc_hd__nor2_1 _21860_ (.A(_05118_),
    .B(_08993_),
    .Y(_01514_));
 sky130_fd_sc_hd__nor2_1 _21861_ (.A(_05192_),
    .B(_08993_),
    .Y(_01515_));
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(_05204_),
    .B(_08993_),
    .Y(_01516_));
 sky130_fd_sc_hd__nor2_1 _21863_ (.A(_05214_),
    .B(_08993_),
    .Y(_01517_));
 sky130_fd_sc_hd__nor2_1 _21864_ (.A(_05221_),
    .B(_08993_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor2_1 _21865_ (.A(net1136),
    .B(_08993_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor2_1 _21866_ (.A(_05238_),
    .B(_08993_),
    .Y(_01520_));
 sky130_fd_sc_hd__nor2_1 _21867_ (.A(_05247_),
    .B(_08993_),
    .Y(_01521_));
 sky130_fd_sc_hd__nor2_1 _21868_ (.A(_05258_),
    .B(_08993_),
    .Y(_01522_));
 sky130_fd_sc_hd__nor2_1 _21869_ (.A(_05267_),
    .B(_08993_),
    .Y(_01523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_810 ();
 sky130_fd_sc_hd__nor2_1 _21871_ (.A(_05280_),
    .B(_08993_),
    .Y(_01524_));
 sky130_fd_sc_hd__nor2_1 _21872_ (.A(_05122_),
    .B(_08993_),
    .Y(_01525_));
 sky130_fd_sc_hd__nor2_1 _21873_ (.A(_05291_),
    .B(_08993_),
    .Y(_01526_));
 sky130_fd_sc_hd__nor2_1 _21874_ (.A(_05301_),
    .B(_08993_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _21875_ (.A(_05309_),
    .B(_08993_),
    .Y(_01528_));
 sky130_fd_sc_hd__nor2_1 _21876_ (.A(_05320_),
    .B(_08993_),
    .Y(_01529_));
 sky130_fd_sc_hd__nor2_1 _21877_ (.A(net1137),
    .B(_08993_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _21878_ (.A(_05339_),
    .B(_08993_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _21879_ (.A(_05347_),
    .B(_08993_),
    .Y(_01532_));
 sky130_fd_sc_hd__nor2_1 _21880_ (.A(net538),
    .B(_08993_),
    .Y(_01533_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_809 ();
 sky130_fd_sc_hd__nor2_1 _21882_ (.A(net1101),
    .B(_08993_),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _21883_ (.A(_05380_),
    .B(_08993_),
    .Y(_01535_));
 sky130_fd_sc_hd__nor2_1 _21884_ (.A(_05126_),
    .B(_08993_),
    .Y(_01536_));
 sky130_fd_sc_hd__nor2_1 _21885_ (.A(net1129),
    .B(_08993_),
    .Y(_01537_));
 sky130_fd_sc_hd__nor2_1 _21886_ (.A(net1042),
    .B(_08993_),
    .Y(_01538_));
 sky130_fd_sc_hd__nor2_1 _21887_ (.A(_05132_),
    .B(_08993_),
    .Y(_01539_));
 sky130_fd_sc_hd__nor2_1 _21888_ (.A(_05140_),
    .B(_08993_),
    .Y(_01540_));
 sky130_fd_sc_hd__nor2_1 _21889_ (.A(_05149_),
    .B(_08993_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _21890_ (.A(_05157_),
    .B(_08993_),
    .Y(_01542_));
 sky130_fd_sc_hd__nor2_1 _21891_ (.A(_05166_),
    .B(_08993_),
    .Y(_01543_));
 sky130_fd_sc_hd__nor2_1 _21892_ (.A(_05173_),
    .B(_08993_),
    .Y(_01544_));
 sky130_fd_sc_hd__nor2_1 _21893_ (.A(_05183_),
    .B(_08993_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_8 _21894_ (.A(_09759_),
    .B(_04784_),
    .Y(_08997_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_808 ();
 sky130_fd_sc_hd__nor2_1 _21896_ (.A(_04790_),
    .B(_08997_),
    .Y(_01546_));
 sky130_fd_sc_hd__nor2_1 _21897_ (.A(_04871_),
    .B(_08997_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_1 _21898_ (.A(_04883_),
    .B(_08997_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _21899_ (.A(_04892_),
    .B(_08997_),
    .Y(_01549_));
 sky130_fd_sc_hd__nor2_1 _21900_ (.A(_04899_),
    .B(_08997_),
    .Y(_01550_));
 sky130_fd_sc_hd__nor2_1 _21901_ (.A(_04906_),
    .B(_08997_),
    .Y(_01551_));
 sky130_fd_sc_hd__nor2_1 _21902_ (.A(_04913_),
    .B(_08997_),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _21903_ (.A(_04923_),
    .B(_08997_),
    .Y(_01553_));
 sky130_fd_sc_hd__nor2_1 _21904_ (.A(_04932_),
    .B(_08997_),
    .Y(_01554_));
 sky130_fd_sc_hd__nor2_1 _21905_ (.A(_04939_),
    .B(_08997_),
    .Y(_01555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_807 ();
 sky130_fd_sc_hd__nor2_1 _21907_ (.A(_04951_),
    .B(_08997_),
    .Y(_01556_));
 sky130_fd_sc_hd__nor2_1 _21908_ (.A(_04794_),
    .B(_08997_),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2_1 _21909_ (.A(_04960_),
    .B(_08997_),
    .Y(_01558_));
 sky130_fd_sc_hd__nor2_1 _21910_ (.A(_04974_),
    .B(_08997_),
    .Y(_01559_));
 sky130_fd_sc_hd__nor2_1 _21911_ (.A(_04984_),
    .B(_08997_),
    .Y(_01560_));
 sky130_fd_sc_hd__nor2_1 _21912_ (.A(_04990_),
    .B(_08997_),
    .Y(_01561_));
 sky130_fd_sc_hd__nor2_1 _21913_ (.A(net1139),
    .B(_08997_),
    .Y(_01562_));
 sky130_fd_sc_hd__nor2_1 _21914_ (.A(_05011_),
    .B(_08997_),
    .Y(_01563_));
 sky130_fd_sc_hd__nor2_1 _21915_ (.A(_05020_),
    .B(_08997_),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_1 _21916_ (.A(_05029_),
    .B(_08997_),
    .Y(_01565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_806 ();
 sky130_fd_sc_hd__nor2_1 _21918_ (.A(net1138),
    .B(_08997_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_1 _21919_ (.A(net1143),
    .B(_08997_),
    .Y(_01567_));
 sky130_fd_sc_hd__nor2_1 _21920_ (.A(_04801_),
    .B(_08997_),
    .Y(_01568_));
 sky130_fd_sc_hd__nor2_1 _21921_ (.A(_05060_),
    .B(_08997_),
    .Y(_01569_));
 sky130_fd_sc_hd__nor2_1 _21922_ (.A(_08895_),
    .B(_08997_),
    .Y(_01570_));
 sky130_fd_sc_hd__nor2_1 _21923_ (.A(_04808_),
    .B(_08997_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_1 _21924_ (.A(_04817_),
    .B(_08997_),
    .Y(_01572_));
 sky130_fd_sc_hd__nor2_1 _21925_ (.A(_04826_),
    .B(_08997_),
    .Y(_01573_));
 sky130_fd_sc_hd__nor2_1 _21926_ (.A(_04834_),
    .B(_08997_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor2_1 _21927_ (.A(_04843_),
    .B(_08997_),
    .Y(_01575_));
 sky130_fd_sc_hd__nor2_1 _21928_ (.A(_04852_),
    .B(_08997_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _21929_ (.A(_04860_),
    .B(_08997_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand2_8 _21930_ (.A(_09811_),
    .B(_05115_),
    .Y(_09001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_805 ();
 sky130_fd_sc_hd__nor2_1 _21932_ (.A(_05118_),
    .B(_09001_),
    .Y(_01578_));
 sky130_fd_sc_hd__nor2_1 _21933_ (.A(_05192_),
    .B(_09001_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _21934_ (.A(_05204_),
    .B(_09001_),
    .Y(_01580_));
 sky130_fd_sc_hd__nor2_1 _21935_ (.A(_05214_),
    .B(_09001_),
    .Y(_01581_));
 sky130_fd_sc_hd__nor2_1 _21936_ (.A(_05221_),
    .B(_09001_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_1 _21937_ (.A(net1136),
    .B(_09001_),
    .Y(_01583_));
 sky130_fd_sc_hd__nor2_1 _21938_ (.A(_05238_),
    .B(_09001_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _21939_ (.A(_05247_),
    .B(_09001_),
    .Y(_01585_));
 sky130_fd_sc_hd__nor2_1 _21940_ (.A(_05258_),
    .B(_09001_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor2_1 _21941_ (.A(_05267_),
    .B(_09001_),
    .Y(_01587_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_804 ();
 sky130_fd_sc_hd__nor2_1 _21943_ (.A(_05280_),
    .B(_09001_),
    .Y(_01588_));
 sky130_fd_sc_hd__nor2_1 _21944_ (.A(_05122_),
    .B(_09001_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_1 _21945_ (.A(_05291_),
    .B(_09001_),
    .Y(_01590_));
 sky130_fd_sc_hd__nor2_1 _21946_ (.A(_05301_),
    .B(_09001_),
    .Y(_01591_));
 sky130_fd_sc_hd__nor2_1 _21947_ (.A(_05309_),
    .B(_09001_),
    .Y(_01592_));
 sky130_fd_sc_hd__nor2_1 _21948_ (.A(_05320_),
    .B(_09001_),
    .Y(_01593_));
 sky130_fd_sc_hd__nor2_1 _21949_ (.A(net1137),
    .B(_09001_),
    .Y(_01594_));
 sky130_fd_sc_hd__nor2_1 _21950_ (.A(_05339_),
    .B(_09001_),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_1 _21951_ (.A(_05347_),
    .B(_09001_),
    .Y(_01596_));
 sky130_fd_sc_hd__nor2_1 _21952_ (.A(net538),
    .B(_09001_),
    .Y(_01597_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_803 ();
 sky130_fd_sc_hd__nor2_1 _21954_ (.A(net1101),
    .B(_09001_),
    .Y(_01598_));
 sky130_fd_sc_hd__nor2_1 _21955_ (.A(_05380_),
    .B(_09001_),
    .Y(_01599_));
 sky130_fd_sc_hd__nor2_1 _21956_ (.A(_05126_),
    .B(_09001_),
    .Y(_01600_));
 sky130_fd_sc_hd__nor2_1 _21957_ (.A(net1129),
    .B(_09001_),
    .Y(_01601_));
 sky130_fd_sc_hd__nor2_1 _21958_ (.A(_05430_),
    .B(_09001_),
    .Y(_01602_));
 sky130_fd_sc_hd__nor2_1 _21959_ (.A(_05132_),
    .B(_09001_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _21960_ (.A(_05140_),
    .B(_09001_),
    .Y(_01604_));
 sky130_fd_sc_hd__nor2_1 _21961_ (.A(_05149_),
    .B(_09001_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _21962_ (.A(_05157_),
    .B(_09001_),
    .Y(_01606_));
 sky130_fd_sc_hd__nor2_1 _21963_ (.A(_05166_),
    .B(_09001_),
    .Y(_01607_));
 sky130_fd_sc_hd__nor2_1 _21964_ (.A(_05173_),
    .B(_09001_),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_1 _21965_ (.A(_05183_),
    .B(_09001_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_8 _21966_ (.A(_09759_),
    .B(_05433_),
    .Y(_09005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_802 ();
 sky130_fd_sc_hd__nor2_1 _21968_ (.A(_04790_),
    .B(_09005_),
    .Y(_01610_));
 sky130_fd_sc_hd__nor2_1 _21969_ (.A(_04871_),
    .B(_09005_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_1 _21970_ (.A(_04883_),
    .B(_09005_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_1 _21971_ (.A(_04892_),
    .B(_09005_),
    .Y(_01613_));
 sky130_fd_sc_hd__nor2_1 _21972_ (.A(_04899_),
    .B(_09005_),
    .Y(_01614_));
 sky130_fd_sc_hd__nor2_1 _21973_ (.A(_04906_),
    .B(_09005_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_1 _21974_ (.A(_04913_),
    .B(_09005_),
    .Y(_01616_));
 sky130_fd_sc_hd__nor2_1 _21975_ (.A(_04923_),
    .B(_09005_),
    .Y(_01617_));
 sky130_fd_sc_hd__nor2_1 _21976_ (.A(_04932_),
    .B(_09005_),
    .Y(_01618_));
 sky130_fd_sc_hd__nor2_1 _21977_ (.A(_04939_),
    .B(_09005_),
    .Y(_01619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_801 ();
 sky130_fd_sc_hd__nor2_1 _21979_ (.A(_04951_),
    .B(_09005_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _21980_ (.A(_04794_),
    .B(_09005_),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_1 _21981_ (.A(_04960_),
    .B(_09005_),
    .Y(_01622_));
 sky130_fd_sc_hd__nor2_1 _21982_ (.A(_04974_),
    .B(_09005_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_1 _21983_ (.A(_04984_),
    .B(_09005_),
    .Y(_01624_));
 sky130_fd_sc_hd__nor2_1 _21984_ (.A(_04990_),
    .B(_09005_),
    .Y(_01625_));
 sky130_fd_sc_hd__nor2_1 _21985_ (.A(net1139),
    .B(_09005_),
    .Y(_01626_));
 sky130_fd_sc_hd__nor2_1 _21986_ (.A(_05011_),
    .B(_09005_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _21987_ (.A(_05020_),
    .B(_09005_),
    .Y(_01628_));
 sky130_fd_sc_hd__nor2_1 _21988_ (.A(_05029_),
    .B(_09005_),
    .Y(_01629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_800 ();
 sky130_fd_sc_hd__nor2_1 _21990_ (.A(net1138),
    .B(_09005_),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_1 _21991_ (.A(net1143),
    .B(_09005_),
    .Y(_01631_));
 sky130_fd_sc_hd__nor2_1 _21992_ (.A(_04801_),
    .B(_09005_),
    .Y(_01632_));
 sky130_fd_sc_hd__nor2_1 _21993_ (.A(_05060_),
    .B(_09005_),
    .Y(_01633_));
 sky130_fd_sc_hd__nor2_1 _21994_ (.A(_08895_),
    .B(_09005_),
    .Y(_01634_));
 sky130_fd_sc_hd__nor2_1 _21995_ (.A(_04808_),
    .B(_09005_),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_1 _21996_ (.A(_04817_),
    .B(_09005_),
    .Y(_01636_));
 sky130_fd_sc_hd__nor2_1 _21997_ (.A(_04826_),
    .B(_09005_),
    .Y(_01637_));
 sky130_fd_sc_hd__nor2_1 _21998_ (.A(_04834_),
    .B(_09005_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor2_1 _21999_ (.A(_04843_),
    .B(_09005_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_1 _22000_ (.A(_04852_),
    .B(_09005_),
    .Y(_01640_));
 sky130_fd_sc_hd__nor2_1 _22001_ (.A(_04860_),
    .B(_09005_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_8 _22002_ (.A(_09811_),
    .B(_05474_),
    .Y(_09009_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_799 ();
 sky130_fd_sc_hd__nor2_1 _22004_ (.A(_05118_),
    .B(_09009_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor2_1 _22005_ (.A(_05192_),
    .B(_09009_),
    .Y(_01643_));
 sky130_fd_sc_hd__nor2_1 _22006_ (.A(_05204_),
    .B(_09009_),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _22007_ (.A(_05214_),
    .B(_09009_),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_1 _22008_ (.A(_05221_),
    .B(_09009_),
    .Y(_01646_));
 sky130_fd_sc_hd__nor2_1 _22009_ (.A(net1136),
    .B(_09009_),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_1 _22010_ (.A(_05238_),
    .B(_09009_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_1 _22011_ (.A(net1135),
    .B(_09009_),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_1 _22012_ (.A(_05258_),
    .B(_09009_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _22013_ (.A(_05267_),
    .B(_09009_),
    .Y(_01651_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_798 ();
 sky130_fd_sc_hd__nor2_1 _22015_ (.A(_05280_),
    .B(_09009_),
    .Y(_01652_));
 sky130_fd_sc_hd__nor2_1 _22016_ (.A(_05122_),
    .B(_09009_),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _22017_ (.A(_05291_),
    .B(_09009_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_1 _22018_ (.A(_05301_),
    .B(_09009_),
    .Y(_01655_));
 sky130_fd_sc_hd__nor2_1 _22019_ (.A(_05309_),
    .B(_09009_),
    .Y(_01656_));
 sky130_fd_sc_hd__nor2_1 _22020_ (.A(_05320_),
    .B(_09009_),
    .Y(_01657_));
 sky130_fd_sc_hd__nor2_1 _22021_ (.A(net1100),
    .B(_09009_),
    .Y(_01658_));
 sky130_fd_sc_hd__nor2_1 _22022_ (.A(_05339_),
    .B(_09009_),
    .Y(_01659_));
 sky130_fd_sc_hd__nor2_1 _22023_ (.A(_05347_),
    .B(_09009_),
    .Y(_01660_));
 sky130_fd_sc_hd__nor2_1 _22024_ (.A(_05358_),
    .B(_09009_),
    .Y(_01661_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_797 ();
 sky130_fd_sc_hd__nor2_1 _22026_ (.A(net1101),
    .B(_09009_),
    .Y(_01662_));
 sky130_fd_sc_hd__nor2_1 _22027_ (.A(_05380_),
    .B(_09009_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor2_1 _22028_ (.A(_05126_),
    .B(_09009_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_1 _22029_ (.A(net1129),
    .B(_09009_),
    .Y(_01665_));
 sky130_fd_sc_hd__nor2_1 _22030_ (.A(net1042),
    .B(_09009_),
    .Y(_01666_));
 sky130_fd_sc_hd__nor2_1 _22031_ (.A(_05132_),
    .B(_09009_),
    .Y(_01667_));
 sky130_fd_sc_hd__nor2_1 _22032_ (.A(_05140_),
    .B(_09009_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _22033_ (.A(_05149_),
    .B(_09009_),
    .Y(_01669_));
 sky130_fd_sc_hd__nor2_1 _22034_ (.A(_05157_),
    .B(_09009_),
    .Y(_01670_));
 sky130_fd_sc_hd__nor2_1 _22035_ (.A(_05166_),
    .B(_09009_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_1 _22036_ (.A(_05173_),
    .B(_09009_),
    .Y(_01672_));
 sky130_fd_sc_hd__nor2_1 _22037_ (.A(_05183_),
    .B(_09009_),
    .Y(_01673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_796 ();
 sky130_fd_sc_hd__nand2_8 _22039_ (.A(_09759_),
    .B(_05516_),
    .Y(_09014_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_795 ();
 sky130_fd_sc_hd__nor2_1 _22041_ (.A(_04790_),
    .B(_09014_),
    .Y(_01674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_794 ();
 sky130_fd_sc_hd__nor2_1 _22043_ (.A(_04871_),
    .B(_09014_),
    .Y(_01675_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_793 ();
 sky130_fd_sc_hd__nor2_1 _22045_ (.A(_04883_),
    .B(_09014_),
    .Y(_01676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_792 ();
 sky130_fd_sc_hd__nor2_1 _22047_ (.A(_04892_),
    .B(_09014_),
    .Y(_01677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_791 ();
 sky130_fd_sc_hd__nor2_1 _22049_ (.A(_04899_),
    .B(_09014_),
    .Y(_01678_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_790 ();
 sky130_fd_sc_hd__nor2_1 _22051_ (.A(_04906_),
    .B(_09014_),
    .Y(_01679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_789 ();
 sky130_fd_sc_hd__nor2_1 _22053_ (.A(_04913_),
    .B(_09014_),
    .Y(_01680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_788 ();
 sky130_fd_sc_hd__nor2_1 _22055_ (.A(_04923_),
    .B(_09014_),
    .Y(_01681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_787 ();
 sky130_fd_sc_hd__nor2_1 _22057_ (.A(_04932_),
    .B(_09014_),
    .Y(_01682_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_786 ();
 sky130_fd_sc_hd__nor2_1 _22059_ (.A(_04939_),
    .B(_09014_),
    .Y(_01683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_784 ();
 sky130_fd_sc_hd__nor2_1 _22062_ (.A(_04951_),
    .B(_09014_),
    .Y(_01684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_783 ();
 sky130_fd_sc_hd__nor2_1 _22064_ (.A(_04794_),
    .B(_09014_),
    .Y(_01685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_782 ();
 sky130_fd_sc_hd__nor2_1 _22066_ (.A(_04960_),
    .B(_09014_),
    .Y(_01686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_781 ();
 sky130_fd_sc_hd__nor2_1 _22068_ (.A(_04974_),
    .B(_09014_),
    .Y(_01687_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_780 ();
 sky130_fd_sc_hd__nor2_1 _22070_ (.A(_04984_),
    .B(_09014_),
    .Y(_01688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_779 ();
 sky130_fd_sc_hd__nor2_1 _22072_ (.A(_04990_),
    .B(_09014_),
    .Y(_01689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_778 ();
 sky130_fd_sc_hd__nor2_1 _22074_ (.A(_05000_),
    .B(_09014_),
    .Y(_01690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_777 ();
 sky130_fd_sc_hd__nor2_1 _22076_ (.A(_05011_),
    .B(_09014_),
    .Y(_01691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_776 ();
 sky130_fd_sc_hd__nor2_1 _22078_ (.A(_05020_),
    .B(_09014_),
    .Y(_01692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_775 ();
 sky130_fd_sc_hd__nor2_1 _22080_ (.A(_05029_),
    .B(_09014_),
    .Y(_01693_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_773 ();
 sky130_fd_sc_hd__nor2_1 _22083_ (.A(net1138),
    .B(_09014_),
    .Y(_01694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_772 ();
 sky130_fd_sc_hd__nor2_1 _22085_ (.A(net1143),
    .B(_09014_),
    .Y(_01695_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_771 ();
 sky130_fd_sc_hd__nor2_1 _22087_ (.A(_04801_),
    .B(_09014_),
    .Y(_01696_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_770 ();
 sky130_fd_sc_hd__nor2_1 _22089_ (.A(_05060_),
    .B(_09014_),
    .Y(_01697_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_769 ();
 sky130_fd_sc_hd__nor2_1 _22091_ (.A(_08895_),
    .B(_09014_),
    .Y(_01698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_768 ();
 sky130_fd_sc_hd__nor2_1 _22093_ (.A(_04808_),
    .B(_09014_),
    .Y(_01699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_767 ();
 sky130_fd_sc_hd__nor2_1 _22095_ (.A(_04817_),
    .B(_09014_),
    .Y(_01700_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_766 ();
 sky130_fd_sc_hd__nor2_1 _22097_ (.A(_04826_),
    .B(_09014_),
    .Y(_01701_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_765 ();
 sky130_fd_sc_hd__nor2_1 _22099_ (.A(_04834_),
    .B(_09014_),
    .Y(_01702_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_764 ();
 sky130_fd_sc_hd__nor2_1 _22101_ (.A(_04843_),
    .B(_09014_),
    .Y(_01703_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_763 ();
 sky130_fd_sc_hd__nor2_1 _22103_ (.A(_04852_),
    .B(_09014_),
    .Y(_01704_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_762 ();
 sky130_fd_sc_hd__nor2_1 _22105_ (.A(_04860_),
    .B(_09014_),
    .Y(_01705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_761 ();
 sky130_fd_sc_hd__nand2_8 _22107_ (.A(_09811_),
    .B(_05557_),
    .Y(_09050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_760 ();
 sky130_fd_sc_hd__nor2_1 _22109_ (.A(_05118_),
    .B(_09050_),
    .Y(_01706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_759 ();
 sky130_fd_sc_hd__nor2_1 _22111_ (.A(_05192_),
    .B(_09050_),
    .Y(_01707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_758 ();
 sky130_fd_sc_hd__nor2_1 _22113_ (.A(_05204_),
    .B(_09050_),
    .Y(_01708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_757 ();
 sky130_fd_sc_hd__nor2_1 _22115_ (.A(_05214_),
    .B(_09050_),
    .Y(_01709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_756 ();
 sky130_fd_sc_hd__nor2_1 _22117_ (.A(_05221_),
    .B(_09050_),
    .Y(_01710_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_755 ();
 sky130_fd_sc_hd__nor2_1 _22119_ (.A(_05228_),
    .B(_09050_),
    .Y(_01711_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_754 ();
 sky130_fd_sc_hd__nor2_1 _22121_ (.A(_05238_),
    .B(_09050_),
    .Y(_01712_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_753 ();
 sky130_fd_sc_hd__nor2_1 _22123_ (.A(_05247_),
    .B(_09050_),
    .Y(_01713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_752 ();
 sky130_fd_sc_hd__nor2_1 _22125_ (.A(_05258_),
    .B(_09050_),
    .Y(_01714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_751 ();
 sky130_fd_sc_hd__nor2_1 _22127_ (.A(net1102),
    .B(_09050_),
    .Y(_01715_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_749 ();
 sky130_fd_sc_hd__nor2_1 _22130_ (.A(_05280_),
    .B(_09050_),
    .Y(_01716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_748 ();
 sky130_fd_sc_hd__nor2_1 _22132_ (.A(_05122_),
    .B(_09050_),
    .Y(_01717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_747 ();
 sky130_fd_sc_hd__nor2_1 _22134_ (.A(_05291_),
    .B(_09050_),
    .Y(_01718_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_746 ();
 sky130_fd_sc_hd__nor2_1 _22136_ (.A(_05301_),
    .B(_09050_),
    .Y(_01719_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_745 ();
 sky130_fd_sc_hd__nor2_1 _22138_ (.A(_05309_),
    .B(_09050_),
    .Y(_01720_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_744 ();
 sky130_fd_sc_hd__nor2_1 _22140_ (.A(_05320_),
    .B(_09050_),
    .Y(_01721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_743 ();
 sky130_fd_sc_hd__nor2_1 _22142_ (.A(net1137),
    .B(_09050_),
    .Y(_01722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_742 ();
 sky130_fd_sc_hd__nor2_1 _22144_ (.A(_05339_),
    .B(_09050_),
    .Y(_01723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_741 ();
 sky130_fd_sc_hd__nor2_1 _22146_ (.A(_05347_),
    .B(_09050_),
    .Y(_01724_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_740 ();
 sky130_fd_sc_hd__nor2_1 _22148_ (.A(net538),
    .B(_09050_),
    .Y(_01725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_738 ();
 sky130_fd_sc_hd__nor2_1 _22151_ (.A(net1101),
    .B(_09050_),
    .Y(_01726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_737 ();
 sky130_fd_sc_hd__nor2_1 _22153_ (.A(_05380_),
    .B(_09050_),
    .Y(_01727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_736 ();
 sky130_fd_sc_hd__nor2_1 _22155_ (.A(_05126_),
    .B(_09050_),
    .Y(_01728_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_735 ();
 sky130_fd_sc_hd__nor2_1 _22157_ (.A(net1129),
    .B(_09050_),
    .Y(_01729_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_734 ();
 sky130_fd_sc_hd__nor2_1 _22159_ (.A(net1042),
    .B(_09050_),
    .Y(_01730_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_733 ();
 sky130_fd_sc_hd__nor2_1 _22161_ (.A(_05132_),
    .B(_09050_),
    .Y(_01731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_732 ();
 sky130_fd_sc_hd__nor2_1 _22163_ (.A(_05140_),
    .B(_09050_),
    .Y(_01732_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_731 ();
 sky130_fd_sc_hd__nor2_1 _22165_ (.A(_05149_),
    .B(_09050_),
    .Y(_01733_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_730 ();
 sky130_fd_sc_hd__nor2_1 _22167_ (.A(_05157_),
    .B(_09050_),
    .Y(_01734_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_729 ();
 sky130_fd_sc_hd__nor2_1 _22169_ (.A(_05166_),
    .B(_09050_),
    .Y(_01735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_728 ();
 sky130_fd_sc_hd__nor2_1 _22171_ (.A(_05173_),
    .B(_09050_),
    .Y(_01736_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_727 ();
 sky130_fd_sc_hd__nor2_1 _22173_ (.A(_05183_),
    .B(_09050_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_8 _22174_ (.A(_09759_),
    .B(_05598_),
    .Y(_09085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_726 ();
 sky130_fd_sc_hd__nor2_1 _22176_ (.A(_04790_),
    .B(_09085_),
    .Y(_01738_));
 sky130_fd_sc_hd__nor2_1 _22177_ (.A(_04871_),
    .B(_09085_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _22178_ (.A(_04883_),
    .B(_09085_),
    .Y(_01740_));
 sky130_fd_sc_hd__nor2_1 _22179_ (.A(_04892_),
    .B(_09085_),
    .Y(_01741_));
 sky130_fd_sc_hd__nor2_1 _22180_ (.A(_04899_),
    .B(_09085_),
    .Y(_01742_));
 sky130_fd_sc_hd__nor2_1 _22181_ (.A(_04906_),
    .B(_09085_),
    .Y(_01743_));
 sky130_fd_sc_hd__nor2_1 _22182_ (.A(_04913_),
    .B(_09085_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _22183_ (.A(_04923_),
    .B(_09085_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor2_1 _22184_ (.A(_04932_),
    .B(_09085_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _22185_ (.A(_04939_),
    .B(_09085_),
    .Y(_01747_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_725 ();
 sky130_fd_sc_hd__nor2_1 _22187_ (.A(_04951_),
    .B(_09085_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _22188_ (.A(_04794_),
    .B(_09085_),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_1 _22189_ (.A(_04960_),
    .B(_09085_),
    .Y(_01750_));
 sky130_fd_sc_hd__nor2_1 _22190_ (.A(_04974_),
    .B(_09085_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor2_1 _22191_ (.A(_04984_),
    .B(_09085_),
    .Y(_01752_));
 sky130_fd_sc_hd__nor2_1 _22192_ (.A(_04990_),
    .B(_09085_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_1 _22193_ (.A(net1139),
    .B(_09085_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _22194_ (.A(_05011_),
    .B(_09085_),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_1 _22195_ (.A(_05020_),
    .B(_09085_),
    .Y(_01756_));
 sky130_fd_sc_hd__nor2_1 _22196_ (.A(_05029_),
    .B(_09085_),
    .Y(_01757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_724 ();
 sky130_fd_sc_hd__nor2_1 _22198_ (.A(net1138),
    .B(_09085_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _22199_ (.A(net1143),
    .B(_09085_),
    .Y(_01759_));
 sky130_fd_sc_hd__nor2_1 _22200_ (.A(_04801_),
    .B(_09085_),
    .Y(_01760_));
 sky130_fd_sc_hd__nor2_1 _22201_ (.A(_05060_),
    .B(_09085_),
    .Y(_01761_));
 sky130_fd_sc_hd__nor2_1 _22202_ (.A(_08895_),
    .B(_09085_),
    .Y(_01762_));
 sky130_fd_sc_hd__nor2_1 _22203_ (.A(_04808_),
    .B(_09085_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _22204_ (.A(_04817_),
    .B(_09085_),
    .Y(_01764_));
 sky130_fd_sc_hd__nor2_1 _22205_ (.A(_04826_),
    .B(_09085_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_1 _22206_ (.A(_04834_),
    .B(_09085_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor2_1 _22207_ (.A(_04843_),
    .B(_09085_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _22208_ (.A(_04852_),
    .B(_09085_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _22209_ (.A(_04860_),
    .B(_09085_),
    .Y(_01769_));
 sky130_fd_sc_hd__or4_4 _22210_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(net1043),
    .D(_09816_),
    .X(_09089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_722 ();
 sky130_fd_sc_hd__nor2_1 _22213_ (.A(_05118_),
    .B(_09089_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor2_1 _22214_ (.A(_05192_),
    .B(_09089_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _22215_ (.A(_05204_),
    .B(_09089_),
    .Y(_01772_));
 sky130_fd_sc_hd__nor2_1 _22216_ (.A(_05214_),
    .B(_09089_),
    .Y(_01773_));
 sky130_fd_sc_hd__nor2_1 _22217_ (.A(_05221_),
    .B(_09089_),
    .Y(_01774_));
 sky130_fd_sc_hd__nor2_1 _22218_ (.A(net1136),
    .B(_09089_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _22219_ (.A(_05238_),
    .B(_09089_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor2_1 _22220_ (.A(net1135),
    .B(_09089_),
    .Y(_01777_));
 sky130_fd_sc_hd__nor2_1 _22221_ (.A(_05258_),
    .B(_09089_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _22222_ (.A(net1102),
    .B(_09089_),
    .Y(_01779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_721 ();
 sky130_fd_sc_hd__nor2_1 _22224_ (.A(_05280_),
    .B(_09089_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _22225_ (.A(_05122_),
    .B(_09089_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _22226_ (.A(_05291_),
    .B(_09089_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor2_1 _22227_ (.A(_05301_),
    .B(_09089_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_1 _22228_ (.A(_05309_),
    .B(_09089_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _22229_ (.A(_05320_),
    .B(_09089_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _22230_ (.A(net1100),
    .B(_09089_),
    .Y(_01786_));
 sky130_fd_sc_hd__nor2_1 _22231_ (.A(_05339_),
    .B(_09089_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _22232_ (.A(_05347_),
    .B(_09089_),
    .Y(_01788_));
 sky130_fd_sc_hd__nor2_1 _22233_ (.A(_05358_),
    .B(_09089_),
    .Y(_01789_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_720 ();
 sky130_fd_sc_hd__nor2_1 _22235_ (.A(net1101),
    .B(_09089_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor2_1 _22236_ (.A(_05380_),
    .B(_09089_),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _22237_ (.A(_05126_),
    .B(_09089_),
    .Y(_01792_));
 sky130_fd_sc_hd__nor2_1 _22238_ (.A(net1129),
    .B(_09089_),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _22239_ (.A(_05430_),
    .B(_09089_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _22240_ (.A(_05132_),
    .B(_09089_),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_1 _22241_ (.A(_05140_),
    .B(_09089_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _22242_ (.A(_05149_),
    .B(_09089_),
    .Y(_01797_));
 sky130_fd_sc_hd__nor2_1 _22243_ (.A(_05157_),
    .B(_09089_),
    .Y(_01798_));
 sky130_fd_sc_hd__nor2_1 _22244_ (.A(_05166_),
    .B(_09089_),
    .Y(_01799_));
 sky130_fd_sc_hd__nor2_1 _22245_ (.A(_05173_),
    .B(_09089_),
    .Y(_01800_));
 sky130_fd_sc_hd__nor2_1 _22246_ (.A(_05183_),
    .B(_09089_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_8 _22247_ (.A(_09764_),
    .B(_04784_),
    .Y(_09094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_719 ();
 sky130_fd_sc_hd__nor2_1 _22249_ (.A(_04790_),
    .B(_09094_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _22250_ (.A(_04871_),
    .B(_09094_),
    .Y(_01803_));
 sky130_fd_sc_hd__nor2_1 _22251_ (.A(_04883_),
    .B(_09094_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _22252_ (.A(_04892_),
    .B(_09094_),
    .Y(_01805_));
 sky130_fd_sc_hd__nor2_1 _22253_ (.A(_04899_),
    .B(_09094_),
    .Y(_01806_));
 sky130_fd_sc_hd__nor2_1 _22254_ (.A(_04906_),
    .B(_09094_),
    .Y(_01807_));
 sky130_fd_sc_hd__nor2_1 _22255_ (.A(_04913_),
    .B(_09094_),
    .Y(_01808_));
 sky130_fd_sc_hd__nor2_1 _22256_ (.A(_04923_),
    .B(_09094_),
    .Y(_01809_));
 sky130_fd_sc_hd__nor2_1 _22257_ (.A(_04932_),
    .B(_09094_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _22258_ (.A(_04939_),
    .B(_09094_),
    .Y(_01811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_718 ();
 sky130_fd_sc_hd__nor2_1 _22260_ (.A(_04951_),
    .B(_09094_),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_1 _22261_ (.A(_04794_),
    .B(_09094_),
    .Y(_01813_));
 sky130_fd_sc_hd__nor2_1 _22262_ (.A(_04960_),
    .B(_09094_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_1 _22263_ (.A(_04974_),
    .B(_09094_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _22264_ (.A(_04984_),
    .B(_09094_),
    .Y(_01816_));
 sky130_fd_sc_hd__nor2_1 _22265_ (.A(_04990_),
    .B(_09094_),
    .Y(_01817_));
 sky130_fd_sc_hd__nor2_1 _22266_ (.A(net1139),
    .B(_09094_),
    .Y(_01818_));
 sky130_fd_sc_hd__nor2_1 _22267_ (.A(_05011_),
    .B(_09094_),
    .Y(_01819_));
 sky130_fd_sc_hd__nor2_1 _22268_ (.A(_05020_),
    .B(_09094_),
    .Y(_01820_));
 sky130_fd_sc_hd__nor2_1 _22269_ (.A(_05029_),
    .B(_09094_),
    .Y(_01821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_717 ();
 sky130_fd_sc_hd__nor2_1 _22271_ (.A(net1138),
    .B(_09094_),
    .Y(_01822_));
 sky130_fd_sc_hd__nor2_1 _22272_ (.A(net1143),
    .B(_09094_),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_1 _22273_ (.A(_04801_),
    .B(_09094_),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _22274_ (.A(_05060_),
    .B(_09094_),
    .Y(_01825_));
 sky130_fd_sc_hd__nor2_1 _22275_ (.A(_08895_),
    .B(_09094_),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _22276_ (.A(_04808_),
    .B(_09094_),
    .Y(_01827_));
 sky130_fd_sc_hd__nor2_1 _22277_ (.A(_04817_),
    .B(_09094_),
    .Y(_01828_));
 sky130_fd_sc_hd__nor2_1 _22278_ (.A(_04826_),
    .B(_09094_),
    .Y(_01829_));
 sky130_fd_sc_hd__nor2_1 _22279_ (.A(_04834_),
    .B(_09094_),
    .Y(_01830_));
 sky130_fd_sc_hd__nor2_1 _22280_ (.A(_04843_),
    .B(_09094_),
    .Y(_01831_));
 sky130_fd_sc_hd__nor2_1 _22281_ (.A(_04852_),
    .B(_09094_),
    .Y(_01832_));
 sky130_fd_sc_hd__nor2_1 _22282_ (.A(_04860_),
    .B(_09094_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_8 _22283_ (.A(_09818_),
    .B(_05115_),
    .Y(_09098_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_716 ();
 sky130_fd_sc_hd__nor2_1 _22285_ (.A(_05118_),
    .B(_09098_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _22286_ (.A(_05192_),
    .B(_09098_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor2_1 _22287_ (.A(_05204_),
    .B(_09098_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _22288_ (.A(_05214_),
    .B(_09098_),
    .Y(_01837_));
 sky130_fd_sc_hd__nor2_1 _22289_ (.A(_05221_),
    .B(_09098_),
    .Y(_01838_));
 sky130_fd_sc_hd__nor2_1 _22290_ (.A(net1136),
    .B(_09098_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _22291_ (.A(_05238_),
    .B(_09098_),
    .Y(_01840_));
 sky130_fd_sc_hd__nor2_1 _22292_ (.A(net1135),
    .B(_09098_),
    .Y(_01841_));
 sky130_fd_sc_hd__nor2_1 _22293_ (.A(_05258_),
    .B(_09098_),
    .Y(_01842_));
 sky130_fd_sc_hd__nor2_1 _22294_ (.A(net1102),
    .B(_09098_),
    .Y(_01843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_715 ();
 sky130_fd_sc_hd__nor2_1 _22296_ (.A(_05280_),
    .B(_09098_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _22297_ (.A(_05122_),
    .B(_09098_),
    .Y(_01845_));
 sky130_fd_sc_hd__nor2_1 _22298_ (.A(_05291_),
    .B(_09098_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_1 _22299_ (.A(_05301_),
    .B(_09098_),
    .Y(_01847_));
 sky130_fd_sc_hd__nor2_1 _22300_ (.A(_05309_),
    .B(_09098_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_1 _22301_ (.A(_05320_),
    .B(_09098_),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _22302_ (.A(net1100),
    .B(_09098_),
    .Y(_01850_));
 sky130_fd_sc_hd__nor2_1 _22303_ (.A(_05339_),
    .B(_09098_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor2_1 _22304_ (.A(_05347_),
    .B(_09098_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _22305_ (.A(_05358_),
    .B(_09098_),
    .Y(_01853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_714 ();
 sky130_fd_sc_hd__nor2_1 _22307_ (.A(net1142),
    .B(_09098_),
    .Y(_01854_));
 sky130_fd_sc_hd__nor2_1 _22308_ (.A(_05380_),
    .B(_09098_),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_1 _22309_ (.A(_05126_),
    .B(_09098_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _22310_ (.A(net1129),
    .B(_09098_),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _22311_ (.A(net1042),
    .B(_09098_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _22312_ (.A(_05132_),
    .B(_09098_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _22313_ (.A(_05140_),
    .B(_09098_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor2_1 _22314_ (.A(_05149_),
    .B(_09098_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _22315_ (.A(_05157_),
    .B(_09098_),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_1 _22316_ (.A(_05166_),
    .B(_09098_),
    .Y(_01863_));
 sky130_fd_sc_hd__nor2_1 _22317_ (.A(_05173_),
    .B(_09098_),
    .Y(_01864_));
 sky130_fd_sc_hd__nor2_1 _22318_ (.A(_05183_),
    .B(_09098_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_8 _22319_ (.A(_09764_),
    .B(_05433_),
    .Y(_09102_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_713 ();
 sky130_fd_sc_hd__nor2_1 _22321_ (.A(_04790_),
    .B(_09102_),
    .Y(_01866_));
 sky130_fd_sc_hd__nor2_1 _22322_ (.A(_04871_),
    .B(_09102_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor2_1 _22323_ (.A(_04883_),
    .B(_09102_),
    .Y(_01868_));
 sky130_fd_sc_hd__nor2_1 _22324_ (.A(_04892_),
    .B(_09102_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _22325_ (.A(_04899_),
    .B(_09102_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _22326_ (.A(_04906_),
    .B(_09102_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _22327_ (.A(_04913_),
    .B(_09102_),
    .Y(_01872_));
 sky130_fd_sc_hd__nor2_1 _22328_ (.A(_04923_),
    .B(_09102_),
    .Y(_01873_));
 sky130_fd_sc_hd__nor2_1 _22329_ (.A(_04932_),
    .B(_09102_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _22330_ (.A(_04939_),
    .B(_09102_),
    .Y(_01875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_712 ();
 sky130_fd_sc_hd__nor2_1 _22332_ (.A(_04951_),
    .B(_09102_),
    .Y(_01876_));
 sky130_fd_sc_hd__nor2_1 _22333_ (.A(_04794_),
    .B(_09102_),
    .Y(_01877_));
 sky130_fd_sc_hd__nor2_1 _22334_ (.A(_04960_),
    .B(_09102_),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _22335_ (.A(_04974_),
    .B(_09102_),
    .Y(_01879_));
 sky130_fd_sc_hd__nor2_1 _22336_ (.A(_04984_),
    .B(_09102_),
    .Y(_01880_));
 sky130_fd_sc_hd__nor2_1 _22337_ (.A(_04990_),
    .B(_09102_),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_1 _22338_ (.A(_05000_),
    .B(_09102_),
    .Y(_01882_));
 sky130_fd_sc_hd__nor2_1 _22339_ (.A(_05011_),
    .B(_09102_),
    .Y(_01883_));
 sky130_fd_sc_hd__nor2_1 _22340_ (.A(_05020_),
    .B(_09102_),
    .Y(_01884_));
 sky130_fd_sc_hd__nor2_1 _22341_ (.A(_05029_),
    .B(_09102_),
    .Y(_01885_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_711 ();
 sky130_fd_sc_hd__nor2_1 _22343_ (.A(net1138),
    .B(_09102_),
    .Y(_01886_));
 sky130_fd_sc_hd__nor2_1 _22344_ (.A(net1143),
    .B(_09102_),
    .Y(_01887_));
 sky130_fd_sc_hd__nor2_1 _22345_ (.A(_04801_),
    .B(_09102_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor2_1 _22346_ (.A(_05060_),
    .B(_09102_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor2_1 _22347_ (.A(_08895_),
    .B(_09102_),
    .Y(_01890_));
 sky130_fd_sc_hd__nor2_1 _22348_ (.A(_04808_),
    .B(_09102_),
    .Y(_01891_));
 sky130_fd_sc_hd__nor2_1 _22349_ (.A(_04817_),
    .B(_09102_),
    .Y(_01892_));
 sky130_fd_sc_hd__nor2_1 _22350_ (.A(_04826_),
    .B(_09102_),
    .Y(_01893_));
 sky130_fd_sc_hd__nor2_1 _22351_ (.A(_04834_),
    .B(_09102_),
    .Y(_01894_));
 sky130_fd_sc_hd__nor2_1 _22352_ (.A(_04843_),
    .B(_09102_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _22353_ (.A(_04852_),
    .B(_09102_),
    .Y(_01896_));
 sky130_fd_sc_hd__nor2_1 _22354_ (.A(_04860_),
    .B(_09102_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_8 _22355_ (.A(_09818_),
    .B(_05474_),
    .Y(_09106_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_710 ();
 sky130_fd_sc_hd__nor2_1 _22357_ (.A(_05118_),
    .B(_09106_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _22358_ (.A(_05192_),
    .B(_09106_),
    .Y(_01899_));
 sky130_fd_sc_hd__nor2_1 _22359_ (.A(_05204_),
    .B(_09106_),
    .Y(_01900_));
 sky130_fd_sc_hd__nor2_1 _22360_ (.A(_05214_),
    .B(_09106_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _22361_ (.A(_05221_),
    .B(_09106_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _22362_ (.A(_05228_),
    .B(_09106_),
    .Y(_01903_));
 sky130_fd_sc_hd__nor2_1 _22363_ (.A(_05238_),
    .B(_09106_),
    .Y(_01904_));
 sky130_fd_sc_hd__nor2_1 _22364_ (.A(net1135),
    .B(_09106_),
    .Y(_01905_));
 sky130_fd_sc_hd__nor2_1 _22365_ (.A(_05258_),
    .B(_09106_),
    .Y(_01906_));
 sky130_fd_sc_hd__nor2_1 _22366_ (.A(net1102),
    .B(_09106_),
    .Y(_01907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_709 ();
 sky130_fd_sc_hd__nor2_1 _22368_ (.A(_05280_),
    .B(_09106_),
    .Y(_01908_));
 sky130_fd_sc_hd__nor2_1 _22369_ (.A(_05122_),
    .B(_09106_),
    .Y(_01909_));
 sky130_fd_sc_hd__nor2_1 _22370_ (.A(_05291_),
    .B(_09106_),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _22371_ (.A(_05301_),
    .B(_09106_),
    .Y(_01911_));
 sky130_fd_sc_hd__nor2_1 _22372_ (.A(_05309_),
    .B(_09106_),
    .Y(_01912_));
 sky130_fd_sc_hd__nor2_1 _22373_ (.A(_05320_),
    .B(_09106_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _22374_ (.A(net1100),
    .B(_09106_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _22375_ (.A(_05339_),
    .B(_09106_),
    .Y(_01915_));
 sky130_fd_sc_hd__nor2_1 _22376_ (.A(_05347_),
    .B(_09106_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _22377_ (.A(_05358_),
    .B(_09106_),
    .Y(_01917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_708 ();
 sky130_fd_sc_hd__nor2_1 _22379_ (.A(net1101),
    .B(_09106_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _22380_ (.A(_05380_),
    .B(_09106_),
    .Y(_01919_));
 sky130_fd_sc_hd__nor2_1 _22381_ (.A(_05126_),
    .B(_09106_),
    .Y(_01920_));
 sky130_fd_sc_hd__nor2_1 _22382_ (.A(net1129),
    .B(_09106_),
    .Y(_01921_));
 sky130_fd_sc_hd__nor2_1 _22383_ (.A(net1042),
    .B(_09106_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _22384_ (.A(_05132_),
    .B(_09106_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_1 _22385_ (.A(_05140_),
    .B(_09106_),
    .Y(_01924_));
 sky130_fd_sc_hd__nor2_1 _22386_ (.A(_05149_),
    .B(_09106_),
    .Y(_01925_));
 sky130_fd_sc_hd__nor2_1 _22387_ (.A(_05157_),
    .B(_09106_),
    .Y(_01926_));
 sky130_fd_sc_hd__nor2_1 _22388_ (.A(_05166_),
    .B(_09106_),
    .Y(_01927_));
 sky130_fd_sc_hd__nor2_1 _22389_ (.A(_05173_),
    .B(_09106_),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _22390_ (.A(_05183_),
    .B(_09106_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_8 _22391_ (.A(_09764_),
    .B(_05516_),
    .Y(_09110_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_707 ();
 sky130_fd_sc_hd__nor2_1 _22393_ (.A(_04790_),
    .B(_09110_),
    .Y(_01930_));
 sky130_fd_sc_hd__nor2_1 _22394_ (.A(_04871_),
    .B(_09110_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _22395_ (.A(_04883_),
    .B(_09110_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_1 _22396_ (.A(_04892_),
    .B(_09110_),
    .Y(_01933_));
 sky130_fd_sc_hd__nor2_1 _22397_ (.A(_04899_),
    .B(_09110_),
    .Y(_01934_));
 sky130_fd_sc_hd__nor2_1 _22398_ (.A(_04906_),
    .B(_09110_),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_1 _22399_ (.A(_04913_),
    .B(_09110_),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _22400_ (.A(_04923_),
    .B(_09110_),
    .Y(_01937_));
 sky130_fd_sc_hd__nor2_1 _22401_ (.A(_04932_),
    .B(_09110_),
    .Y(_01938_));
 sky130_fd_sc_hd__nor2_1 _22402_ (.A(_04939_),
    .B(_09110_),
    .Y(_01939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_706 ();
 sky130_fd_sc_hd__nor2_1 _22404_ (.A(_04951_),
    .B(_09110_),
    .Y(_01940_));
 sky130_fd_sc_hd__nor2_1 _22405_ (.A(_04794_),
    .B(_09110_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor2_1 _22406_ (.A(_04960_),
    .B(_09110_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_1 _22407_ (.A(_04974_),
    .B(_09110_),
    .Y(_01943_));
 sky130_fd_sc_hd__nor2_1 _22408_ (.A(_04984_),
    .B(_09110_),
    .Y(_01944_));
 sky130_fd_sc_hd__nor2_1 _22409_ (.A(_04990_),
    .B(_09110_),
    .Y(_01945_));
 sky130_fd_sc_hd__nor2_1 _22410_ (.A(net1139),
    .B(_09110_),
    .Y(_01946_));
 sky130_fd_sc_hd__nor2_1 _22411_ (.A(_05011_),
    .B(_09110_),
    .Y(_01947_));
 sky130_fd_sc_hd__nor2_1 _22412_ (.A(_05020_),
    .B(_09110_),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_1 _22413_ (.A(_05029_),
    .B(_09110_),
    .Y(_01949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_705 ();
 sky130_fd_sc_hd__nor2_1 _22415_ (.A(net1138),
    .B(_09110_),
    .Y(_01950_));
 sky130_fd_sc_hd__nor2_1 _22416_ (.A(_05044_),
    .B(_09110_),
    .Y(_01951_));
 sky130_fd_sc_hd__nor2_1 _22417_ (.A(_04801_),
    .B(_09110_),
    .Y(_01952_));
 sky130_fd_sc_hd__nor2_1 _22418_ (.A(_05060_),
    .B(_09110_),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _22419_ (.A(_08895_),
    .B(_09110_),
    .Y(_01954_));
 sky130_fd_sc_hd__nor2_1 _22420_ (.A(_04808_),
    .B(_09110_),
    .Y(_01955_));
 sky130_fd_sc_hd__nor2_1 _22421_ (.A(_04817_),
    .B(_09110_),
    .Y(_01956_));
 sky130_fd_sc_hd__nor2_1 _22422_ (.A(_04826_),
    .B(_09110_),
    .Y(_01957_));
 sky130_fd_sc_hd__nor2_1 _22423_ (.A(_04834_),
    .B(_09110_),
    .Y(_01958_));
 sky130_fd_sc_hd__nor2_1 _22424_ (.A(_04843_),
    .B(_09110_),
    .Y(_01959_));
 sky130_fd_sc_hd__nor2_1 _22425_ (.A(_04852_),
    .B(_09110_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2_1 _22426_ (.A(_04860_),
    .B(_09110_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_8 _22427_ (.A(_09818_),
    .B(_05557_),
    .Y(_09114_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_704 ();
 sky130_fd_sc_hd__nor2_1 _22429_ (.A(_05118_),
    .B(_09114_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _22430_ (.A(_05192_),
    .B(_09114_),
    .Y(_01963_));
 sky130_fd_sc_hd__nor2_1 _22431_ (.A(_05204_),
    .B(_09114_),
    .Y(_01964_));
 sky130_fd_sc_hd__nor2_1 _22432_ (.A(_05214_),
    .B(_09114_),
    .Y(_01965_));
 sky130_fd_sc_hd__nor2_1 _22433_ (.A(_05221_),
    .B(_09114_),
    .Y(_01966_));
 sky130_fd_sc_hd__nor2_1 _22434_ (.A(net1136),
    .B(_09114_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _22435_ (.A(_05238_),
    .B(_09114_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor2_1 _22436_ (.A(net1135),
    .B(_09114_),
    .Y(_01969_));
 sky130_fd_sc_hd__nor2_1 _22437_ (.A(_05258_),
    .B(_09114_),
    .Y(_01970_));
 sky130_fd_sc_hd__nor2_1 _22438_ (.A(net1102),
    .B(_09114_),
    .Y(_01971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_703 ();
 sky130_fd_sc_hd__nor2_1 _22440_ (.A(_05280_),
    .B(_09114_),
    .Y(_01972_));
 sky130_fd_sc_hd__nor2_1 _22441_ (.A(_05122_),
    .B(_09114_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_1 _22442_ (.A(_05291_),
    .B(_09114_),
    .Y(_01974_));
 sky130_fd_sc_hd__nor2_1 _22443_ (.A(_05301_),
    .B(_09114_),
    .Y(_01975_));
 sky130_fd_sc_hd__nor2_1 _22444_ (.A(_05309_),
    .B(_09114_),
    .Y(_01976_));
 sky130_fd_sc_hd__nor2_1 _22445_ (.A(_05320_),
    .B(_09114_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_1 _22446_ (.A(net1100),
    .B(_09114_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _22447_ (.A(_05339_),
    .B(_09114_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _22448_ (.A(_05347_),
    .B(_09114_),
    .Y(_01980_));
 sky130_fd_sc_hd__nor2_1 _22449_ (.A(_05358_),
    .B(_09114_),
    .Y(_01981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_702 ();
 sky130_fd_sc_hd__nor2_1 _22451_ (.A(net1142),
    .B(_09114_),
    .Y(_01982_));
 sky130_fd_sc_hd__nor2_1 _22452_ (.A(_05380_),
    .B(_09114_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _22453_ (.A(_05126_),
    .B(_09114_),
    .Y(_01984_));
 sky130_fd_sc_hd__nor2_1 _22454_ (.A(net1129),
    .B(_09114_),
    .Y(_01985_));
 sky130_fd_sc_hd__nor2_1 _22455_ (.A(net1042),
    .B(_09114_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_1 _22456_ (.A(_05132_),
    .B(_09114_),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2_1 _22457_ (.A(_05140_),
    .B(_09114_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor2_1 _22458_ (.A(_05149_),
    .B(_09114_),
    .Y(_01989_));
 sky130_fd_sc_hd__nor2_1 _22459_ (.A(_05157_),
    .B(_09114_),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_1 _22460_ (.A(_05166_),
    .B(_09114_),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_1 _22461_ (.A(_05173_),
    .B(_09114_),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _22462_ (.A(_05183_),
    .B(_09114_),
    .Y(_01993_));
 sky130_fd_sc_hd__nand2_8 _22463_ (.A(_09764_),
    .B(_05598_),
    .Y(_09118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_701 ();
 sky130_fd_sc_hd__nor2_1 _22465_ (.A(_04790_),
    .B(_09118_),
    .Y(_01994_));
 sky130_fd_sc_hd__nor2_1 _22466_ (.A(_04871_),
    .B(_09118_),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_1 _22467_ (.A(_04883_),
    .B(_09118_),
    .Y(_01996_));
 sky130_fd_sc_hd__nor2_1 _22468_ (.A(_04892_),
    .B(_09118_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _22469_ (.A(_04899_),
    .B(_09118_),
    .Y(_01998_));
 sky130_fd_sc_hd__nor2_1 _22470_ (.A(_04906_),
    .B(_09118_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor2_1 _22471_ (.A(_04913_),
    .B(_09118_),
    .Y(_02000_));
 sky130_fd_sc_hd__nor2_1 _22472_ (.A(_04923_),
    .B(_09118_),
    .Y(_02001_));
 sky130_fd_sc_hd__nor2_1 _22473_ (.A(_04932_),
    .B(_09118_),
    .Y(_02002_));
 sky130_fd_sc_hd__nor2_1 _22474_ (.A(_04939_),
    .B(_09118_),
    .Y(_02003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_700 ();
 sky130_fd_sc_hd__nor2_1 _22476_ (.A(_04951_),
    .B(_09118_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_1 _22477_ (.A(_04794_),
    .B(_09118_),
    .Y(_02005_));
 sky130_fd_sc_hd__nor2_1 _22478_ (.A(_04960_),
    .B(_09118_),
    .Y(_02006_));
 sky130_fd_sc_hd__nor2_1 _22479_ (.A(_04974_),
    .B(_09118_),
    .Y(_02007_));
 sky130_fd_sc_hd__nor2_1 _22480_ (.A(_04984_),
    .B(_09118_),
    .Y(_02008_));
 sky130_fd_sc_hd__nor2_1 _22481_ (.A(_04990_),
    .B(_09118_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _22482_ (.A(_05000_),
    .B(_09118_),
    .Y(_02010_));
 sky130_fd_sc_hd__nor2_1 _22483_ (.A(_05011_),
    .B(_09118_),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _22484_ (.A(_05020_),
    .B(_09118_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_1 _22485_ (.A(_05029_),
    .B(_09118_),
    .Y(_02013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_699 ();
 sky130_fd_sc_hd__nor2_1 _22487_ (.A(net1138),
    .B(_09118_),
    .Y(_02014_));
 sky130_fd_sc_hd__nor2_1 _22488_ (.A(_05044_),
    .B(_09118_),
    .Y(_02015_));
 sky130_fd_sc_hd__nor2_1 _22489_ (.A(_04801_),
    .B(_09118_),
    .Y(_02016_));
 sky130_fd_sc_hd__nor2_1 _22490_ (.A(_05060_),
    .B(_09118_),
    .Y(_02017_));
 sky130_fd_sc_hd__nor2_1 _22491_ (.A(_08895_),
    .B(_09118_),
    .Y(_02018_));
 sky130_fd_sc_hd__nor2_1 _22492_ (.A(_04808_),
    .B(_09118_),
    .Y(_02019_));
 sky130_fd_sc_hd__nor2_1 _22493_ (.A(_04817_),
    .B(_09118_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _22494_ (.A(_04826_),
    .B(_09118_),
    .Y(_02021_));
 sky130_fd_sc_hd__nor2_1 _22495_ (.A(_04834_),
    .B(_09118_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_1 _22496_ (.A(_04843_),
    .B(_09118_),
    .Y(_02023_));
 sky130_fd_sc_hd__nor2_1 _22497_ (.A(_04852_),
    .B(_09118_),
    .Y(_02024_));
 sky130_fd_sc_hd__nor2_1 _22498_ (.A(_04860_),
    .B(_09118_),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_8 _22499_ (.A(_09818_),
    .B(_05951_),
    .Y(_09122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_698 ();
 sky130_fd_sc_hd__nor2_1 _22501_ (.A(_05118_),
    .B(_09122_),
    .Y(_02026_));
 sky130_fd_sc_hd__nor2_1 _22502_ (.A(_05192_),
    .B(_09122_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _22503_ (.A(_05204_),
    .B(_09122_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _22504_ (.A(_05214_),
    .B(_09122_),
    .Y(_02029_));
 sky130_fd_sc_hd__nor2_1 _22505_ (.A(_05221_),
    .B(_09122_),
    .Y(_02030_));
 sky130_fd_sc_hd__nor2_1 _22506_ (.A(net1136),
    .B(_09122_),
    .Y(_02031_));
 sky130_fd_sc_hd__nor2_1 _22507_ (.A(_05238_),
    .B(_09122_),
    .Y(_02032_));
 sky130_fd_sc_hd__nor2_1 _22508_ (.A(net1135),
    .B(_09122_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_1 _22509_ (.A(_05258_),
    .B(_09122_),
    .Y(_02034_));
 sky130_fd_sc_hd__nor2_1 _22510_ (.A(net1102),
    .B(_09122_),
    .Y(_02035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_697 ();
 sky130_fd_sc_hd__nor2_1 _22512_ (.A(_05280_),
    .B(_09122_),
    .Y(_02036_));
 sky130_fd_sc_hd__nor2_1 _22513_ (.A(_05122_),
    .B(_09122_),
    .Y(_02037_));
 sky130_fd_sc_hd__nor2_1 _22514_ (.A(_05291_),
    .B(_09122_),
    .Y(_02038_));
 sky130_fd_sc_hd__nor2_1 _22515_ (.A(_05301_),
    .B(_09122_),
    .Y(_02039_));
 sky130_fd_sc_hd__nor2_1 _22516_ (.A(_05309_),
    .B(_09122_),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _22517_ (.A(_05320_),
    .B(_09122_),
    .Y(_02041_));
 sky130_fd_sc_hd__nor2_1 _22518_ (.A(net1100),
    .B(_09122_),
    .Y(_02042_));
 sky130_fd_sc_hd__nor2_1 _22519_ (.A(_05339_),
    .B(_09122_),
    .Y(_02043_));
 sky130_fd_sc_hd__nor2_1 _22520_ (.A(_05347_),
    .B(_09122_),
    .Y(_02044_));
 sky130_fd_sc_hd__nor2_1 _22521_ (.A(_05358_),
    .B(_09122_),
    .Y(_02045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_696 ();
 sky130_fd_sc_hd__nor2_1 _22523_ (.A(net1101),
    .B(_09122_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_1 _22524_ (.A(_05380_),
    .B(_09122_),
    .Y(_02047_));
 sky130_fd_sc_hd__nor2_1 _22525_ (.A(_05126_),
    .B(_09122_),
    .Y(_02048_));
 sky130_fd_sc_hd__nor2_1 _22526_ (.A(net1134),
    .B(_09122_),
    .Y(_02049_));
 sky130_fd_sc_hd__nor2_1 _22527_ (.A(net1042),
    .B(_09122_),
    .Y(_02050_));
 sky130_fd_sc_hd__nor2_1 _22528_ (.A(_05132_),
    .B(_09122_),
    .Y(_02051_));
 sky130_fd_sc_hd__nor2_1 _22529_ (.A(_05140_),
    .B(_09122_),
    .Y(_02052_));
 sky130_fd_sc_hd__nor2_1 _22530_ (.A(_05149_),
    .B(_09122_),
    .Y(_02053_));
 sky130_fd_sc_hd__nor2_1 _22531_ (.A(_05157_),
    .B(_09122_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _22532_ (.A(_05166_),
    .B(_09122_),
    .Y(_02055_));
 sky130_fd_sc_hd__nor2_1 _22533_ (.A(_05173_),
    .B(_09122_),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_1 _22534_ (.A(_05183_),
    .B(_09122_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_8 _22535_ (.A(_09771_),
    .B(_04784_),
    .Y(_09126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_695 ();
 sky130_fd_sc_hd__nor2_1 _22537_ (.A(_04790_),
    .B(_09126_),
    .Y(_02058_));
 sky130_fd_sc_hd__nor2_1 _22538_ (.A(_04871_),
    .B(_09126_),
    .Y(_02059_));
 sky130_fd_sc_hd__nor2_1 _22539_ (.A(_04883_),
    .B(_09126_),
    .Y(_02060_));
 sky130_fd_sc_hd__nor2_1 _22540_ (.A(_04892_),
    .B(_09126_),
    .Y(_02061_));
 sky130_fd_sc_hd__nor2_1 _22541_ (.A(_04899_),
    .B(_09126_),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _22542_ (.A(_04906_),
    .B(_09126_),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_1 _22543_ (.A(_04913_),
    .B(_09126_),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _22544_ (.A(_04923_),
    .B(_09126_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor2_1 _22545_ (.A(_04932_),
    .B(_09126_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _22546_ (.A(_04939_),
    .B(_09126_),
    .Y(_02067_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_694 ();
 sky130_fd_sc_hd__nor2_1 _22548_ (.A(_04951_),
    .B(_09126_),
    .Y(_02068_));
 sky130_fd_sc_hd__nor2_1 _22549_ (.A(_04794_),
    .B(_09126_),
    .Y(_02069_));
 sky130_fd_sc_hd__nor2_1 _22550_ (.A(_04960_),
    .B(_09126_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_1 _22551_ (.A(_04974_),
    .B(_09126_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_1 _22552_ (.A(_04984_),
    .B(_09126_),
    .Y(_02072_));
 sky130_fd_sc_hd__nor2_1 _22553_ (.A(_04990_),
    .B(_09126_),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_1 _22554_ (.A(_05000_),
    .B(_09126_),
    .Y(_02074_));
 sky130_fd_sc_hd__nor2_1 _22555_ (.A(_05011_),
    .B(_09126_),
    .Y(_02075_));
 sky130_fd_sc_hd__nor2_1 _22556_ (.A(_05020_),
    .B(_09126_),
    .Y(_02076_));
 sky130_fd_sc_hd__nor2_1 _22557_ (.A(_05029_),
    .B(_09126_),
    .Y(_02077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_693 ();
 sky130_fd_sc_hd__nor2_1 _22559_ (.A(_05035_),
    .B(_09126_),
    .Y(_02078_));
 sky130_fd_sc_hd__nor2_1 _22560_ (.A(_05044_),
    .B(_09126_),
    .Y(_02079_));
 sky130_fd_sc_hd__nor2_1 _22561_ (.A(_04801_),
    .B(_09126_),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _22562_ (.A(_05060_),
    .B(_09126_),
    .Y(_02081_));
 sky130_fd_sc_hd__nor2_1 _22563_ (.A(_08895_),
    .B(_09126_),
    .Y(_02082_));
 sky130_fd_sc_hd__nor2_1 _22564_ (.A(_04808_),
    .B(_09126_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_1 _22565_ (.A(_04817_),
    .B(_09126_),
    .Y(_02084_));
 sky130_fd_sc_hd__nor2_1 _22566_ (.A(_04826_),
    .B(_09126_),
    .Y(_02085_));
 sky130_fd_sc_hd__nor2_1 _22567_ (.A(_04834_),
    .B(_09126_),
    .Y(_02086_));
 sky130_fd_sc_hd__nor2_1 _22568_ (.A(_04843_),
    .B(_09126_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor2_1 _22569_ (.A(_04852_),
    .B(_09126_),
    .Y(_02088_));
 sky130_fd_sc_hd__nor2_1 _22570_ (.A(_04860_),
    .B(_09126_),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_8 _22571_ (.A(_09825_),
    .B(_05115_),
    .Y(_09130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_692 ();
 sky130_fd_sc_hd__nor2_1 _22573_ (.A(_05118_),
    .B(_09130_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _22574_ (.A(_05192_),
    .B(_09130_),
    .Y(_02091_));
 sky130_fd_sc_hd__nor2_1 _22575_ (.A(_05204_),
    .B(_09130_),
    .Y(_02092_));
 sky130_fd_sc_hd__nor2_1 _22576_ (.A(_05214_),
    .B(_09130_),
    .Y(_02093_));
 sky130_fd_sc_hd__nor2_1 _22577_ (.A(_05221_),
    .B(_09130_),
    .Y(_02094_));
 sky130_fd_sc_hd__nor2_1 _22578_ (.A(_05228_),
    .B(_09130_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor2_1 _22579_ (.A(_05238_),
    .B(_09130_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_1 _22580_ (.A(_05247_),
    .B(_09130_),
    .Y(_02097_));
 sky130_fd_sc_hd__nor2_1 _22581_ (.A(_05258_),
    .B(_09130_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_1 _22582_ (.A(net1102),
    .B(_09130_),
    .Y(_02099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_691 ();
 sky130_fd_sc_hd__nor2_1 _22584_ (.A(_05280_),
    .B(_09130_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_1 _22585_ (.A(_05122_),
    .B(_09130_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor2_1 _22586_ (.A(_05291_),
    .B(_09130_),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _22587_ (.A(_05301_),
    .B(_09130_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _22588_ (.A(_05309_),
    .B(_09130_),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _22589_ (.A(_05320_),
    .B(_09130_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _22590_ (.A(net1100),
    .B(_09130_),
    .Y(_02106_));
 sky130_fd_sc_hd__nor2_1 _22591_ (.A(_05339_),
    .B(_09130_),
    .Y(_02107_));
 sky130_fd_sc_hd__nor2_1 _22592_ (.A(_05347_),
    .B(_09130_),
    .Y(_02108_));
 sky130_fd_sc_hd__nor2_1 _22593_ (.A(_05358_),
    .B(_09130_),
    .Y(_02109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_690 ();
 sky130_fd_sc_hd__nor2_1 _22595_ (.A(net1101),
    .B(_09130_),
    .Y(_02110_));
 sky130_fd_sc_hd__nor2_1 _22596_ (.A(_05380_),
    .B(_09130_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor2_1 _22597_ (.A(_05126_),
    .B(_09130_),
    .Y(_02112_));
 sky130_fd_sc_hd__nor2_1 _22598_ (.A(net1134),
    .B(_09130_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor2_1 _22599_ (.A(net1042),
    .B(_09130_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _22600_ (.A(_05132_),
    .B(_09130_),
    .Y(_02115_));
 sky130_fd_sc_hd__nor2_1 _22601_ (.A(_05140_),
    .B(_09130_),
    .Y(_02116_));
 sky130_fd_sc_hd__nor2_1 _22602_ (.A(_05149_),
    .B(_09130_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _22603_ (.A(_05157_),
    .B(_09130_),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_1 _22604_ (.A(_05166_),
    .B(_09130_),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _22605_ (.A(_05173_),
    .B(_09130_),
    .Y(_02120_));
 sky130_fd_sc_hd__nor2_1 _22606_ (.A(_05183_),
    .B(_09130_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_8 _22607_ (.A(_09771_),
    .B(_05433_),
    .Y(_09134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_689 ();
 sky130_fd_sc_hd__nor2_1 _22609_ (.A(_04790_),
    .B(_09134_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _22610_ (.A(_04871_),
    .B(_09134_),
    .Y(_02123_));
 sky130_fd_sc_hd__nor2_1 _22611_ (.A(_04883_),
    .B(_09134_),
    .Y(_02124_));
 sky130_fd_sc_hd__nor2_1 _22612_ (.A(_04892_),
    .B(_09134_),
    .Y(_02125_));
 sky130_fd_sc_hd__nor2_1 _22613_ (.A(_04899_),
    .B(_09134_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor2_1 _22614_ (.A(_04906_),
    .B(_09134_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _22615_ (.A(_04913_),
    .B(_09134_),
    .Y(_02128_));
 sky130_fd_sc_hd__nor2_1 _22616_ (.A(_04923_),
    .B(_09134_),
    .Y(_02129_));
 sky130_fd_sc_hd__nor2_1 _22617_ (.A(_04932_),
    .B(_09134_),
    .Y(_02130_));
 sky130_fd_sc_hd__nor2_1 _22618_ (.A(_04939_),
    .B(_09134_),
    .Y(_02131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_688 ();
 sky130_fd_sc_hd__nor2_1 _22620_ (.A(_04951_),
    .B(_09134_),
    .Y(_02132_));
 sky130_fd_sc_hd__nor2_1 _22621_ (.A(_04794_),
    .B(_09134_),
    .Y(_02133_));
 sky130_fd_sc_hd__nor2_1 _22622_ (.A(_04960_),
    .B(_09134_),
    .Y(_02134_));
 sky130_fd_sc_hd__nor2_1 _22623_ (.A(_04974_),
    .B(_09134_),
    .Y(_02135_));
 sky130_fd_sc_hd__nor2_1 _22624_ (.A(_04984_),
    .B(_09134_),
    .Y(_02136_));
 sky130_fd_sc_hd__nor2_1 _22625_ (.A(_04990_),
    .B(_09134_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _22626_ (.A(net1139),
    .B(_09134_),
    .Y(_02138_));
 sky130_fd_sc_hd__nor2_1 _22627_ (.A(_05011_),
    .B(_09134_),
    .Y(_02139_));
 sky130_fd_sc_hd__nor2_1 _22628_ (.A(_05020_),
    .B(_09134_),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2_1 _22629_ (.A(_05029_),
    .B(_09134_),
    .Y(_02141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_687 ();
 sky130_fd_sc_hd__nor2_1 _22631_ (.A(net1138),
    .B(_09134_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _22632_ (.A(net1143),
    .B(_09134_),
    .Y(_02143_));
 sky130_fd_sc_hd__nor2_1 _22633_ (.A(_04801_),
    .B(_09134_),
    .Y(_02144_));
 sky130_fd_sc_hd__nor2_1 _22634_ (.A(_05060_),
    .B(_09134_),
    .Y(_02145_));
 sky130_fd_sc_hd__nor2_1 _22635_ (.A(_08895_),
    .B(_09134_),
    .Y(_02146_));
 sky130_fd_sc_hd__nor2_1 _22636_ (.A(_04808_),
    .B(_09134_),
    .Y(_02147_));
 sky130_fd_sc_hd__nor2_1 _22637_ (.A(_04817_),
    .B(_09134_),
    .Y(_02148_));
 sky130_fd_sc_hd__nor2_1 _22638_ (.A(_04826_),
    .B(_09134_),
    .Y(_02149_));
 sky130_fd_sc_hd__nor2_1 _22639_ (.A(_04834_),
    .B(_09134_),
    .Y(_02150_));
 sky130_fd_sc_hd__nor2_1 _22640_ (.A(_04843_),
    .B(_09134_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_1 _22641_ (.A(_04852_),
    .B(_09134_),
    .Y(_02152_));
 sky130_fd_sc_hd__nor2_1 _22642_ (.A(_04860_),
    .B(_09134_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_8 _22643_ (.A(_09825_),
    .B(_05474_),
    .Y(_09138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_686 ();
 sky130_fd_sc_hd__nor2_1 _22645_ (.A(_05118_),
    .B(_09138_),
    .Y(_02154_));
 sky130_fd_sc_hd__nor2_1 _22646_ (.A(_05192_),
    .B(_09138_),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _22647_ (.A(_05204_),
    .B(_09138_),
    .Y(_02156_));
 sky130_fd_sc_hd__nor2_1 _22648_ (.A(_05214_),
    .B(_09138_),
    .Y(_02157_));
 sky130_fd_sc_hd__nor2_1 _22649_ (.A(_05221_),
    .B(_09138_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _22650_ (.A(_05228_),
    .B(_09138_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _22651_ (.A(_05238_),
    .B(_09138_),
    .Y(_02160_));
 sky130_fd_sc_hd__nor2_1 _22652_ (.A(net1135),
    .B(_09138_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_1 _22653_ (.A(_05258_),
    .B(_09138_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _22654_ (.A(net1102),
    .B(_09138_),
    .Y(_02163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_685 ();
 sky130_fd_sc_hd__nor2_1 _22656_ (.A(_05280_),
    .B(_09138_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _22657_ (.A(_05122_),
    .B(_09138_),
    .Y(_02165_));
 sky130_fd_sc_hd__nor2_1 _22658_ (.A(_05291_),
    .B(_09138_),
    .Y(_02166_));
 sky130_fd_sc_hd__nor2_1 _22659_ (.A(_05301_),
    .B(_09138_),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _22660_ (.A(_05309_),
    .B(_09138_),
    .Y(_02168_));
 sky130_fd_sc_hd__nor2_1 _22661_ (.A(_05320_),
    .B(_09138_),
    .Y(_02169_));
 sky130_fd_sc_hd__nor2_1 _22662_ (.A(net1100),
    .B(_09138_),
    .Y(_02170_));
 sky130_fd_sc_hd__nor2_1 _22663_ (.A(_05339_),
    .B(_09138_),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_1 _22664_ (.A(_05347_),
    .B(_09138_),
    .Y(_02172_));
 sky130_fd_sc_hd__nor2_1 _22665_ (.A(_05358_),
    .B(_09138_),
    .Y(_02173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_684 ();
 sky130_fd_sc_hd__nor2_1 _22667_ (.A(net1101),
    .B(_09138_),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_1 _22668_ (.A(_05380_),
    .B(_09138_),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _22669_ (.A(_05126_),
    .B(_09138_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _22670_ (.A(net1134),
    .B(_09138_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _22671_ (.A(net1042),
    .B(_09138_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _22672_ (.A(_05132_),
    .B(_09138_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_1 _22673_ (.A(_05140_),
    .B(_09138_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _22674_ (.A(_05149_),
    .B(_09138_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_1 _22675_ (.A(_05157_),
    .B(_09138_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_1 _22676_ (.A(_05166_),
    .B(_09138_),
    .Y(_02183_));
 sky130_fd_sc_hd__nor2_1 _22677_ (.A(_05173_),
    .B(_09138_),
    .Y(_02184_));
 sky130_fd_sc_hd__nor2_1 _22678_ (.A(_05183_),
    .B(_09138_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand2_8 _22679_ (.A(_09771_),
    .B(_05516_),
    .Y(_09142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_683 ();
 sky130_fd_sc_hd__nor2_1 _22681_ (.A(_04790_),
    .B(_09142_),
    .Y(_02186_));
 sky130_fd_sc_hd__nor2_1 _22682_ (.A(_04871_),
    .B(_09142_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _22683_ (.A(_04883_),
    .B(_09142_),
    .Y(_02188_));
 sky130_fd_sc_hd__nor2_1 _22684_ (.A(_04892_),
    .B(_09142_),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _22685_ (.A(_04899_),
    .B(_09142_),
    .Y(_02190_));
 sky130_fd_sc_hd__nor2_1 _22686_ (.A(_04906_),
    .B(_09142_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _22687_ (.A(_04913_),
    .B(_09142_),
    .Y(_02192_));
 sky130_fd_sc_hd__nor2_1 _22688_ (.A(_04923_),
    .B(_09142_),
    .Y(_02193_));
 sky130_fd_sc_hd__nor2_1 _22689_ (.A(_04932_),
    .B(_09142_),
    .Y(_02194_));
 sky130_fd_sc_hd__nor2_1 _22690_ (.A(_04939_),
    .B(_09142_),
    .Y(_02195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_682 ();
 sky130_fd_sc_hd__nor2_1 _22692_ (.A(_04951_),
    .B(_09142_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _22693_ (.A(_04794_),
    .B(_09142_),
    .Y(_02197_));
 sky130_fd_sc_hd__nor2_1 _22694_ (.A(_04960_),
    .B(_09142_),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _22695_ (.A(_04974_),
    .B(_09142_),
    .Y(_02199_));
 sky130_fd_sc_hd__nor2_1 _22696_ (.A(_04984_),
    .B(_09142_),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_1 _22697_ (.A(_04990_),
    .B(_09142_),
    .Y(_02201_));
 sky130_fd_sc_hd__nor2_1 _22698_ (.A(net1139),
    .B(_09142_),
    .Y(_02202_));
 sky130_fd_sc_hd__nor2_1 _22699_ (.A(_05011_),
    .B(_09142_),
    .Y(_02203_));
 sky130_fd_sc_hd__nor2_1 _22700_ (.A(_05020_),
    .B(_09142_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _22701_ (.A(_05029_),
    .B(_09142_),
    .Y(_02205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_681 ();
 sky130_fd_sc_hd__nor2_1 _22703_ (.A(_05035_),
    .B(_09142_),
    .Y(_02206_));
 sky130_fd_sc_hd__nor2_1 _22704_ (.A(net1143),
    .B(_09142_),
    .Y(_02207_));
 sky130_fd_sc_hd__nor2_1 _22705_ (.A(_04801_),
    .B(_09142_),
    .Y(_02208_));
 sky130_fd_sc_hd__nor2_1 _22706_ (.A(_05060_),
    .B(_09142_),
    .Y(_02209_));
 sky130_fd_sc_hd__nor2_1 _22707_ (.A(_08895_),
    .B(_09142_),
    .Y(_02210_));
 sky130_fd_sc_hd__nor2_1 _22708_ (.A(_04808_),
    .B(_09142_),
    .Y(_02211_));
 sky130_fd_sc_hd__nor2_1 _22709_ (.A(_04817_),
    .B(_09142_),
    .Y(_02212_));
 sky130_fd_sc_hd__nor2_1 _22710_ (.A(_04826_),
    .B(_09142_),
    .Y(_02213_));
 sky130_fd_sc_hd__nor2_1 _22711_ (.A(_04834_),
    .B(_09142_),
    .Y(_02214_));
 sky130_fd_sc_hd__nor2_1 _22712_ (.A(_04843_),
    .B(_09142_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _22713_ (.A(_04852_),
    .B(_09142_),
    .Y(_02216_));
 sky130_fd_sc_hd__nor2_1 _22714_ (.A(_04860_),
    .B(_09142_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_8 _22715_ (.A(_09825_),
    .B(_05557_),
    .Y(_09146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_680 ();
 sky130_fd_sc_hd__nor2_1 _22717_ (.A(_05118_),
    .B(_09146_),
    .Y(_02218_));
 sky130_fd_sc_hd__nor2_1 _22718_ (.A(_05192_),
    .B(_09146_),
    .Y(_02219_));
 sky130_fd_sc_hd__nor2_1 _22719_ (.A(_05204_),
    .B(_09146_),
    .Y(_02220_));
 sky130_fd_sc_hd__nor2_1 _22720_ (.A(_05214_),
    .B(_09146_),
    .Y(_02221_));
 sky130_fd_sc_hd__nor2_1 _22721_ (.A(_05221_),
    .B(_09146_),
    .Y(_02222_));
 sky130_fd_sc_hd__nor2_1 _22722_ (.A(net1136),
    .B(_09146_),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _22723_ (.A(_05238_),
    .B(_09146_),
    .Y(_02224_));
 sky130_fd_sc_hd__nor2_1 _22724_ (.A(net1135),
    .B(_09146_),
    .Y(_02225_));
 sky130_fd_sc_hd__nor2_1 _22725_ (.A(_05258_),
    .B(_09146_),
    .Y(_02226_));
 sky130_fd_sc_hd__nor2_1 _22726_ (.A(net1102),
    .B(_09146_),
    .Y(_02227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_679 ();
 sky130_fd_sc_hd__nor2_1 _22728_ (.A(_05280_),
    .B(_09146_),
    .Y(_02228_));
 sky130_fd_sc_hd__nor2_1 _22729_ (.A(_05122_),
    .B(_09146_),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _22730_ (.A(_05291_),
    .B(_09146_),
    .Y(_02230_));
 sky130_fd_sc_hd__nor2_1 _22731_ (.A(_05301_),
    .B(_09146_),
    .Y(_02231_));
 sky130_fd_sc_hd__nor2_1 _22732_ (.A(_05309_),
    .B(_09146_),
    .Y(_02232_));
 sky130_fd_sc_hd__nor2_1 _22733_ (.A(_05320_),
    .B(_09146_),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_1 _22734_ (.A(net1100),
    .B(_09146_),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _22735_ (.A(_05339_),
    .B(_09146_),
    .Y(_02235_));
 sky130_fd_sc_hd__nor2_1 _22736_ (.A(_05347_),
    .B(_09146_),
    .Y(_02236_));
 sky130_fd_sc_hd__nor2_1 _22737_ (.A(_05358_),
    .B(_09146_),
    .Y(_02237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_678 ();
 sky130_fd_sc_hd__nor2_1 _22739_ (.A(net1101),
    .B(_09146_),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_1 _22740_ (.A(_05380_),
    .B(_09146_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _22741_ (.A(_05126_),
    .B(_09146_),
    .Y(_02240_));
 sky130_fd_sc_hd__nor2_1 _22742_ (.A(net1129),
    .B(_09146_),
    .Y(_02241_));
 sky130_fd_sc_hd__nor2_1 _22743_ (.A(net1042),
    .B(_09146_),
    .Y(_02242_));
 sky130_fd_sc_hd__nor2_1 _22744_ (.A(_05132_),
    .B(_09146_),
    .Y(_02243_));
 sky130_fd_sc_hd__nor2_1 _22745_ (.A(_05140_),
    .B(_09146_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_1 _22746_ (.A(_05149_),
    .B(_09146_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _22747_ (.A(_05157_),
    .B(_09146_),
    .Y(_02246_));
 sky130_fd_sc_hd__nor2_1 _22748_ (.A(_05166_),
    .B(_09146_),
    .Y(_02247_));
 sky130_fd_sc_hd__nor2_1 _22749_ (.A(_05173_),
    .B(_09146_),
    .Y(_02248_));
 sky130_fd_sc_hd__nor2_1 _22750_ (.A(_05183_),
    .B(_09146_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_8 _22751_ (.A(_09771_),
    .B(_05598_),
    .Y(_09150_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_677 ();
 sky130_fd_sc_hd__nor2_1 _22753_ (.A(_04790_),
    .B(_09150_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _22754_ (.A(_04871_),
    .B(_09150_),
    .Y(_02251_));
 sky130_fd_sc_hd__nor2_1 _22755_ (.A(_04883_),
    .B(_09150_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor2_1 _22756_ (.A(_04892_),
    .B(_09150_),
    .Y(_02253_));
 sky130_fd_sc_hd__nor2_1 _22757_ (.A(_04899_),
    .B(_09150_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor2_1 _22758_ (.A(_04906_),
    .B(_09150_),
    .Y(_02255_));
 sky130_fd_sc_hd__nor2_1 _22759_ (.A(_04913_),
    .B(_09150_),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_1 _22760_ (.A(_04923_),
    .B(_09150_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _22761_ (.A(_04932_),
    .B(_09150_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _22762_ (.A(_04939_),
    .B(_09150_),
    .Y(_02259_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_676 ();
 sky130_fd_sc_hd__nor2_1 _22764_ (.A(_04951_),
    .B(_09150_),
    .Y(_02260_));
 sky130_fd_sc_hd__nor2_1 _22765_ (.A(_04794_),
    .B(_09150_),
    .Y(_02261_));
 sky130_fd_sc_hd__nor2_1 _22766_ (.A(_04960_),
    .B(_09150_),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_1 _22767_ (.A(_04974_),
    .B(_09150_),
    .Y(_02263_));
 sky130_fd_sc_hd__nor2_1 _22768_ (.A(_04984_),
    .B(_09150_),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _22769_ (.A(_04990_),
    .B(_09150_),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _22770_ (.A(net1139),
    .B(_09150_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_1 _22771_ (.A(_05011_),
    .B(_09150_),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _22772_ (.A(_05020_),
    .B(_09150_),
    .Y(_02268_));
 sky130_fd_sc_hd__nor2_1 _22773_ (.A(_05029_),
    .B(_09150_),
    .Y(_02269_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_675 ();
 sky130_fd_sc_hd__nor2_1 _22775_ (.A(net1138),
    .B(_09150_),
    .Y(_02270_));
 sky130_fd_sc_hd__nor2_1 _22776_ (.A(net1143),
    .B(_09150_),
    .Y(_02271_));
 sky130_fd_sc_hd__nor2_1 _22777_ (.A(_04801_),
    .B(_09150_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _22778_ (.A(_05060_),
    .B(_09150_),
    .Y(_02273_));
 sky130_fd_sc_hd__nor2_1 _22779_ (.A(_08895_),
    .B(_09150_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _22780_ (.A(_04808_),
    .B(_09150_),
    .Y(_02275_));
 sky130_fd_sc_hd__nor2_1 _22781_ (.A(_04817_),
    .B(_09150_),
    .Y(_02276_));
 sky130_fd_sc_hd__nor2_1 _22782_ (.A(_04826_),
    .B(_09150_),
    .Y(_02277_));
 sky130_fd_sc_hd__nor2_1 _22783_ (.A(_04834_),
    .B(_09150_),
    .Y(_02278_));
 sky130_fd_sc_hd__nor2_1 _22784_ (.A(_04843_),
    .B(_09150_),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_1 _22785_ (.A(_04852_),
    .B(_09150_),
    .Y(_02280_));
 sky130_fd_sc_hd__nor2_1 _22786_ (.A(_04860_),
    .B(_09150_),
    .Y(_02281_));
 sky130_fd_sc_hd__or3_4 _22787_ (.A(net1043),
    .B(_09816_),
    .C(_09793_),
    .X(_09154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_673 ();
 sky130_fd_sc_hd__nor2_1 _22790_ (.A(_05118_),
    .B(_09154_),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2_1 _22791_ (.A(_05192_),
    .B(_09154_),
    .Y(_02283_));
 sky130_fd_sc_hd__nor2_1 _22792_ (.A(_05204_),
    .B(_09154_),
    .Y(_02284_));
 sky130_fd_sc_hd__nor2_1 _22793_ (.A(_05214_),
    .B(_09154_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _22794_ (.A(_05221_),
    .B(_09154_),
    .Y(_02286_));
 sky130_fd_sc_hd__nor2_1 _22795_ (.A(net1136),
    .B(_09154_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_1 _22796_ (.A(_05238_),
    .B(_09154_),
    .Y(_02288_));
 sky130_fd_sc_hd__nor2_1 _22797_ (.A(_05247_),
    .B(_09154_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _22798_ (.A(_05258_),
    .B(_09154_),
    .Y(_02290_));
 sky130_fd_sc_hd__nor2_1 _22799_ (.A(net1102),
    .B(_09154_),
    .Y(_02291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_672 ();
 sky130_fd_sc_hd__nor2_1 _22801_ (.A(_05280_),
    .B(_09154_),
    .Y(_02292_));
 sky130_fd_sc_hd__nor2_1 _22802_ (.A(_05122_),
    .B(_09154_),
    .Y(_02293_));
 sky130_fd_sc_hd__nor2_1 _22803_ (.A(_05291_),
    .B(_09154_),
    .Y(_02294_));
 sky130_fd_sc_hd__nor2_1 _22804_ (.A(_05301_),
    .B(_09154_),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_1 _22805_ (.A(_05309_),
    .B(_09154_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor2_1 _22806_ (.A(_05320_),
    .B(_09154_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _22807_ (.A(net1100),
    .B(_09154_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _22808_ (.A(_05339_),
    .B(_09154_),
    .Y(_02299_));
 sky130_fd_sc_hd__nor2_1 _22809_ (.A(_05347_),
    .B(_09154_),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _22810_ (.A(_05358_),
    .B(_09154_),
    .Y(_02301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_671 ();
 sky130_fd_sc_hd__nor2_1 _22812_ (.A(net1101),
    .B(_09154_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _22813_ (.A(_05380_),
    .B(_09154_),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _22814_ (.A(_05126_),
    .B(_09154_),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _22815_ (.A(net1134),
    .B(_09154_),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _22816_ (.A(net1042),
    .B(_09154_),
    .Y(_02306_));
 sky130_fd_sc_hd__nor2_1 _22817_ (.A(_05132_),
    .B(_09154_),
    .Y(_02307_));
 sky130_fd_sc_hd__nor2_1 _22818_ (.A(_05140_),
    .B(_09154_),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2_1 _22819_ (.A(_05149_),
    .B(_09154_),
    .Y(_02309_));
 sky130_fd_sc_hd__nor2_1 _22820_ (.A(_05157_),
    .B(_09154_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor2_1 _22821_ (.A(_05166_),
    .B(_09154_),
    .Y(_02311_));
 sky130_fd_sc_hd__nor2_1 _22822_ (.A(_05173_),
    .B(_09154_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _22823_ (.A(_05183_),
    .B(_09154_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_8 _22824_ (.A(_09778_),
    .B(_04784_),
    .Y(_09159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_670 ();
 sky130_fd_sc_hd__nor2_1 _22826_ (.A(_04790_),
    .B(_09159_),
    .Y(_02314_));
 sky130_fd_sc_hd__nor2_1 _22827_ (.A(_04871_),
    .B(_09159_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _22828_ (.A(_04883_),
    .B(_09159_),
    .Y(_02316_));
 sky130_fd_sc_hd__nor2_1 _22829_ (.A(_04892_),
    .B(_09159_),
    .Y(_02317_));
 sky130_fd_sc_hd__nor2_1 _22830_ (.A(_04899_),
    .B(_09159_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_1 _22831_ (.A(_04906_),
    .B(_09159_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _22832_ (.A(_04913_),
    .B(_09159_),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _22833_ (.A(_04923_),
    .B(_09159_),
    .Y(_02321_));
 sky130_fd_sc_hd__nor2_1 _22834_ (.A(_04932_),
    .B(_09159_),
    .Y(_02322_));
 sky130_fd_sc_hd__nor2_1 _22835_ (.A(_04939_),
    .B(_09159_),
    .Y(_02323_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_669 ();
 sky130_fd_sc_hd__nor2_1 _22837_ (.A(_04951_),
    .B(_09159_),
    .Y(_02324_));
 sky130_fd_sc_hd__nor2_1 _22838_ (.A(_04794_),
    .B(_09159_),
    .Y(_02325_));
 sky130_fd_sc_hd__nor2_1 _22839_ (.A(_04960_),
    .B(_09159_),
    .Y(_02326_));
 sky130_fd_sc_hd__nor2_1 _22840_ (.A(_04974_),
    .B(_09159_),
    .Y(_02327_));
 sky130_fd_sc_hd__nor2_1 _22841_ (.A(_04984_),
    .B(_09159_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_1 _22842_ (.A(_04990_),
    .B(_09159_),
    .Y(_02329_));
 sky130_fd_sc_hd__nor2_1 _22843_ (.A(net1139),
    .B(_09159_),
    .Y(_02330_));
 sky130_fd_sc_hd__nor2_1 _22844_ (.A(_05011_),
    .B(_09159_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_1 _22845_ (.A(_05020_),
    .B(_09159_),
    .Y(_02332_));
 sky130_fd_sc_hd__nor2_1 _22846_ (.A(_05029_),
    .B(_09159_),
    .Y(_02333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_668 ();
 sky130_fd_sc_hd__nor2_1 _22848_ (.A(_05035_),
    .B(_09159_),
    .Y(_02334_));
 sky130_fd_sc_hd__nor2_1 _22849_ (.A(net1143),
    .B(_09159_),
    .Y(_02335_));
 sky130_fd_sc_hd__nor2_1 _22850_ (.A(_04801_),
    .B(_09159_),
    .Y(_02336_));
 sky130_fd_sc_hd__nor2_1 _22851_ (.A(_05060_),
    .B(_09159_),
    .Y(_02337_));
 sky130_fd_sc_hd__nor2_1 _22852_ (.A(_08895_),
    .B(_09159_),
    .Y(_02338_));
 sky130_fd_sc_hd__nor2_1 _22853_ (.A(_04808_),
    .B(_09159_),
    .Y(_02339_));
 sky130_fd_sc_hd__nor2_1 _22854_ (.A(_04817_),
    .B(_09159_),
    .Y(_02340_));
 sky130_fd_sc_hd__nor2_1 _22855_ (.A(_04826_),
    .B(_09159_),
    .Y(_02341_));
 sky130_fd_sc_hd__nor2_1 _22856_ (.A(_04834_),
    .B(_09159_),
    .Y(_02342_));
 sky130_fd_sc_hd__nor2_1 _22857_ (.A(_04843_),
    .B(_09159_),
    .Y(_02343_));
 sky130_fd_sc_hd__nor2_1 _22858_ (.A(_04852_),
    .B(_09159_),
    .Y(_02344_));
 sky130_fd_sc_hd__nor2_1 _22859_ (.A(_04860_),
    .B(_09159_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand2_8 _22860_ (.A(_09830_),
    .B(_05115_),
    .Y(_09163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_667 ();
 sky130_fd_sc_hd__nor2_1 _22862_ (.A(_05118_),
    .B(_09163_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _22863_ (.A(_05192_),
    .B(_09163_),
    .Y(_02347_));
 sky130_fd_sc_hd__nor2_1 _22864_ (.A(_05204_),
    .B(_09163_),
    .Y(_02348_));
 sky130_fd_sc_hd__nor2_1 _22865_ (.A(_05214_),
    .B(_09163_),
    .Y(_02349_));
 sky130_fd_sc_hd__nor2_1 _22866_ (.A(_05221_),
    .B(_09163_),
    .Y(_02350_));
 sky130_fd_sc_hd__nor2_1 _22867_ (.A(net1136),
    .B(_09163_),
    .Y(_02351_));
 sky130_fd_sc_hd__nor2_1 _22868_ (.A(_05238_),
    .B(_09163_),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_1 _22869_ (.A(_05247_),
    .B(_09163_),
    .Y(_02353_));
 sky130_fd_sc_hd__nor2_1 _22870_ (.A(_05258_),
    .B(_09163_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _22871_ (.A(net1102),
    .B(_09163_),
    .Y(_02355_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_666 ();
 sky130_fd_sc_hd__nor2_1 _22873_ (.A(_05280_),
    .B(_09163_),
    .Y(_02356_));
 sky130_fd_sc_hd__nor2_1 _22874_ (.A(_05122_),
    .B(_09163_),
    .Y(_02357_));
 sky130_fd_sc_hd__nor2_1 _22875_ (.A(_05291_),
    .B(_09163_),
    .Y(_02358_));
 sky130_fd_sc_hd__nor2_1 _22876_ (.A(_05301_),
    .B(_09163_),
    .Y(_02359_));
 sky130_fd_sc_hd__nor2_1 _22877_ (.A(_05309_),
    .B(_09163_),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_1 _22878_ (.A(_05320_),
    .B(_09163_),
    .Y(_02361_));
 sky130_fd_sc_hd__nor2_1 _22879_ (.A(net1100),
    .B(_09163_),
    .Y(_02362_));
 sky130_fd_sc_hd__nor2_1 _22880_ (.A(_05339_),
    .B(_09163_),
    .Y(_02363_));
 sky130_fd_sc_hd__nor2_1 _22881_ (.A(_05347_),
    .B(_09163_),
    .Y(_02364_));
 sky130_fd_sc_hd__nor2_1 _22882_ (.A(_05358_),
    .B(_09163_),
    .Y(_02365_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_665 ();
 sky130_fd_sc_hd__nor2_1 _22884_ (.A(net1101),
    .B(_09163_),
    .Y(_02366_));
 sky130_fd_sc_hd__nor2_1 _22885_ (.A(_05380_),
    .B(_09163_),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_1 _22886_ (.A(_05126_),
    .B(_09163_),
    .Y(_02368_));
 sky130_fd_sc_hd__nor2_1 _22887_ (.A(net1134),
    .B(_09163_),
    .Y(_02369_));
 sky130_fd_sc_hd__nor2_1 _22888_ (.A(net1042),
    .B(_09163_),
    .Y(_02370_));
 sky130_fd_sc_hd__nor2_1 _22889_ (.A(_05132_),
    .B(_09163_),
    .Y(_02371_));
 sky130_fd_sc_hd__nor2_1 _22890_ (.A(_05140_),
    .B(_09163_),
    .Y(_02372_));
 sky130_fd_sc_hd__nor2_1 _22891_ (.A(_05149_),
    .B(_09163_),
    .Y(_02373_));
 sky130_fd_sc_hd__nor2_1 _22892_ (.A(_05157_),
    .B(_09163_),
    .Y(_02374_));
 sky130_fd_sc_hd__nor2_1 _22893_ (.A(_05166_),
    .B(_09163_),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2_1 _22894_ (.A(_05173_),
    .B(_09163_),
    .Y(_02376_));
 sky130_fd_sc_hd__nor2_1 _22895_ (.A(_05183_),
    .B(_09163_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_8 _22896_ (.A(_09778_),
    .B(_05433_),
    .Y(_09167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_664 ();
 sky130_fd_sc_hd__nor2_1 _22898_ (.A(_04790_),
    .B(_09167_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _22899_ (.A(_04871_),
    .B(_09167_),
    .Y(_02379_));
 sky130_fd_sc_hd__nor2_1 _22900_ (.A(_04883_),
    .B(_09167_),
    .Y(_02380_));
 sky130_fd_sc_hd__nor2_1 _22901_ (.A(_04892_),
    .B(_09167_),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_1 _22902_ (.A(_04899_),
    .B(_09167_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor2_1 _22903_ (.A(_04906_),
    .B(_09167_),
    .Y(_02383_));
 sky130_fd_sc_hd__nor2_1 _22904_ (.A(_04913_),
    .B(_09167_),
    .Y(_02384_));
 sky130_fd_sc_hd__nor2_1 _22905_ (.A(_04923_),
    .B(_09167_),
    .Y(_02385_));
 sky130_fd_sc_hd__nor2_1 _22906_ (.A(_04932_),
    .B(_09167_),
    .Y(_02386_));
 sky130_fd_sc_hd__nor2_1 _22907_ (.A(_04939_),
    .B(_09167_),
    .Y(_02387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_663 ();
 sky130_fd_sc_hd__nor2_1 _22909_ (.A(_04951_),
    .B(_09167_),
    .Y(_02388_));
 sky130_fd_sc_hd__nor2_1 _22910_ (.A(_04794_),
    .B(_09167_),
    .Y(_02389_));
 sky130_fd_sc_hd__nor2_1 _22911_ (.A(_04960_),
    .B(_09167_),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_1 _22912_ (.A(_04974_),
    .B(_09167_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_1 _22913_ (.A(_04984_),
    .B(_09167_),
    .Y(_02392_));
 sky130_fd_sc_hd__nor2_1 _22914_ (.A(_04990_),
    .B(_09167_),
    .Y(_02393_));
 sky130_fd_sc_hd__nor2_1 _22915_ (.A(net1139),
    .B(_09167_),
    .Y(_02394_));
 sky130_fd_sc_hd__nor2_1 _22916_ (.A(_05011_),
    .B(_09167_),
    .Y(_02395_));
 sky130_fd_sc_hd__nor2_1 _22917_ (.A(_05020_),
    .B(_09167_),
    .Y(_02396_));
 sky130_fd_sc_hd__nor2_1 _22918_ (.A(_05029_),
    .B(_09167_),
    .Y(_02397_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_662 ();
 sky130_fd_sc_hd__nor2_1 _22920_ (.A(net1138),
    .B(_09167_),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _22921_ (.A(net1143),
    .B(_09167_),
    .Y(_02399_));
 sky130_fd_sc_hd__nor2_1 _22922_ (.A(_04801_),
    .B(_09167_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _22923_ (.A(_05060_),
    .B(_09167_),
    .Y(_02401_));
 sky130_fd_sc_hd__nor2_1 _22924_ (.A(_08895_),
    .B(_09167_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_1 _22925_ (.A(_04808_),
    .B(_09167_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _22926_ (.A(_04817_),
    .B(_09167_),
    .Y(_02404_));
 sky130_fd_sc_hd__nor2_1 _22927_ (.A(_04826_),
    .B(_09167_),
    .Y(_02405_));
 sky130_fd_sc_hd__nor2_1 _22928_ (.A(_04834_),
    .B(_09167_),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _22929_ (.A(_04843_),
    .B(_09167_),
    .Y(_02407_));
 sky130_fd_sc_hd__nor2_1 _22930_ (.A(_04852_),
    .B(_09167_),
    .Y(_02408_));
 sky130_fd_sc_hd__nor2_1 _22931_ (.A(_04860_),
    .B(_09167_),
    .Y(_02409_));
 sky130_fd_sc_hd__nand2_8 _22932_ (.A(_09830_),
    .B(_05474_),
    .Y(_09171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_661 ();
 sky130_fd_sc_hd__nor2_1 _22934_ (.A(_05118_),
    .B(_09171_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor2_1 _22935_ (.A(_05192_),
    .B(_09171_),
    .Y(_02411_));
 sky130_fd_sc_hd__nor2_1 _22936_ (.A(_05204_),
    .B(_09171_),
    .Y(_02412_));
 sky130_fd_sc_hd__nor2_1 _22937_ (.A(_05214_),
    .B(_09171_),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _22938_ (.A(_05221_),
    .B(_09171_),
    .Y(_02414_));
 sky130_fd_sc_hd__nor2_1 _22939_ (.A(net1136),
    .B(_09171_),
    .Y(_02415_));
 sky130_fd_sc_hd__nor2_1 _22940_ (.A(_05238_),
    .B(_09171_),
    .Y(_02416_));
 sky130_fd_sc_hd__nor2_1 _22941_ (.A(_05247_),
    .B(_09171_),
    .Y(_02417_));
 sky130_fd_sc_hd__nor2_1 _22942_ (.A(_05258_),
    .B(_09171_),
    .Y(_02418_));
 sky130_fd_sc_hd__nor2_1 _22943_ (.A(net1102),
    .B(_09171_),
    .Y(_02419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_660 ();
 sky130_fd_sc_hd__nor2_1 _22945_ (.A(_05280_),
    .B(_09171_),
    .Y(_02420_));
 sky130_fd_sc_hd__nor2_1 _22946_ (.A(_05122_),
    .B(_09171_),
    .Y(_02421_));
 sky130_fd_sc_hd__nor2_1 _22947_ (.A(_05291_),
    .B(_09171_),
    .Y(_02422_));
 sky130_fd_sc_hd__nor2_1 _22948_ (.A(_05301_),
    .B(_09171_),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_1 _22949_ (.A(_05309_),
    .B(_09171_),
    .Y(_02424_));
 sky130_fd_sc_hd__nor2_1 _22950_ (.A(_05320_),
    .B(_09171_),
    .Y(_02425_));
 sky130_fd_sc_hd__nor2_1 _22951_ (.A(net1100),
    .B(_09171_),
    .Y(_02426_));
 sky130_fd_sc_hd__nor2_1 _22952_ (.A(_05339_),
    .B(_09171_),
    .Y(_02427_));
 sky130_fd_sc_hd__nor2_1 _22953_ (.A(_05347_),
    .B(_09171_),
    .Y(_02428_));
 sky130_fd_sc_hd__nor2_1 _22954_ (.A(_05358_),
    .B(_09171_),
    .Y(_02429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_659 ();
 sky130_fd_sc_hd__nor2_1 _22956_ (.A(net1101),
    .B(_09171_),
    .Y(_02430_));
 sky130_fd_sc_hd__nor2_1 _22957_ (.A(_05380_),
    .B(_09171_),
    .Y(_02431_));
 sky130_fd_sc_hd__nor2_1 _22958_ (.A(_05126_),
    .B(_09171_),
    .Y(_02432_));
 sky130_fd_sc_hd__nor2_1 _22959_ (.A(net1129),
    .B(_09171_),
    .Y(_02433_));
 sky130_fd_sc_hd__nor2_1 _22960_ (.A(net1042),
    .B(_09171_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_1 _22961_ (.A(_05132_),
    .B(_09171_),
    .Y(_02435_));
 sky130_fd_sc_hd__nor2_1 _22962_ (.A(_05140_),
    .B(_09171_),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _22963_ (.A(_05149_),
    .B(_09171_),
    .Y(_02437_));
 sky130_fd_sc_hd__nor2_1 _22964_ (.A(_05157_),
    .B(_09171_),
    .Y(_02438_));
 sky130_fd_sc_hd__nor2_1 _22965_ (.A(_05166_),
    .B(_09171_),
    .Y(_02439_));
 sky130_fd_sc_hd__nor2_1 _22966_ (.A(_05173_),
    .B(_09171_),
    .Y(_02440_));
 sky130_fd_sc_hd__nor2_1 _22967_ (.A(_05183_),
    .B(_09171_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_8 _22968_ (.A(_09778_),
    .B(_05516_),
    .Y(_09175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_658 ();
 sky130_fd_sc_hd__nor2_1 _22970_ (.A(_04790_),
    .B(_09175_),
    .Y(_02442_));
 sky130_fd_sc_hd__nor2_1 _22971_ (.A(_04871_),
    .B(_09175_),
    .Y(_02443_));
 sky130_fd_sc_hd__nor2_1 _22972_ (.A(_04883_),
    .B(_09175_),
    .Y(_02444_));
 sky130_fd_sc_hd__nor2_1 _22973_ (.A(_04892_),
    .B(_09175_),
    .Y(_02445_));
 sky130_fd_sc_hd__nor2_1 _22974_ (.A(_04899_),
    .B(_09175_),
    .Y(_02446_));
 sky130_fd_sc_hd__nor2_1 _22975_ (.A(_04906_),
    .B(_09175_),
    .Y(_02447_));
 sky130_fd_sc_hd__nor2_1 _22976_ (.A(_04913_),
    .B(_09175_),
    .Y(_02448_));
 sky130_fd_sc_hd__nor2_1 _22977_ (.A(_04923_),
    .B(_09175_),
    .Y(_02449_));
 sky130_fd_sc_hd__nor2_1 _22978_ (.A(_04932_),
    .B(_09175_),
    .Y(_02450_));
 sky130_fd_sc_hd__nor2_1 _22979_ (.A(_04939_),
    .B(_09175_),
    .Y(_02451_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_657 ();
 sky130_fd_sc_hd__nor2_1 _22981_ (.A(_04951_),
    .B(_09175_),
    .Y(_02452_));
 sky130_fd_sc_hd__nor2_1 _22982_ (.A(_04794_),
    .B(_09175_),
    .Y(_02453_));
 sky130_fd_sc_hd__nor2_1 _22983_ (.A(_04960_),
    .B(_09175_),
    .Y(_02454_));
 sky130_fd_sc_hd__nor2_1 _22984_ (.A(_04974_),
    .B(_09175_),
    .Y(_02455_));
 sky130_fd_sc_hd__nor2_1 _22985_ (.A(_04984_),
    .B(_09175_),
    .Y(_02456_));
 sky130_fd_sc_hd__nor2_1 _22986_ (.A(_04990_),
    .B(_09175_),
    .Y(_02457_));
 sky130_fd_sc_hd__nor2_1 _22987_ (.A(net1139),
    .B(_09175_),
    .Y(_02458_));
 sky130_fd_sc_hd__nor2_1 _22988_ (.A(_05011_),
    .B(_09175_),
    .Y(_02459_));
 sky130_fd_sc_hd__nor2_1 _22989_ (.A(_05020_),
    .B(_09175_),
    .Y(_02460_));
 sky130_fd_sc_hd__nor2_1 _22990_ (.A(_05029_),
    .B(_09175_),
    .Y(_02461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_656 ();
 sky130_fd_sc_hd__nor2_1 _22992_ (.A(net1138),
    .B(_09175_),
    .Y(_02462_));
 sky130_fd_sc_hd__nor2_1 _22993_ (.A(_05044_),
    .B(_09175_),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _22994_ (.A(_04801_),
    .B(_09175_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor2_1 _22995_ (.A(_05060_),
    .B(_09175_),
    .Y(_02465_));
 sky130_fd_sc_hd__nor2_1 _22996_ (.A(_08895_),
    .B(_09175_),
    .Y(_02466_));
 sky130_fd_sc_hd__nor2_1 _22997_ (.A(_04808_),
    .B(_09175_),
    .Y(_02467_));
 sky130_fd_sc_hd__nor2_1 _22998_ (.A(_04817_),
    .B(_09175_),
    .Y(_02468_));
 sky130_fd_sc_hd__nor2_1 _22999_ (.A(_04826_),
    .B(_09175_),
    .Y(_02469_));
 sky130_fd_sc_hd__nor2_1 _23000_ (.A(_04834_),
    .B(_09175_),
    .Y(_02470_));
 sky130_fd_sc_hd__nor2_1 _23001_ (.A(_04843_),
    .B(_09175_),
    .Y(_02471_));
 sky130_fd_sc_hd__nor2_1 _23002_ (.A(_04852_),
    .B(_09175_),
    .Y(_02472_));
 sky130_fd_sc_hd__nor2_1 _23003_ (.A(_04860_),
    .B(_09175_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand2_8 _23004_ (.A(_09830_),
    .B(_05557_),
    .Y(_09179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_655 ();
 sky130_fd_sc_hd__nor2_1 _23006_ (.A(_05118_),
    .B(_09179_),
    .Y(_02474_));
 sky130_fd_sc_hd__nor2_1 _23007_ (.A(_05192_),
    .B(_09179_),
    .Y(_02475_));
 sky130_fd_sc_hd__nor2_1 _23008_ (.A(_05204_),
    .B(_09179_),
    .Y(_02476_));
 sky130_fd_sc_hd__nor2_1 _23009_ (.A(_05214_),
    .B(_09179_),
    .Y(_02477_));
 sky130_fd_sc_hd__nor2_1 _23010_ (.A(_05221_),
    .B(_09179_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_1 _23011_ (.A(net1136),
    .B(_09179_),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _23012_ (.A(_05238_),
    .B(_09179_),
    .Y(_02480_));
 sky130_fd_sc_hd__nor2_1 _23013_ (.A(net1135),
    .B(_09179_),
    .Y(_02481_));
 sky130_fd_sc_hd__nor2_1 _23014_ (.A(_05258_),
    .B(_09179_),
    .Y(_02482_));
 sky130_fd_sc_hd__nor2_1 _23015_ (.A(net1102),
    .B(_09179_),
    .Y(_02483_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_654 ();
 sky130_fd_sc_hd__nor2_1 _23017_ (.A(_05280_),
    .B(_09179_),
    .Y(_02484_));
 sky130_fd_sc_hd__nor2_1 _23018_ (.A(_05122_),
    .B(_09179_),
    .Y(_02485_));
 sky130_fd_sc_hd__nor2_1 _23019_ (.A(_05291_),
    .B(_09179_),
    .Y(_02486_));
 sky130_fd_sc_hd__nor2_1 _23020_ (.A(_05301_),
    .B(_09179_),
    .Y(_02487_));
 sky130_fd_sc_hd__nor2_1 _23021_ (.A(_05309_),
    .B(_09179_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_1 _23022_ (.A(_05320_),
    .B(_09179_),
    .Y(_02489_));
 sky130_fd_sc_hd__nor2_1 _23023_ (.A(net1100),
    .B(_09179_),
    .Y(_02490_));
 sky130_fd_sc_hd__nor2_1 _23024_ (.A(_05339_),
    .B(_09179_),
    .Y(_02491_));
 sky130_fd_sc_hd__nor2_1 _23025_ (.A(_05347_),
    .B(_09179_),
    .Y(_02492_));
 sky130_fd_sc_hd__nor2_1 _23026_ (.A(_05358_),
    .B(_09179_),
    .Y(_02493_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_653 ();
 sky130_fd_sc_hd__nor2_1 _23028_ (.A(net1142),
    .B(_09179_),
    .Y(_02494_));
 sky130_fd_sc_hd__nor2_1 _23029_ (.A(_05380_),
    .B(_09179_),
    .Y(_02495_));
 sky130_fd_sc_hd__nor2_1 _23030_ (.A(_05126_),
    .B(_09179_),
    .Y(_02496_));
 sky130_fd_sc_hd__nor2_1 _23031_ (.A(net1134),
    .B(_09179_),
    .Y(_02497_));
 sky130_fd_sc_hd__nor2_1 _23032_ (.A(net1042),
    .B(_09179_),
    .Y(_02498_));
 sky130_fd_sc_hd__nor2_1 _23033_ (.A(_05132_),
    .B(_09179_),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_1 _23034_ (.A(_05140_),
    .B(_09179_),
    .Y(_02500_));
 sky130_fd_sc_hd__nor2_1 _23035_ (.A(_05149_),
    .B(_09179_),
    .Y(_02501_));
 sky130_fd_sc_hd__nor2_1 _23036_ (.A(_05157_),
    .B(_09179_),
    .Y(_02502_));
 sky130_fd_sc_hd__nor2_1 _23037_ (.A(_05166_),
    .B(_09179_),
    .Y(_02503_));
 sky130_fd_sc_hd__nor2_1 _23038_ (.A(_05173_),
    .B(_09179_),
    .Y(_02504_));
 sky130_fd_sc_hd__nor2_1 _23039_ (.A(_05183_),
    .B(_09179_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_8 _23040_ (.A(_09778_),
    .B(_05598_),
    .Y(_09183_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_652 ();
 sky130_fd_sc_hd__nor2_1 _23042_ (.A(_04790_),
    .B(_09183_),
    .Y(_02506_));
 sky130_fd_sc_hd__nor2_1 _23043_ (.A(_04871_),
    .B(_09183_),
    .Y(_02507_));
 sky130_fd_sc_hd__nor2_1 _23044_ (.A(_04883_),
    .B(_09183_),
    .Y(_02508_));
 sky130_fd_sc_hd__nor2_1 _23045_ (.A(_04892_),
    .B(_09183_),
    .Y(_02509_));
 sky130_fd_sc_hd__nor2_1 _23046_ (.A(_04899_),
    .B(_09183_),
    .Y(_02510_));
 sky130_fd_sc_hd__nor2_1 _23047_ (.A(_04906_),
    .B(_09183_),
    .Y(_02511_));
 sky130_fd_sc_hd__nor2_1 _23048_ (.A(_04913_),
    .B(_09183_),
    .Y(_02512_));
 sky130_fd_sc_hd__nor2_1 _23049_ (.A(_04923_),
    .B(_09183_),
    .Y(_02513_));
 sky130_fd_sc_hd__nor2_1 _23050_ (.A(_04932_),
    .B(_09183_),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _23051_ (.A(_04939_),
    .B(_09183_),
    .Y(_02515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_651 ();
 sky130_fd_sc_hd__nor2_1 _23053_ (.A(_04951_),
    .B(_09183_),
    .Y(_02516_));
 sky130_fd_sc_hd__nor2_1 _23054_ (.A(_04794_),
    .B(_09183_),
    .Y(_02517_));
 sky130_fd_sc_hd__nor2_1 _23055_ (.A(_04960_),
    .B(_09183_),
    .Y(_02518_));
 sky130_fd_sc_hd__nor2_1 _23056_ (.A(_04974_),
    .B(_09183_),
    .Y(_02519_));
 sky130_fd_sc_hd__nor2_1 _23057_ (.A(_04984_),
    .B(_09183_),
    .Y(_02520_));
 sky130_fd_sc_hd__nor2_1 _23058_ (.A(_04990_),
    .B(_09183_),
    .Y(_02521_));
 sky130_fd_sc_hd__nor2_1 _23059_ (.A(net1139),
    .B(_09183_),
    .Y(_02522_));
 sky130_fd_sc_hd__nor2_1 _23060_ (.A(_05011_),
    .B(_09183_),
    .Y(_02523_));
 sky130_fd_sc_hd__nor2_1 _23061_ (.A(_05020_),
    .B(_09183_),
    .Y(_02524_));
 sky130_fd_sc_hd__nor2_1 _23062_ (.A(_05029_),
    .B(_09183_),
    .Y(_02525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_650 ();
 sky130_fd_sc_hd__nor2_1 _23064_ (.A(net1138),
    .B(_09183_),
    .Y(_02526_));
 sky130_fd_sc_hd__nor2_1 _23065_ (.A(net1143),
    .B(_09183_),
    .Y(_02527_));
 sky130_fd_sc_hd__nor2_1 _23066_ (.A(_04801_),
    .B(_09183_),
    .Y(_02528_));
 sky130_fd_sc_hd__nor2_1 _23067_ (.A(_05060_),
    .B(_09183_),
    .Y(_02529_));
 sky130_fd_sc_hd__nor2_1 _23068_ (.A(_08895_),
    .B(_09183_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_1 _23069_ (.A(_04808_),
    .B(_09183_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_1 _23070_ (.A(_04817_),
    .B(_09183_),
    .Y(_02532_));
 sky130_fd_sc_hd__nor2_1 _23071_ (.A(_04826_),
    .B(_09183_),
    .Y(_02533_));
 sky130_fd_sc_hd__nor2_1 _23072_ (.A(_04834_),
    .B(_09183_),
    .Y(_02534_));
 sky130_fd_sc_hd__nor2_1 _23073_ (.A(_04843_),
    .B(_09183_),
    .Y(_02535_));
 sky130_fd_sc_hd__nor2_1 _23074_ (.A(_04852_),
    .B(_09183_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor2_1 _23075_ (.A(_04860_),
    .B(_09183_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2b_4 _23076_ (.A_N(_09726_),
    .B(_09731_),
    .Y(_09187_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_649 ();
 sky130_fd_sc_hd__nor2_1 _23078_ (.A(_05118_),
    .B(_09187_),
    .Y(_02538_));
 sky130_fd_sc_hd__nor2_1 _23079_ (.A(_05192_),
    .B(_09187_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor2_1 _23080_ (.A(_05204_),
    .B(_09187_),
    .Y(_02540_));
 sky130_fd_sc_hd__nor2_1 _23081_ (.A(_05214_),
    .B(_09187_),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _23082_ (.A(_05221_),
    .B(_09187_),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_1 _23083_ (.A(net1136),
    .B(_09187_),
    .Y(_02543_));
 sky130_fd_sc_hd__nor2_1 _23084_ (.A(_05238_),
    .B(_09187_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _23085_ (.A(net1135),
    .B(_09187_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _23086_ (.A(_05258_),
    .B(_09187_),
    .Y(_02546_));
 sky130_fd_sc_hd__nor2_1 _23087_ (.A(net1102),
    .B(_09187_),
    .Y(_02547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_648 ();
 sky130_fd_sc_hd__nor2_1 _23089_ (.A(_05280_),
    .B(_09187_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor2_1 _23090_ (.A(_05122_),
    .B(_09187_),
    .Y(_02549_));
 sky130_fd_sc_hd__nor2_1 _23091_ (.A(_05291_),
    .B(_09187_),
    .Y(_02550_));
 sky130_fd_sc_hd__nor2_1 _23092_ (.A(_05301_),
    .B(_09187_),
    .Y(_02551_));
 sky130_fd_sc_hd__nor2_1 _23093_ (.A(_05309_),
    .B(_09187_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _23094_ (.A(_05320_),
    .B(_09187_),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _23095_ (.A(net1100),
    .B(_09187_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_1 _23096_ (.A(_05339_),
    .B(_09187_),
    .Y(_02555_));
 sky130_fd_sc_hd__nor2_1 _23097_ (.A(_05347_),
    .B(_09187_),
    .Y(_02556_));
 sky130_fd_sc_hd__nor2_1 _23098_ (.A(_05358_),
    .B(_09187_),
    .Y(_02557_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_647 ();
 sky130_fd_sc_hd__nor2_1 _23100_ (.A(net1142),
    .B(_09187_),
    .Y(_02558_));
 sky130_fd_sc_hd__nor2_1 _23101_ (.A(_05380_),
    .B(_09187_),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2_1 _23102_ (.A(_05126_),
    .B(_09187_),
    .Y(_02560_));
 sky130_fd_sc_hd__nor2_1 _23103_ (.A(net1129),
    .B(_09187_),
    .Y(_02561_));
 sky130_fd_sc_hd__nor2_1 _23104_ (.A(_05430_),
    .B(_09187_),
    .Y(_02562_));
 sky130_fd_sc_hd__nor2_1 _23105_ (.A(_05132_),
    .B(_09187_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_1 _23106_ (.A(_05140_),
    .B(_09187_),
    .Y(_02564_));
 sky130_fd_sc_hd__nor2_1 _23107_ (.A(_05149_),
    .B(_09187_),
    .Y(_02565_));
 sky130_fd_sc_hd__nor2_1 _23108_ (.A(_05157_),
    .B(_09187_),
    .Y(_02566_));
 sky130_fd_sc_hd__nor2_1 _23109_ (.A(_05166_),
    .B(_09187_),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_1 _23110_ (.A(_05173_),
    .B(_09187_),
    .Y(_02568_));
 sky130_fd_sc_hd__nor2_1 _23111_ (.A(_05183_),
    .B(_09187_),
    .Y(_02569_));
 sky130_fd_sc_hd__nor2b_4 _23112_ (.A(net349),
    .B_N(\hash.CA2.b_dash[0] ),
    .Y(\hash.CA1.d[0] ));
 sky130_fd_sc_hd__clkinv_1 _23113_ (.A(_13581_),
    .Y(_09191_));
 sky130_fd_sc_hd__inv_2 _23114_ (.A(_13573_),
    .Y(_09192_));
 sky130_fd_sc_hd__inv_1 _23115_ (.A(_13565_),
    .Y(_09193_));
 sky130_fd_sc_hd__inv_1 _23116_ (.A(_13557_),
    .Y(_09194_));
 sky130_fd_sc_hd__nor2b_2 _23117_ (.A(_12882_),
    .B_N(_13554_),
    .Y(_09195_));
 sky130_fd_sc_hd__o21ai_2 _23118_ (.A1(_13553_),
    .A2(_09195_),
    .B1(_13558_),
    .Y(_09196_));
 sky130_fd_sc_hd__a21boi_2 _23119_ (.A1(_09194_),
    .A2(_09196_),
    .B1_N(_13562_),
    .Y(_09197_));
 sky130_fd_sc_hd__o21ai_2 _23120_ (.A1(_13561_),
    .A2(_09197_),
    .B1(_13566_),
    .Y(_09198_));
 sky130_fd_sc_hd__a21boi_2 _23121_ (.A1(_09193_),
    .A2(_09198_),
    .B1_N(_13570_),
    .Y(_09199_));
 sky130_fd_sc_hd__o21ai_2 _23122_ (.A1(_13569_),
    .A2(_09199_),
    .B1(_13574_),
    .Y(_09200_));
 sky130_fd_sc_hd__a21boi_2 _23123_ (.A1(_09192_),
    .A2(_09200_),
    .B1_N(_13578_),
    .Y(_09201_));
 sky130_fd_sc_hd__o21ai_2 _23124_ (.A1(_13577_),
    .A2(_09201_),
    .B1(_13582_),
    .Y(_09202_));
 sky130_fd_sc_hd__a21boi_4 _23125_ (.A1(_09191_),
    .A2(_09202_),
    .B1_N(_13586_),
    .Y(_09203_));
 sky130_fd_sc_hd__nand2_1 _23126_ (.A(_09191_),
    .B(_09202_),
    .Y(_09204_));
 sky130_fd_sc_hd__nor2_1 _23127_ (.A(_13586_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__nor2_1 _23128_ (.A(_09203_),
    .B(_09205_),
    .Y(\hash.CA1.p1[10] ));
 sky130_fd_sc_hd__o21a_1 _23129_ (.A1(_13582_),
    .A2(_13581_),
    .B1(_13586_),
    .X(_09206_));
 sky130_fd_sc_hd__nor2_2 _23130_ (.A(_13585_),
    .B(_09206_),
    .Y(_09207_));
 sky130_fd_sc_hd__inv_1 _23131_ (.A(_13558_),
    .Y(_09208_));
 sky130_fd_sc_hd__a21o_1 _23132_ (.A1(_14204_),
    .A2(_13550_),
    .B1(_13549_),
    .X(_09209_));
 sky130_fd_sc_hd__a21oi_2 _23133_ (.A1(_13554_),
    .A2(_09209_),
    .B1(_13553_),
    .Y(_09210_));
 sky130_fd_sc_hd__nor3_1 _23134_ (.A(_13557_),
    .B(_13561_),
    .C(_13565_),
    .Y(_09211_));
 sky130_fd_sc_hd__o21ai_1 _23135_ (.A1(_09208_),
    .A2(_09210_),
    .B1(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__o21ai_0 _23136_ (.A1(_13562_),
    .A2(_13561_),
    .B1(_13566_),
    .Y(_09213_));
 sky130_fd_sc_hd__nand2_1 _23137_ (.A(_09193_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__and3_4 _23138_ (.A(_13570_),
    .B(_13574_),
    .C(_13578_),
    .X(_09215_));
 sky130_fd_sc_hd__and3_4 _23139_ (.A(_09212_),
    .B(_09214_),
    .C(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__nand2_1 _23140_ (.A(_13574_),
    .B(_13569_),
    .Y(_09217_));
 sky130_fd_sc_hd__nand2_1 _23141_ (.A(_09192_),
    .B(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__a21oi_1 _23142_ (.A1(_13578_),
    .A2(_09218_),
    .B1(_13577_),
    .Y(_09219_));
 sky130_fd_sc_hd__nor4b_4 _23143_ (.A(_13581_),
    .B(_13585_),
    .C(_09216_),
    .D_N(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__nor2_2 _23144_ (.A(_09207_),
    .B(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__xor2_1 _23145_ (.A(_13590_),
    .B(_09221_),
    .X(\hash.CA1.p1[11] ));
 sky130_fd_sc_hd__o21a_1 _23146_ (.A1(_13585_),
    .A2(_09203_),
    .B1(_13590_),
    .X(_09222_));
 sky130_fd_sc_hd__nor2_1 _23147_ (.A(_13589_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__xnor2_1 _23148_ (.A(_13594_),
    .B(_09223_),
    .Y(\hash.CA1.p1[12] ));
 sky130_fd_sc_hd__a21o_4 _23149_ (.A1(_13594_),
    .A2(_13589_),
    .B1(_13593_),
    .X(_09224_));
 sky130_fd_sc_hd__and3_4 _23150_ (.A(_13590_),
    .B(_13594_),
    .C(_09221_),
    .X(_09225_));
 sky130_fd_sc_hd__nor2_1 _23151_ (.A(_09224_),
    .B(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__xnor2_1 _23152_ (.A(_13598_),
    .B(_09226_),
    .Y(\hash.CA1.p1[13] ));
 sky130_fd_sc_hd__or3_4 _23153_ (.A(_13585_),
    .B(_13597_),
    .C(_09224_),
    .X(_09227_));
 sky130_fd_sc_hd__a211oi_1 _23154_ (.A1(_13590_),
    .A2(_13594_),
    .B1(_13597_),
    .C1(_09224_),
    .Y(_09228_));
 sky130_fd_sc_hd__nor2_1 _23155_ (.A(_13598_),
    .B(_13597_),
    .Y(_09229_));
 sky130_fd_sc_hd__nor2_1 _23156_ (.A(_09228_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__o21ai_4 _23157_ (.A1(_09227_),
    .A2(_09203_),
    .B1(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__xnor2_1 _23158_ (.A(_13602_),
    .B(_09231_),
    .Y(\hash.CA1.p1[14] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_646 ();
 sky130_fd_sc_hd__o21ai_2 _23160_ (.A1(_09225_),
    .A2(_09224_),
    .B1(_13598_),
    .Y(_09233_));
 sky130_fd_sc_hd__nand2b_1 _23161_ (.A_N(_13597_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__a21oi_2 _23162_ (.A1(_09234_),
    .A2(_13602_),
    .B1(_13601_),
    .Y(_09235_));
 sky130_fd_sc_hd__xnor2_1 _23163_ (.A(_13606_),
    .B(_09235_),
    .Y(\hash.CA1.p1[15] ));
 sky130_fd_sc_hd__inv_1 _23164_ (.A(_13602_),
    .Y(_09236_));
 sky130_fd_sc_hd__o21bai_4 _23165_ (.A1(_09231_),
    .A2(_09236_),
    .B1_N(_13601_),
    .Y(_09237_));
 sky130_fd_sc_hd__a21oi_2 _23166_ (.A1(_09237_),
    .A2(_13606_),
    .B1(_13605_),
    .Y(_09238_));
 sky130_fd_sc_hd__xnor2_1 _23167_ (.A(_13610_),
    .B(_09238_),
    .Y(\hash.CA1.p1[16] ));
 sky130_fd_sc_hd__inv_1 _23168_ (.A(_13606_),
    .Y(_09239_));
 sky130_fd_sc_hd__o21bai_1 _23169_ (.A1(_09239_),
    .A2(_09235_),
    .B1_N(_13605_),
    .Y(_09240_));
 sky130_fd_sc_hd__a21oi_1 _23170_ (.A1(_09240_),
    .A2(_13610_),
    .B1(_13609_),
    .Y(_09241_));
 sky130_fd_sc_hd__xnor2_1 _23171_ (.A(_09241_),
    .B(_13614_),
    .Y(\hash.CA1.p1[17] ));
 sky130_fd_sc_hd__inv_1 _23172_ (.A(_13614_),
    .Y(_09242_));
 sky130_fd_sc_hd__and2_0 _23173_ (.A(_13610_),
    .B(_13605_),
    .X(_09243_));
 sky130_fd_sc_hd__a311oi_2 _23174_ (.A1(_13606_),
    .A2(_09237_),
    .A3(_13610_),
    .B1(_09243_),
    .C1(_13609_),
    .Y(_09244_));
 sky130_fd_sc_hd__o21bai_1 _23175_ (.A1(_09244_),
    .A2(_09242_),
    .B1_N(_13613_),
    .Y(_09245_));
 sky130_fd_sc_hd__xor2_1 _23176_ (.A(_09245_),
    .B(_13618_),
    .X(\hash.CA1.p1[18] ));
 sky130_fd_sc_hd__and3_4 _23177_ (.A(_13610_),
    .B(_13614_),
    .C(_13618_),
    .X(_09246_));
 sky130_fd_sc_hd__a21o_1 _23178_ (.A1(_13606_),
    .A2(_13601_),
    .B1(_13605_),
    .X(_09247_));
 sky130_fd_sc_hd__a21o_1 _23179_ (.A1(_13614_),
    .A2(_13609_),
    .B1(_13613_),
    .X(_09248_));
 sky130_fd_sc_hd__a221oi_4 _23180_ (.A1(_09246_),
    .A2(_09247_),
    .B1(_09248_),
    .B2(_13618_),
    .C1(_13617_),
    .Y(_09249_));
 sky130_fd_sc_hd__clkinv_2 _23181_ (.A(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand3_1 _23182_ (.A(_13602_),
    .B(_13606_),
    .C(_09246_),
    .Y(_09251_));
 sky130_fd_sc_hd__a21oi_1 _23183_ (.A1(_13598_),
    .A2(_09224_),
    .B1(_13597_),
    .Y(_09252_));
 sky130_fd_sc_hd__nor2_1 _23184_ (.A(_09251_),
    .B(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__and3_4 _23185_ (.A(_13602_),
    .B(_13606_),
    .C(_09246_),
    .X(_09254_));
 sky130_fd_sc_hd__nand4_1 _23186_ (.A(_09254_),
    .B(_13590_),
    .C(_13594_),
    .D(_13598_),
    .Y(_09255_));
 sky130_fd_sc_hd__nor3_4 _23187_ (.A(_09207_),
    .B(_09220_),
    .C(_09255_),
    .Y(_09256_));
 sky130_fd_sc_hd__nor3_1 _23188_ (.A(_09250_),
    .B(_09253_),
    .C(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__xnor2_1 _23189_ (.A(_13622_),
    .B(_09257_),
    .Y(\hash.CA1.p1[19] ));
 sky130_fd_sc_hd__o21ai_2 _23190_ (.A1(_09251_),
    .A2(_09231_),
    .B1(_09249_),
    .Y(_09258_));
 sky130_fd_sc_hd__a21oi_2 _23191_ (.A1(_09258_),
    .A2(_13622_),
    .B1(_13621_),
    .Y(_09259_));
 sky130_fd_sc_hd__xnor2_1 _23192_ (.A(_13626_),
    .B(_09259_),
    .Y(\hash.CA1.p1[20] ));
 sky130_fd_sc_hd__o31ai_4 _23193_ (.A1(_09250_),
    .A2(_09253_),
    .A3(_09256_),
    .B1(_13622_),
    .Y(_09260_));
 sky130_fd_sc_hd__nor2_2 _23194_ (.A(_13621_),
    .B(_13625_),
    .Y(_09261_));
 sky130_fd_sc_hd__nor2_1 _23195_ (.A(_13626_),
    .B(_13625_),
    .Y(_09262_));
 sky130_fd_sc_hd__a21oi_4 _23196_ (.A1(_09261_),
    .A2(_09260_),
    .B1(_09262_),
    .Y(_09263_));
 sky130_fd_sc_hd__xor2_1 _23197_ (.A(_13630_),
    .B(_09263_),
    .X(\hash.CA1.p1[21] ));
 sky130_fd_sc_hd__and3_4 _23198_ (.A(_13622_),
    .B(_13626_),
    .C(_09254_),
    .X(_09264_));
 sky130_fd_sc_hd__o211ai_1 _23199_ (.A1(_09203_),
    .A2(_09227_),
    .B1(_09230_),
    .C1(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__and3_1 _23200_ (.A(_13622_),
    .B(_13626_),
    .C(_09250_),
    .X(_09266_));
 sky130_fd_sc_hd__a21oi_2 _23201_ (.A1(_13626_),
    .A2(_13621_),
    .B1(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__nand3b_1 _23202_ (.A_N(_13625_),
    .B(_09267_),
    .C(_09265_),
    .Y(_09268_));
 sky130_fd_sc_hd__a21oi_2 _23203_ (.A1(_09268_),
    .A2(_13630_),
    .B1(_13629_),
    .Y(_09269_));
 sky130_fd_sc_hd__xnor2_1 _23204_ (.A(_13634_),
    .B(_09269_),
    .Y(\hash.CA1.p1[22] ));
 sky130_fd_sc_hd__a21o_1 _23205_ (.A1(_09263_),
    .A2(_13630_),
    .B1(_13629_),
    .X(_09270_));
 sky130_fd_sc_hd__a21oi_2 _23206_ (.A1(_09270_),
    .A2(_13634_),
    .B1(_13633_),
    .Y(_09271_));
 sky130_fd_sc_hd__xnor2_1 _23207_ (.A(_09271_),
    .B(_13638_),
    .Y(\hash.CA1.p1[23] ));
 sky130_fd_sc_hd__and3_4 _23208_ (.A(_13630_),
    .B(_13634_),
    .C(_13638_),
    .X(_09272_));
 sky130_fd_sc_hd__a21o_1 _23209_ (.A1(_13634_),
    .A2(_13629_),
    .B1(_13633_),
    .X(_09273_));
 sky130_fd_sc_hd__a21oi_2 _23210_ (.A1(_13638_),
    .A2(_09273_),
    .B1(_13637_),
    .Y(_09274_));
 sky130_fd_sc_hd__a21boi_2 _23211_ (.A1(_09268_),
    .A2(_09272_),
    .B1_N(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__xnor2_1 _23212_ (.A(_13642_),
    .B(_09275_),
    .Y(\hash.CA1.p1[24] ));
 sky130_fd_sc_hd__nand2_1 _23213_ (.A(_13642_),
    .B(_13646_),
    .Y(_09276_));
 sky130_fd_sc_hd__nand2_1 _23214_ (.A(_13646_),
    .B(_13641_),
    .Y(_09277_));
 sky130_fd_sc_hd__o21ai_0 _23215_ (.A1(_09274_),
    .A2(_09276_),
    .B1(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__a41o_4 _23216_ (.A1(_09263_),
    .A2(_13646_),
    .A3(_13642_),
    .A4(_09272_),
    .B1(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__nand2_1 _23217_ (.A(_09263_),
    .B(_09272_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_1 _23218_ (.A(_09274_),
    .B(_09280_),
    .Y(_09281_));
 sky130_fd_sc_hd__a211oi_2 _23219_ (.A1(_09281_),
    .A2(_13642_),
    .B1(_13641_),
    .C1(_13646_),
    .Y(_09282_));
 sky130_fd_sc_hd__nor2_1 _23220_ (.A(_09279_),
    .B(_09282_),
    .Y(\hash.CA1.p1[25] ));
 sky130_fd_sc_hd__nand4b_1 _23221_ (.A_N(_13625_),
    .B(_09265_),
    .C(_09267_),
    .D(_09274_),
    .Y(_09283_));
 sky130_fd_sc_hd__nand2b_1 _23222_ (.A_N(_09272_),
    .B(_09274_),
    .Y(_09284_));
 sky130_fd_sc_hd__a31o_1 _23223_ (.A1(_13642_),
    .A2(_09283_),
    .A3(_09284_),
    .B1(_13641_),
    .X(_09285_));
 sky130_fd_sc_hd__a21oi_2 _23224_ (.A1(_13646_),
    .A2(_09285_),
    .B1(_13645_),
    .Y(_09286_));
 sky130_fd_sc_hd__xnor2_1 _23225_ (.A(_09286_),
    .B(_13650_),
    .Y(\hash.CA1.p1[26] ));
 sky130_fd_sc_hd__o21a_1 _23226_ (.A1(_09279_),
    .A2(_13645_),
    .B1(_13650_),
    .X(_09287_));
 sky130_fd_sc_hd__nor2_2 _23227_ (.A(_13649_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__xnor2_2 _23228_ (.A(_09288_),
    .B(_13654_),
    .Y(\hash.CA1.p1[27] ));
 sky130_fd_sc_hd__a21o_1 _23229_ (.A1(_13638_),
    .A2(_13633_),
    .B1(_13637_),
    .X(_09289_));
 sky130_fd_sc_hd__a21oi_1 _23230_ (.A1(_13642_),
    .A2(_09289_),
    .B1(_13641_),
    .Y(_09290_));
 sky130_fd_sc_hd__nor2b_1 _23231_ (.A(_09290_),
    .B_N(_13646_),
    .Y(_09291_));
 sky130_fd_sc_hd__o21ai_0 _23232_ (.A1(_13645_),
    .A2(_09291_),
    .B1(_13650_),
    .Y(_09292_));
 sky130_fd_sc_hd__nand2b_1 _23233_ (.A_N(_13649_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__a21oi_1 _23234_ (.A1(_13654_),
    .A2(_09293_),
    .B1(_13653_),
    .Y(_09294_));
 sky130_fd_sc_hd__nor2_1 _23235_ (.A(_13625_),
    .B(_13629_),
    .Y(_09295_));
 sky130_fd_sc_hd__nand4_1 _23236_ (.A(net1123),
    .B(_09267_),
    .C(_09294_),
    .D(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__nand2_1 _23237_ (.A(_13634_),
    .B(_13638_),
    .Y(_09297_));
 sky130_fd_sc_hd__nand2_1 _23238_ (.A(_13650_),
    .B(_13654_),
    .Y(_09298_));
 sky130_fd_sc_hd__nor2_1 _23239_ (.A(_13630_),
    .B(_13629_),
    .Y(_09299_));
 sky130_fd_sc_hd__o41ai_1 _23240_ (.A1(_09297_),
    .A2(_09276_),
    .A3(_09298_),
    .A4(_09299_),
    .B1(_09294_),
    .Y(_09300_));
 sky130_fd_sc_hd__nand2_2 _23241_ (.A(_09296_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__xnor2_2 _23242_ (.A(_13658_),
    .B(_09301_),
    .Y(\hash.CA1.p1[28] ));
 sky130_fd_sc_hd__a21o_1 _23243_ (.A1(_13658_),
    .A2(_13653_),
    .B1(_13657_),
    .X(_09302_));
 sky130_fd_sc_hd__or4_4 _23244_ (.A(_13645_),
    .B(_13649_),
    .C(_09302_),
    .D(_09279_),
    .X(_09303_));
 sky130_fd_sc_hd__a21oi_1 _23245_ (.A1(_13654_),
    .A2(_13658_),
    .B1(_09302_),
    .Y(_09304_));
 sky130_fd_sc_hd__nor3_1 _23246_ (.A(_13650_),
    .B(_13649_),
    .C(_09302_),
    .Y(_09305_));
 sky130_fd_sc_hd__nor2_1 _23247_ (.A(_09304_),
    .B(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand2_4 _23248_ (.A(_09303_),
    .B(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__xnor2_2 _23249_ (.A(_13662_),
    .B(_09307_),
    .Y(\hash.CA1.p1[29] ));
 sky130_fd_sc_hd__xnor2_1 _23250_ (.A(_12882_),
    .B(_13554_),
    .Y(\hash.CA1.p1[2] ));
 sky130_fd_sc_hd__a31o_1 _23251_ (.A1(_13658_),
    .A2(_09296_),
    .A3(_09300_),
    .B1(_13657_),
    .X(_09308_));
 sky130_fd_sc_hd__a21oi_2 _23252_ (.A1(_09308_),
    .A2(_13662_),
    .B1(_13661_),
    .Y(_09309_));
 sky130_fd_sc_hd__xnor2_1 _23253_ (.A(_09309_),
    .B(_13666_),
    .Y(\hash.CA1.p1[30] ));
 sky130_fd_sc_hd__xor2_1 _23254_ (.A(_13241_),
    .B(_06073_),
    .X(_09310_));
 sky130_fd_sc_hd__xnor3_1 _23255_ (.A(\hash.CA2.b_dash[31] ),
    .B(_06248_),
    .C(_06266_),
    .X(_09311_));
 sky130_fd_sc_hd__maj3_1 _23256_ (.A(\hash.CA2.a_dash[31] ),
    .B(_04612_),
    .C(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__xnor2_1 _23257_ (.A(_09310_),
    .B(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__nor2_1 _23258_ (.A(net350),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__inv_1 _23259_ (.A(_13666_),
    .Y(_09315_));
 sky130_fd_sc_hd__a31oi_2 _23260_ (.A1(_09303_),
    .A2(_13662_),
    .A3(_09306_),
    .B1(_13661_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21bai_1 _23261_ (.A1(_09316_),
    .A2(_09315_),
    .B1_N(_13665_),
    .Y(_09317_));
 sky130_fd_sc_hd__xor2_1 _23262_ (.A(_09317_),
    .B(_06156_),
    .X(_09318_));
 sky130_fd_sc_hd__xnor2_1 _23263_ (.A(_09318_),
    .B(_09314_),
    .Y(\hash.CA1.p1[31] ));
 sky130_fd_sc_hd__xnor2_1 _23264_ (.A(_13558_),
    .B(_09210_),
    .Y(\hash.CA1.p1[3] ));
 sky130_fd_sc_hd__nand2_1 _23265_ (.A(_09194_),
    .B(_09196_),
    .Y(_09319_));
 sky130_fd_sc_hd__nor2_1 _23266_ (.A(_13562_),
    .B(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__nor2_2 _23267_ (.A(_09197_),
    .B(_09320_),
    .Y(\hash.CA1.p1[4] ));
 sky130_fd_sc_hd__o21ai_0 _23268_ (.A1(_09208_),
    .A2(_09210_),
    .B1(_09194_),
    .Y(_09321_));
 sky130_fd_sc_hd__a21oi_1 _23269_ (.A1(_13562_),
    .A2(_09321_),
    .B1(_13561_),
    .Y(_09322_));
 sky130_fd_sc_hd__xnor2_1 _23270_ (.A(_13566_),
    .B(_09322_),
    .Y(\hash.CA1.p1[5] ));
 sky130_fd_sc_hd__nand2_1 _23271_ (.A(_09193_),
    .B(_09198_),
    .Y(_09323_));
 sky130_fd_sc_hd__nor2_1 _23272_ (.A(_13570_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__nor2_1 _23273_ (.A(_09199_),
    .B(_09324_),
    .Y(\hash.CA1.p1[6] ));
 sky130_fd_sc_hd__a31oi_1 _23274_ (.A1(_13570_),
    .A2(_09212_),
    .A3(_09214_),
    .B1(_13569_),
    .Y(_09325_));
 sky130_fd_sc_hd__xnor2_1 _23275_ (.A(_13574_),
    .B(_09325_),
    .Y(\hash.CA1.p1[7] ));
 sky130_fd_sc_hd__nand2_1 _23276_ (.A(_09192_),
    .B(_09200_),
    .Y(_09326_));
 sky130_fd_sc_hd__nor2_1 _23277_ (.A(_13578_),
    .B(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__nor2_1 _23278_ (.A(_09201_),
    .B(_09327_),
    .Y(\hash.CA1.p1[8] ));
 sky130_fd_sc_hd__nand2b_1 _23279_ (.A_N(_09216_),
    .B(_09219_),
    .Y(_09328_));
 sky130_fd_sc_hd__xor2_1 _23280_ (.A(_13582_),
    .B(_09328_),
    .X(\hash.CA1.p1[9] ));
 sky130_fd_sc_hd__inv_1 _23281_ (.A(_14155_),
    .Y(_09329_));
 sky130_fd_sc_hd__inv_1 _23282_ (.A(_14147_),
    .Y(_09330_));
 sky130_fd_sc_hd__a21o_1 _23283_ (.A1(_14207_),
    .A2(_14131_),
    .B1(_14130_),
    .X(_09331_));
 sky130_fd_sc_hd__a21o_4 _23284_ (.A1(_14135_),
    .A2(_09331_),
    .B1(_14134_),
    .X(_09332_));
 sky130_fd_sc_hd__a21oi_1 _23285_ (.A1(_14139_),
    .A2(_09332_),
    .B1(_14138_),
    .Y(_09333_));
 sky130_fd_sc_hd__nor2b_1 _23286_ (.A(_09333_),
    .B_N(_14143_),
    .Y(_09334_));
 sky130_fd_sc_hd__nor2_2 _23287_ (.A(_14142_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__o21bai_1 _23288_ (.A1(_09330_),
    .A2(_09335_),
    .B1_N(_14146_),
    .Y(_09336_));
 sky130_fd_sc_hd__a21oi_2 _23289_ (.A1(_14151_),
    .A2(_09336_),
    .B1(_14150_),
    .Y(_09337_));
 sky130_fd_sc_hd__o21bai_1 _23290_ (.A1(_09329_),
    .A2(_09337_),
    .B1_N(_14154_),
    .Y(_09338_));
 sky130_fd_sc_hd__a21oi_1 _23291_ (.A1(_14158_),
    .A2(_09338_),
    .B1(_14157_),
    .Y(_09339_));
 sky130_fd_sc_hd__xnor2_2 _23292_ (.A(_14160_),
    .B(_09339_),
    .Y(\hash.CA1.p2[10] ));
 sky130_fd_sc_hd__a21o_1 _23293_ (.A1(_14158_),
    .A2(_14154_),
    .B1(_14157_),
    .X(_09340_));
 sky130_fd_sc_hd__a21o_4 _23294_ (.A1(_14160_),
    .A2(_09340_),
    .B1(_14159_),
    .X(_09341_));
 sky130_fd_sc_hd__nor2b_1 _23295_ (.A(_12885_),
    .B_N(_14135_),
    .Y(_09342_));
 sky130_fd_sc_hd__o21a_1 _23296_ (.A1(_14134_),
    .A2(_09342_),
    .B1(_14139_),
    .X(_09343_));
 sky130_fd_sc_hd__o21ai_2 _23297_ (.A1(_14138_),
    .A2(_09343_),
    .B1(_14143_),
    .Y(_09344_));
 sky130_fd_sc_hd__nor3_1 _23298_ (.A(_14142_),
    .B(_14146_),
    .C(_14150_),
    .Y(_09345_));
 sky130_fd_sc_hd__inv_1 _23299_ (.A(_14151_),
    .Y(_09346_));
 sky130_fd_sc_hd__nor2_1 _23300_ (.A(_14147_),
    .B(_14146_),
    .Y(_09347_));
 sky130_fd_sc_hd__nor2_1 _23301_ (.A(_09346_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__and3_4 _23302_ (.A(_14158_),
    .B(_14155_),
    .C(_14160_),
    .X(_09349_));
 sky130_fd_sc_hd__o21ai_2 _23303_ (.A1(_14150_),
    .A2(_09348_),
    .B1(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__a21oi_4 _23304_ (.A1(_09344_),
    .A2(_09345_),
    .B1(_09350_),
    .Y(_09351_));
 sky130_fd_sc_hd__nor2_2 _23305_ (.A(_09341_),
    .B(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__xnor2_2 _23306_ (.A(_14162_),
    .B(_09352_),
    .Y(\hash.CA1.p2[11] ));
 sky130_fd_sc_hd__a211oi_1 _23307_ (.A1(_14139_),
    .A2(_09332_),
    .B1(_14142_),
    .C1(_14138_),
    .Y(_09353_));
 sky130_fd_sc_hd__o2111ai_4 _23308_ (.A1(_14143_),
    .A2(_14142_),
    .B1(_14151_),
    .C1(_14147_),
    .D1(_09349_),
    .Y(_09354_));
 sky130_fd_sc_hd__a21o_1 _23309_ (.A1(_14151_),
    .A2(_14146_),
    .B1(_14150_),
    .X(_09355_));
 sky130_fd_sc_hd__a21oi_4 _23310_ (.A1(_09349_),
    .A2(_09355_),
    .B1(_09341_),
    .Y(_09356_));
 sky130_fd_sc_hd__o21ai_4 _23311_ (.A1(_09353_),
    .A2(_09354_),
    .B1(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__a21oi_1 _23312_ (.A1(_14162_),
    .A2(_09357_),
    .B1(_14161_),
    .Y(_09358_));
 sky130_fd_sc_hd__xnor2_1 _23313_ (.A(_14164_),
    .B(_09358_),
    .Y(\hash.CA1.p2[12] ));
 sky130_fd_sc_hd__inv_1 _23314_ (.A(_14161_),
    .Y(_09359_));
 sky130_fd_sc_hd__o21ai_4 _23315_ (.A1(_09351_),
    .A2(_09341_),
    .B1(_14162_),
    .Y(_09360_));
 sky130_fd_sc_hd__nand2_1 _23316_ (.A(_09359_),
    .B(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__a21o_1 _23317_ (.A1(_14164_),
    .A2(_09361_),
    .B1(_14163_),
    .X(_09362_));
 sky130_fd_sc_hd__xor2_1 _23318_ (.A(_14166_),
    .B(_09362_),
    .X(\hash.CA1.p2[13] ));
 sky130_fd_sc_hd__nor3_2 _23319_ (.A(_14161_),
    .B(_09357_),
    .C(_14163_),
    .Y(_09363_));
 sky130_fd_sc_hd__o21a_1 _23320_ (.A1(_14162_),
    .A2(_14161_),
    .B1(_14164_),
    .X(_09364_));
 sky130_fd_sc_hd__nor2_1 _23321_ (.A(_14163_),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__nor2_1 _23322_ (.A(_09363_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__a21oi_1 _23323_ (.A1(_14166_),
    .A2(_09366_),
    .B1(_14165_),
    .Y(_09367_));
 sky130_fd_sc_hd__xnor2_1 _23324_ (.A(_14168_),
    .B(_09367_),
    .Y(\hash.CA1.p2[14] ));
 sky130_fd_sc_hd__a21o_1 _23325_ (.A1(_14166_),
    .A2(_09362_),
    .B1(_14165_),
    .X(_09368_));
 sky130_fd_sc_hd__a21oi_1 _23326_ (.A1(_14168_),
    .A2(_09368_),
    .B1(_14167_),
    .Y(_09369_));
 sky130_fd_sc_hd__xnor2_1 _23327_ (.A(_14170_),
    .B(_09369_),
    .Y(\hash.CA1.p2[15] ));
 sky130_fd_sc_hd__nand3_1 _23328_ (.A(_14166_),
    .B(_14168_),
    .C(_14170_),
    .Y(_09370_));
 sky130_fd_sc_hd__or3_4 _23329_ (.A(_09363_),
    .B(_09365_),
    .C(_09370_),
    .X(_09371_));
 sky130_fd_sc_hd__a21o_1 _23330_ (.A1(_14168_),
    .A2(_14165_),
    .B1(_14167_),
    .X(_09372_));
 sky130_fd_sc_hd__a21oi_4 _23331_ (.A1(_14170_),
    .A2(_09372_),
    .B1(_14169_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand2_1 _23332_ (.A(_09371_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__xor2_1 _23333_ (.A(_14172_),
    .B(_09374_),
    .X(\hash.CA1.p2[16] ));
 sky130_fd_sc_hd__nand4_1 _23334_ (.A(_14164_),
    .B(_14166_),
    .C(_14168_),
    .D(_14170_),
    .Y(_09375_));
 sky130_fd_sc_hd__a21oi_4 _23335_ (.A1(_09360_),
    .A2(_09359_),
    .B1(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand4_1 _23336_ (.A(_14166_),
    .B(_14168_),
    .C(_14170_),
    .D(_14163_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand2_1 _23337_ (.A(_09373_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__o21a_1 _23338_ (.A1(_09376_),
    .A2(_09378_),
    .B1(_14172_),
    .X(_09379_));
 sky130_fd_sc_hd__nor2_1 _23339_ (.A(_14171_),
    .B(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__xnor2_1 _23340_ (.A(_14174_),
    .B(_09380_),
    .Y(\hash.CA1.p2[17] ));
 sky130_fd_sc_hd__nor2_1 _23341_ (.A(_14171_),
    .B(_14173_),
    .Y(_09381_));
 sky130_fd_sc_hd__o21a_1 _23342_ (.A1(_14172_),
    .A2(_14171_),
    .B1(_14174_),
    .X(_09382_));
 sky130_fd_sc_hd__nor2_1 _23343_ (.A(_14173_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__a31oi_4 _23344_ (.A1(_09371_),
    .A2(_09373_),
    .A3(_09381_),
    .B1(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__xor2_1 _23345_ (.A(_14176_),
    .B(_09384_),
    .X(\hash.CA1.p2[18] ));
 sky130_fd_sc_hd__o2111ai_2 _23346_ (.A1(_09378_),
    .A2(_09376_),
    .B1(_14172_),
    .C1(_14174_),
    .D1(_14176_),
    .Y(_09385_));
 sky130_fd_sc_hd__and3_1 _23347_ (.A(_14174_),
    .B(_14176_),
    .C(_14171_),
    .X(_09386_));
 sky130_fd_sc_hd__a21oi_1 _23348_ (.A1(_14176_),
    .A2(_14173_),
    .B1(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand3b_1 _23349_ (.A_N(_14175_),
    .B(_09385_),
    .C(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__xor2_1 _23350_ (.A(_14178_),
    .B(_09388_),
    .X(\hash.CA1.p2[19] ));
 sky130_fd_sc_hd__nand2_1 _23351_ (.A(_14180_),
    .B(_14177_),
    .Y(_09389_));
 sky130_fd_sc_hd__nand3_1 _23352_ (.A(_14178_),
    .B(_14180_),
    .C(_14175_),
    .Y(_09390_));
 sky130_fd_sc_hd__nand2_1 _23353_ (.A(_09389_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__a41o_4 _23354_ (.A1(_14176_),
    .A2(_14178_),
    .A3(_14180_),
    .A4(_09384_),
    .B1(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__a21o_1 _23355_ (.A1(_09384_),
    .A2(_14176_),
    .B1(_14175_),
    .X(_09393_));
 sky130_fd_sc_hd__a211oi_2 _23356_ (.A1(_09393_),
    .A2(_14178_),
    .B1(_14177_),
    .C1(_14180_),
    .Y(_09394_));
 sky130_fd_sc_hd__nor2_1 _23357_ (.A(_09392_),
    .B(_09394_),
    .Y(\hash.CA1.p2[20] ));
 sky130_fd_sc_hd__nor3_1 _23358_ (.A(_14175_),
    .B(_14177_),
    .C(_14179_),
    .Y(_09395_));
 sky130_fd_sc_hd__or2_0 _23359_ (.A(_14178_),
    .B(_14177_),
    .X(_09396_));
 sky130_fd_sc_hd__a21oi_2 _23360_ (.A1(_14180_),
    .A2(_09396_),
    .B1(_14179_),
    .Y(_09397_));
 sky130_fd_sc_hd__a31oi_2 _23361_ (.A1(_09395_),
    .A2(_09387_),
    .A3(_09385_),
    .B1(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__and2_4 _23362_ (.A(_09398_),
    .B(_14182_),
    .X(_09399_));
 sky130_fd_sc_hd__nor2_1 _23363_ (.A(_14182_),
    .B(_09398_),
    .Y(_09400_));
 sky130_fd_sc_hd__nor2_1 _23364_ (.A(_09399_),
    .B(_09400_),
    .Y(\hash.CA1.p2[21] ));
 sky130_fd_sc_hd__o21a_1 _23365_ (.A1(_14179_),
    .A2(_09392_),
    .B1(_14182_),
    .X(_09401_));
 sky130_fd_sc_hd__nor2_1 _23366_ (.A(_14181_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__xnor2_1 _23367_ (.A(_14184_),
    .B(_09402_),
    .Y(\hash.CA1.p2[22] ));
 sky130_fd_sc_hd__inv_1 _23368_ (.A(_14183_),
    .Y(_09403_));
 sky130_fd_sc_hd__o21ai_4 _23369_ (.A1(_14181_),
    .A2(_09399_),
    .B1(_14184_),
    .Y(_09404_));
 sky130_fd_sc_hd__clkinv_1 _23370_ (.A(_14186_),
    .Y(_09405_));
 sky130_fd_sc_hd__a21oi_4 _23371_ (.A1(_09404_),
    .A2(_09403_),
    .B1(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__and3_1 _23372_ (.A(_09405_),
    .B(_09403_),
    .C(_09404_),
    .X(_09407_));
 sky130_fd_sc_hd__nor2_1 _23373_ (.A(_09407_),
    .B(_09406_),
    .Y(\hash.CA1.p2[23] ));
 sky130_fd_sc_hd__inv_1 _23374_ (.A(_14184_),
    .Y(_09408_));
 sky130_fd_sc_hd__nor2_1 _23375_ (.A(_14182_),
    .B(_14181_),
    .Y(_09409_));
 sky130_fd_sc_hd__o21ai_0 _23376_ (.A1(_09408_),
    .A2(_09409_),
    .B1(_09403_),
    .Y(_09410_));
 sky130_fd_sc_hd__o41ai_4 _23377_ (.A1(_14179_),
    .A2(_14181_),
    .A3(_14183_),
    .A4(_09392_),
    .B1(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__o21bai_1 _23378_ (.A1(_09405_),
    .A2(_09411_),
    .B1_N(_14185_),
    .Y(_09412_));
 sky130_fd_sc_hd__xor2_1 _23379_ (.A(_14188_),
    .B(_09412_),
    .X(\hash.CA1.p2[24] ));
 sky130_fd_sc_hd__o21a_1 _23380_ (.A1(_14185_),
    .A2(_09406_),
    .B1(_14188_),
    .X(_09413_));
 sky130_fd_sc_hd__nor2_1 _23381_ (.A(_14187_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__xnor2_1 _23382_ (.A(_14190_),
    .B(_09414_),
    .Y(\hash.CA1.p2[25] ));
 sky130_fd_sc_hd__nand3_1 _23383_ (.A(_14186_),
    .B(_14188_),
    .C(_14190_),
    .Y(_09415_));
 sky130_fd_sc_hd__a21oi_2 _23384_ (.A1(_14188_),
    .A2(_14185_),
    .B1(_14187_),
    .Y(_09416_));
 sky130_fd_sc_hd__inv_2 _23385_ (.A(_14190_),
    .Y(_09417_));
 sky130_fd_sc_hd__o22ai_2 _23386_ (.A1(_09411_),
    .A2(_09415_),
    .B1(_09416_),
    .B2(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__nor2_2 _23387_ (.A(_14189_),
    .B(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__xnor2_2 _23388_ (.A(_14192_),
    .B(_09419_),
    .Y(\hash.CA1.p2[26] ));
 sky130_fd_sc_hd__nor2_1 _23389_ (.A(_14188_),
    .B(_14187_),
    .Y(_09420_));
 sky130_fd_sc_hd__o21bai_1 _23390_ (.A1(_09417_),
    .A2(_09420_),
    .B1_N(_14189_),
    .Y(_09421_));
 sky130_fd_sc_hd__o41a_1 _23391_ (.A1(_14185_),
    .A2(_14187_),
    .A3(_09406_),
    .A4(_14189_),
    .B1(_09421_),
    .X(_09422_));
 sky130_fd_sc_hd__a21oi_2 _23392_ (.A1(_09422_),
    .A2(_14192_),
    .B1(_14191_),
    .Y(_09423_));
 sky130_fd_sc_hd__xnor2_2 _23393_ (.A(_09423_),
    .B(_14194_),
    .Y(\hash.CA1.p2[27] ));
 sky130_fd_sc_hd__nor3_1 _23394_ (.A(_14192_),
    .B(_14191_),
    .C(_14193_),
    .Y(_09424_));
 sky130_fd_sc_hd__nor2_1 _23395_ (.A(_14194_),
    .B(_14193_),
    .Y(_09425_));
 sky130_fd_sc_hd__nor2_1 _23396_ (.A(_09424_),
    .B(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__o41ai_4 _23397_ (.A1(_14189_),
    .A2(_14191_),
    .A3(_14193_),
    .A4(_09418_),
    .B1(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__xnor2_1 _23398_ (.A(_09427_),
    .B(_14196_),
    .Y(\hash.CA1.p2[28] ));
 sky130_fd_sc_hd__inv_1 _23399_ (.A(_14196_),
    .Y(_09428_));
 sky130_fd_sc_hd__a21oi_1 _23400_ (.A1(_14194_),
    .A2(_14191_),
    .B1(_14193_),
    .Y(_09429_));
 sky130_fd_sc_hd__o21bai_1 _23401_ (.A1(_09428_),
    .A2(_09429_),
    .B1_N(_14195_),
    .Y(_09430_));
 sky130_fd_sc_hd__a41o_1 _23402_ (.A1(_09422_),
    .A2(_14194_),
    .A3(_14196_),
    .A4(_14192_),
    .B1(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__xor2_2 _23403_ (.A(_14198_),
    .B(_09431_),
    .X(\hash.CA1.p2[29] ));
 sky130_fd_sc_hd__o21bai_1 _23404_ (.A1(_09428_),
    .A2(_09427_),
    .B1_N(_14195_),
    .Y(_09432_));
 sky130_fd_sc_hd__a21oi_2 _23405_ (.A1(_09432_),
    .A2(_14198_),
    .B1(_14197_),
    .Y(_09433_));
 sky130_fd_sc_hd__xnor2_1 _23406_ (.A(_14201_),
    .B(_09433_),
    .Y(\hash.CA1.p2[30] ));
 sky130_fd_sc_hd__xnor2_1 _23407_ (.A(\hash.CA2.f_dash[31] ),
    .B(_08094_),
    .Y(_09434_));
 sky130_fd_sc_hd__nor2_1 _23408_ (.A(net353),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__xor2_4 _23409_ (.A(\hash.CA1.w_i1[31] ),
    .B(\hash.CA1.k_i1[31] ),
    .X(_09436_));
 sky130_fd_sc_hd__xnor2_1 _23410_ (.A(_09435_),
    .B(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__xnor2_1 _23411_ (.A(\hash.CA1.S1.X[10] ),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__xnor2_1 _23412_ (.A(_06673_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__nand2_1 _23413_ (.A(_14115_),
    .B(_14124_),
    .Y(_09440_));
 sky130_fd_sc_hd__a21oi_1 _23414_ (.A1(_14124_),
    .A2(_14114_),
    .B1(_14123_),
    .Y(_09441_));
 sky130_fd_sc_hd__o21ai_0 _23415_ (.A1(_07134_),
    .A2(_09440_),
    .B1(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__xnor2_1 _23416_ (.A(_09439_),
    .B(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__nor2b_1 _23417_ (.A(_07108_),
    .B_N(_14120_),
    .Y(_09444_));
 sky130_fd_sc_hd__a311oi_1 _23418_ (.A1(_14111_),
    .A2(_14120_),
    .A3(_08101_),
    .B1(_09444_),
    .C1(_14119_),
    .Y(_09445_));
 sky130_fd_sc_hd__xnor2_1 _23419_ (.A(_09443_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__nor2b_2 _23420_ (.A(net352),
    .B_N(\hash.CA2.S1.X[31] ),
    .Y(_09447_));
 sky130_fd_sc_hd__mux2i_4 _23421_ (.A0(_09447_),
    .A1(_06418_),
    .S(net1069),
    .Y(_09448_));
 sky130_fd_sc_hd__xnor2_2 _23422_ (.A(_09446_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__xor2_1 _23423_ (.A(_12877_),
    .B(_12873_),
    .X(_09450_));
 sky130_fd_sc_hd__nor2_1 _23424_ (.A(net353),
    .B(\hash.CA2.b_dash[31] ),
    .Y(_09451_));
 sky130_fd_sc_hd__xnor2_1 _23425_ (.A(_09450_),
    .B(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__nand3_1 _23426_ (.A(_14192_),
    .B(_14194_),
    .C(_14196_),
    .Y(_09453_));
 sky130_fd_sc_hd__nand4_1 _23427_ (.A(_14188_),
    .B(_14190_),
    .C(_14198_),
    .D(_14201_),
    .Y(_09454_));
 sky130_fd_sc_hd__nor2_1 _23428_ (.A(_09453_),
    .B(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__nor2_1 _23429_ (.A(_09417_),
    .B(_09416_),
    .Y(_09456_));
 sky130_fd_sc_hd__o21ai_0 _23430_ (.A1(_14189_),
    .A2(_09456_),
    .B1(_14192_),
    .Y(_09457_));
 sky130_fd_sc_hd__nand2b_1 _23431_ (.A_N(_14191_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__a21oi_1 _23432_ (.A1(_14194_),
    .A2(_09458_),
    .B1(_14193_),
    .Y(_09459_));
 sky130_fd_sc_hd__o21bai_1 _23433_ (.A1(_09428_),
    .A2(_09459_),
    .B1_N(_14195_),
    .Y(_09460_));
 sky130_fd_sc_hd__a21oi_1 _23434_ (.A1(_14198_),
    .A2(_09460_),
    .B1(_14197_),
    .Y(_09461_));
 sky130_fd_sc_hd__nor2b_1 _23435_ (.A(_09461_),
    .B_N(_14201_),
    .Y(_09462_));
 sky130_fd_sc_hd__a211oi_2 _23436_ (.A1(_09406_),
    .A2(_09455_),
    .B1(_09462_),
    .C1(_14200_),
    .Y(_09463_));
 sky130_fd_sc_hd__xnor2_1 _23437_ (.A(_09452_),
    .B(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__xnor2_1 _23438_ (.A(_09449_),
    .B(_09464_),
    .Y(\hash.CA1.p2[31] ));
 sky130_fd_sc_hd__xnor2_1 _23439_ (.A(_12885_),
    .B(_14135_),
    .Y(\hash.CA1.p2[3] ));
 sky130_fd_sc_hd__xor2_1 _23440_ (.A(_14139_),
    .B(_09332_),
    .X(\hash.CA1.p2[4] ));
 sky130_fd_sc_hd__nor2_1 _23441_ (.A(_14138_),
    .B(_09343_),
    .Y(_09465_));
 sky130_fd_sc_hd__xnor2_1 _23442_ (.A(_14143_),
    .B(_09465_),
    .Y(\hash.CA1.p2[5] ));
 sky130_fd_sc_hd__xnor2_2 _23443_ (.A(_14147_),
    .B(_09335_),
    .Y(\hash.CA1.p2[6] ));
 sky130_fd_sc_hd__nand2b_1 _23444_ (.A_N(_14142_),
    .B(_09344_),
    .Y(_09466_));
 sky130_fd_sc_hd__a21oi_2 _23445_ (.A1(_14147_),
    .A2(_09466_),
    .B1(_14146_),
    .Y(_09467_));
 sky130_fd_sc_hd__xnor2_2 _23446_ (.A(_14151_),
    .B(_09467_),
    .Y(\hash.CA1.p2[7] ));
 sky130_fd_sc_hd__xnor2_2 _23447_ (.A(_14155_),
    .B(_09337_),
    .Y(\hash.CA1.p2[8] ));
 sky130_fd_sc_hd__o21bai_1 _23448_ (.A1(_09346_),
    .A2(_09467_),
    .B1_N(_14150_),
    .Y(_09468_));
 sky130_fd_sc_hd__a21oi_2 _23449_ (.A1(_14155_),
    .A2(_09468_),
    .B1(_14154_),
    .Y(_09469_));
 sky130_fd_sc_hd__xnor2_2 _23450_ (.A(_14158_),
    .B(_09469_),
    .Y(\hash.CA1.p2[9] ));
 sky130_fd_sc_hd__inv_2 _23451_ (.A(_13918_),
    .Y(_09470_));
 sky130_fd_sc_hd__inv_1 _23452_ (.A(_13893_),
    .Y(_09471_));
 sky130_fd_sc_hd__a21o_4 _23453_ (.A1(_14208_),
    .A2(_13874_),
    .B1(_13873_),
    .X(_09472_));
 sky130_fd_sc_hd__a21oi_4 _23454_ (.A1(_13883_),
    .A2(_09472_),
    .B1(_13882_),
    .Y(_09473_));
 sky130_fd_sc_hd__inv_2 _23455_ (.A(_13892_),
    .Y(_09474_));
 sky130_fd_sc_hd__o21ai_1 _23456_ (.A1(_09471_),
    .A2(_09473_),
    .B1(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__a21o_4 _23457_ (.A1(_13902_),
    .A2(_09475_),
    .B1(_13901_),
    .X(_09476_));
 sky130_fd_sc_hd__a21oi_2 _23458_ (.A1(_13910_),
    .A2(_09476_),
    .B1(_13909_),
    .Y(_09477_));
 sky130_fd_sc_hd__nor2_1 _23459_ (.A(_09470_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__o21ai_0 _23460_ (.A1(_13917_),
    .A2(_09478_),
    .B1(_13927_),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2b_1 _23461_ (.A_N(_13926_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__a21oi_2 _23462_ (.A1(_13936_),
    .A2(_09480_),
    .B1(_13935_),
    .Y(_09481_));
 sky130_fd_sc_hd__xnor2_4 _23463_ (.A(_13945_),
    .B(_09481_),
    .Y(\hash.CA1.p3[10] ));
 sky130_fd_sc_hd__nor2b_1 _23464_ (.A(_12892_),
    .B_N(_13883_),
    .Y(_09482_));
 sky130_fd_sc_hd__o21ai_2 _23465_ (.A1(_13882_),
    .A2(_09482_),
    .B1(_13893_),
    .Y(_09483_));
 sky130_fd_sc_hd__a21boi_4 _23466_ (.A1(_09474_),
    .A2(_09483_),
    .B1_N(_13902_),
    .Y(_09484_));
 sky130_fd_sc_hd__nor2_2 _23467_ (.A(_13901_),
    .B(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__nand2_1 _23468_ (.A(_13910_),
    .B(_13918_),
    .Y(_09486_));
 sky130_fd_sc_hd__a21oi_1 _23469_ (.A1(_13918_),
    .A2(_13909_),
    .B1(_13917_),
    .Y(_09487_));
 sky130_fd_sc_hd__o21ai_2 _23470_ (.A1(_09485_),
    .A2(_09486_),
    .B1(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__and2_4 _23471_ (.A(_13927_),
    .B(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__o21a_4 _23472_ (.A1(_13926_),
    .A2(_09489_),
    .B1(_13936_),
    .X(_09490_));
 sky130_fd_sc_hd__o21a_4 _23473_ (.A1(_13935_),
    .A2(_09490_),
    .B1(_13945_),
    .X(_09491_));
 sky130_fd_sc_hd__nor2_4 _23474_ (.A(_13944_),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__xnor2_4 _23475_ (.A(_13955_),
    .B(_09492_),
    .Y(\hash.CA1.p3[11] ));
 sky130_fd_sc_hd__nand4_1 _23476_ (.A(_13945_),
    .B(_13955_),
    .C(_13927_),
    .D(_13936_),
    .Y(_09493_));
 sky130_fd_sc_hd__inv_1 _23477_ (.A(_13955_),
    .Y(_09494_));
 sky130_fd_sc_hd__a21o_1 _23478_ (.A1(_13936_),
    .A2(_13926_),
    .B1(_13935_),
    .X(_09495_));
 sky130_fd_sc_hd__a21oi_2 _23479_ (.A1(_13945_),
    .A2(_09495_),
    .B1(_13944_),
    .Y(_09496_));
 sky130_fd_sc_hd__nor2_2 _23480_ (.A(_09494_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__inv_1 _23481_ (.A(_13917_),
    .Y(_09498_));
 sky130_fd_sc_hd__nor2_1 _23482_ (.A(_09498_),
    .B(_09493_),
    .Y(_09499_));
 sky130_fd_sc_hd__nor2_2 _23483_ (.A(_09499_),
    .B(_09497_),
    .Y(_09500_));
 sky130_fd_sc_hd__o31ai_4 _23484_ (.A1(_09470_),
    .A2(_09477_),
    .A3(_09493_),
    .B1(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__nor2_1 _23485_ (.A(_13954_),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__xnor2_2 _23486_ (.A(_13964_),
    .B(_09502_),
    .Y(\hash.CA1.p3[12] ));
 sky130_fd_sc_hd__o21bai_1 _23487_ (.A1(_09494_),
    .A2(_09492_),
    .B1_N(_13954_),
    .Y(_09503_));
 sky130_fd_sc_hd__a21oi_1 _23488_ (.A1(_13964_),
    .A2(_09503_),
    .B1(_13963_),
    .Y(_09504_));
 sky130_fd_sc_hd__xnor2_2 _23489_ (.A(_13972_),
    .B(_09504_),
    .Y(\hash.CA1.p3[13] ));
 sky130_fd_sc_hd__o21ai_0 _23490_ (.A1(_13954_),
    .A2(_09501_),
    .B1(_13964_),
    .Y(_09505_));
 sky130_fd_sc_hd__nand2b_1 _23491_ (.A_N(_13963_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__a21oi_1 _23492_ (.A1(_13972_),
    .A2(_09506_),
    .B1(_13971_),
    .Y(_09507_));
 sky130_fd_sc_hd__xnor2_1 _23493_ (.A(_13981_),
    .B(_09507_),
    .Y(\hash.CA1.p3[14] ));
 sky130_fd_sc_hd__o211ai_1 _23494_ (.A1(_13963_),
    .A2(_13964_),
    .B1(_13972_),
    .C1(_13981_),
    .Y(_09508_));
 sky130_fd_sc_hd__nor3_2 _23495_ (.A(_13954_),
    .B(_13963_),
    .C(_09497_),
    .Y(_09509_));
 sky130_fd_sc_hd__a21oi_2 _23496_ (.A1(_13981_),
    .A2(_13971_),
    .B1(_13980_),
    .Y(_09510_));
 sky130_fd_sc_hd__o21ai_2 _23497_ (.A1(_09508_),
    .A2(_09509_),
    .B1(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__nor3b_2 _23498_ (.A(_09493_),
    .B(_09508_),
    .C_N(_09488_),
    .Y(_09512_));
 sky130_fd_sc_hd__o21a_4 _23499_ (.A1(_09511_),
    .A2(_09512_),
    .B1(_13991_),
    .X(_09513_));
 sky130_fd_sc_hd__nor3_2 _23500_ (.A(_13991_),
    .B(_09511_),
    .C(_09512_),
    .Y(_09514_));
 sky130_fd_sc_hd__nor2_4 _23501_ (.A(_09513_),
    .B(_09514_),
    .Y(\hash.CA1.p3[15] ));
 sky130_fd_sc_hd__nor3_1 _23502_ (.A(_13954_),
    .B(_13963_),
    .C(_13990_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand2_1 _23503_ (.A(_09510_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__a21boi_1 _23504_ (.A1(_09510_),
    .A2(_09508_),
    .B1_N(_13991_),
    .Y(_09517_));
 sky130_fd_sc_hd__o22ai_1 _23505_ (.A1(_09501_),
    .A2(_09516_),
    .B1(_09517_),
    .B2(_13990_),
    .Y(_09518_));
 sky130_fd_sc_hd__xnor2_1 _23506_ (.A(_14000_),
    .B(_09518_),
    .Y(\hash.CA1.p3[16] ));
 sky130_fd_sc_hd__o21a_1 _23507_ (.A1(_14000_),
    .A2(_13999_),
    .B1(_14008_),
    .X(_09519_));
 sky130_fd_sc_hd__o31a_1 _23508_ (.A1(_13990_),
    .A2(_13999_),
    .A3(_09513_),
    .B1(_09519_),
    .X(_09520_));
 sky130_fd_sc_hd__o21ai_0 _23509_ (.A1(_13990_),
    .A2(_09513_),
    .B1(_14000_),
    .Y(_09521_));
 sky130_fd_sc_hd__nor3b_1 _23510_ (.A(_14008_),
    .B(_13999_),
    .C_N(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__nor2_1 _23511_ (.A(_09520_),
    .B(_09522_),
    .Y(\hash.CA1.p3[17] ));
 sky130_fd_sc_hd__o221a_4 _23512_ (.A1(_09516_),
    .A2(_09501_),
    .B1(_09517_),
    .B2(_13990_),
    .C1(_14000_),
    .X(_09523_));
 sky130_fd_sc_hd__o21a_1 _23513_ (.A1(_13999_),
    .A2(_09523_),
    .B1(_14008_),
    .X(_09524_));
 sky130_fd_sc_hd__nor2_1 _23514_ (.A(_14007_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__xnor2_1 _23515_ (.A(_14016_),
    .B(_09525_),
    .Y(\hash.CA1.p3[18] ));
 sky130_fd_sc_hd__o21a_1 _23516_ (.A1(_14007_),
    .A2(_09520_),
    .B1(_14016_),
    .X(_09526_));
 sky130_fd_sc_hd__nor2_1 _23517_ (.A(_14015_),
    .B(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__xnor2_1 _23518_ (.A(_14024_),
    .B(_09527_),
    .Y(\hash.CA1.p3[19] ));
 sky130_fd_sc_hd__o21a_1 _23519_ (.A1(_14008_),
    .A2(_14007_),
    .B1(_14016_),
    .X(_09528_));
 sky130_fd_sc_hd__o31ai_4 _23520_ (.A1(_09523_),
    .A2(_14007_),
    .A3(_13999_),
    .B1(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__nand2b_1 _23521_ (.A_N(_14015_),
    .B(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__a21oi_1 _23522_ (.A1(_14024_),
    .A2(_09530_),
    .B1(_14023_),
    .Y(_09531_));
 sky130_fd_sc_hd__xnor2_1 _23523_ (.A(_14032_),
    .B(_09531_),
    .Y(\hash.CA1.p3[20] ));
 sky130_fd_sc_hd__or3_4 _23524_ (.A(_14007_),
    .B(_14015_),
    .C(_14023_),
    .X(_09532_));
 sky130_fd_sc_hd__or2_0 _23525_ (.A(_09520_),
    .B(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__or3_4 _23526_ (.A(_14016_),
    .B(_14015_),
    .C(_14023_),
    .X(_09534_));
 sky130_fd_sc_hd__or2_4 _23527_ (.A(_14024_),
    .B(_14023_),
    .X(_09535_));
 sky130_fd_sc_hd__a41o_1 _23528_ (.A1(_14032_),
    .A2(_09533_),
    .A3(_09534_),
    .A4(_09535_),
    .B1(_14031_),
    .X(_09536_));
 sky130_fd_sc_hd__xor2_1 _23529_ (.A(_14041_),
    .B(_09536_),
    .X(\hash.CA1.p3[21] ));
 sky130_fd_sc_hd__nor3_1 _23530_ (.A(_14015_),
    .B(_14023_),
    .C(_14031_),
    .Y(_09537_));
 sky130_fd_sc_hd__a21oi_1 _23531_ (.A1(_14032_),
    .A2(_09535_),
    .B1(_14031_),
    .Y(_09538_));
 sky130_fd_sc_hd__a21oi_2 _23532_ (.A1(_09537_),
    .A2(_09529_),
    .B1(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__a21oi_1 _23533_ (.A1(_14041_),
    .A2(_09539_),
    .B1(_14040_),
    .Y(_09540_));
 sky130_fd_sc_hd__xnor2_1 _23534_ (.A(_14051_),
    .B(_09540_),
    .Y(\hash.CA1.p3[22] ));
 sky130_fd_sc_hd__and3_1 _23535_ (.A(_14032_),
    .B(_14041_),
    .C(_14051_),
    .X(_09541_));
 sky130_fd_sc_hd__o2111ai_2 _23536_ (.A1(_09520_),
    .A2(_09532_),
    .B1(_09534_),
    .C1(_09535_),
    .D1(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__and3_1 _23537_ (.A(_14041_),
    .B(_14051_),
    .C(_14031_),
    .X(_09543_));
 sky130_fd_sc_hd__a21oi_1 _23538_ (.A1(_14051_),
    .A2(_14040_),
    .B1(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nand3b_1 _23539_ (.A_N(_14050_),
    .B(_09542_),
    .C(_09544_),
    .Y(_09545_));
 sky130_fd_sc_hd__xor2_1 _23540_ (.A(_14061_),
    .B(_09545_),
    .X(\hash.CA1.p3[23] ));
 sky130_fd_sc_hd__nand2_1 _23541_ (.A(_14061_),
    .B(_14050_),
    .Y(_09546_));
 sky130_fd_sc_hd__nand3_1 _23542_ (.A(_14051_),
    .B(_14061_),
    .C(_14040_),
    .Y(_09547_));
 sky130_fd_sc_hd__nand2_1 _23543_ (.A(_09546_),
    .B(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__a41oi_2 _23544_ (.A1(_09539_),
    .A2(_14051_),
    .A3(_14061_),
    .A4(_14041_),
    .B1(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__nor2b_2 _23545_ (.A(_14060_),
    .B_N(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__xnor2_1 _23546_ (.A(_14071_),
    .B(_09550_),
    .Y(\hash.CA1.p3[24] ));
 sky130_fd_sc_hd__nor3_1 _23547_ (.A(_14050_),
    .B(_14060_),
    .C(_14070_),
    .Y(_09551_));
 sky130_fd_sc_hd__or2_4 _23548_ (.A(_14071_),
    .B(_14070_),
    .X(_09552_));
 sky130_fd_sc_hd__o31ai_1 _23549_ (.A1(_14061_),
    .A2(_14060_),
    .A3(_14070_),
    .B1(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__a31o_4 _23550_ (.A1(_09542_),
    .A2(_09544_),
    .A3(_09551_),
    .B1(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__xnor2_1 _23551_ (.A(_14081_),
    .B(_09554_),
    .Y(\hash.CA1.p3[25] ));
 sky130_fd_sc_hd__nor3_1 _23552_ (.A(_14060_),
    .B(_14070_),
    .C(_14080_),
    .Y(_09555_));
 sky130_fd_sc_hd__a21oi_1 _23553_ (.A1(_14081_),
    .A2(_09552_),
    .B1(_14080_),
    .Y(_09556_));
 sky130_fd_sc_hd__a21oi_2 _23554_ (.A1(_09555_),
    .A2(_09549_),
    .B1(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__xor2_1 _23555_ (.A(_14090_),
    .B(_09557_),
    .X(\hash.CA1.p3[26] ));
 sky130_fd_sc_hd__nand2_1 _23556_ (.A(_14081_),
    .B(_14090_),
    .Y(_09558_));
 sky130_fd_sc_hd__a21oi_1 _23557_ (.A1(_14090_),
    .A2(_14080_),
    .B1(_14089_),
    .Y(_09559_));
 sky130_fd_sc_hd__o21ai_4 _23558_ (.A1(_09554_),
    .A2(_09558_),
    .B1(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__xor2_1 _23559_ (.A(_14099_),
    .B(_09560_),
    .X(\hash.CA1.p3[27] ));
 sky130_fd_sc_hd__a21o_1 _23560_ (.A1(_09557_),
    .A2(_14090_),
    .B1(_14089_),
    .X(_09561_));
 sky130_fd_sc_hd__a21oi_2 _23561_ (.A1(_09561_),
    .A2(_14099_),
    .B1(_14098_),
    .Y(_09562_));
 sky130_fd_sc_hd__xnor2_1 _23562_ (.A(_09562_),
    .B(_14109_),
    .Y(\hash.CA1.p3[28] ));
 sky130_fd_sc_hd__a21o_1 _23563_ (.A1(_14099_),
    .A2(_09560_),
    .B1(_14098_),
    .X(_09563_));
 sky130_fd_sc_hd__a21oi_2 _23564_ (.A1(_09563_),
    .A2(_14109_),
    .B1(_14108_),
    .Y(_09564_));
 sky130_fd_sc_hd__xnor2_1 _23565_ (.A(_14118_),
    .B(_09564_),
    .Y(\hash.CA1.p3[29] ));
 sky130_fd_sc_hd__nand2_1 _23566_ (.A(_09557_),
    .B(_14090_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand3_1 _23567_ (.A(_14099_),
    .B(_14109_),
    .C(_14118_),
    .Y(_09566_));
 sky130_fd_sc_hd__a21o_1 _23568_ (.A1(_14099_),
    .A2(_14089_),
    .B1(_14098_),
    .X(_09567_));
 sky130_fd_sc_hd__a21o_1 _23569_ (.A1(_14109_),
    .A2(_09567_),
    .B1(_14108_),
    .X(_09568_));
 sky130_fd_sc_hd__a21oi_1 _23570_ (.A1(_14118_),
    .A2(_09568_),
    .B1(_14117_),
    .Y(_09569_));
 sky130_fd_sc_hd__o21ai_1 _23571_ (.A1(_09566_),
    .A2(_09565_),
    .B1(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__xor2_1 _23572_ (.A(_14127_),
    .B(_09570_),
    .X(\hash.CA1.p3[30] ));
 sky130_fd_sc_hd__nor3b_1 _23573_ (.A(_09566_),
    .B(_12651_),
    .C_N(_14127_),
    .Y(_09571_));
 sky130_fd_sc_hd__a21o_1 _23574_ (.A1(_14109_),
    .A2(_14098_),
    .B1(_14108_),
    .X(_09572_));
 sky130_fd_sc_hd__a21o_1 _23575_ (.A1(_14118_),
    .A2(_09572_),
    .B1(_14117_),
    .X(_09573_));
 sky130_fd_sc_hd__nor4b_1 _23576_ (.A(_14126_),
    .B(_09560_),
    .C(_09573_),
    .D_N(_12651_),
    .Y(_09574_));
 sky130_fd_sc_hd__a21oi_1 _23577_ (.A1(_14127_),
    .A2(_09573_),
    .B1(_14126_),
    .Y(_09575_));
 sky130_fd_sc_hd__nand2b_1 _23578_ (.A_N(_09573_),
    .B(_09566_),
    .Y(_09576_));
 sky130_fd_sc_hd__a21oi_1 _23579_ (.A1(_14127_),
    .A2(_09576_),
    .B1(_14126_),
    .Y(_09577_));
 sky130_fd_sc_hd__nand2_1 _23580_ (.A(_12651_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__o21ai_0 _23581_ (.A1(_12651_),
    .A2(_09575_),
    .B1(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__a211o_1 _23582_ (.A1(net1075),
    .A2(_09571_),
    .B1(_09574_),
    .C1(_09579_),
    .X(_09580_));
 sky130_fd_sc_hd__xnor2_2 _23583_ (.A(_09449_),
    .B(_09580_),
    .Y(\hash.CA1.p3[31] ));
 sky130_fd_sc_hd__xnor2_2 _23584_ (.A(_12892_),
    .B(_13883_),
    .Y(\hash.CA1.p3[3] ));
 sky130_fd_sc_hd__xnor2_4 _23585_ (.A(_13893_),
    .B(_09473_),
    .Y(\hash.CA1.p3[4] ));
 sky130_fd_sc_hd__nand2_1 _23586_ (.A(_09474_),
    .B(_09483_),
    .Y(_09581_));
 sky130_fd_sc_hd__nor2_1 _23587_ (.A(_13902_),
    .B(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__nor2_4 _23588_ (.A(_09484_),
    .B(_09582_),
    .Y(\hash.CA1.p3[5] ));
 sky130_fd_sc_hd__xor2_4 _23589_ (.A(_13910_),
    .B(_09476_),
    .X(\hash.CA1.p3[6] ));
 sky130_fd_sc_hd__inv_1 _23590_ (.A(_09485_),
    .Y(_09583_));
 sky130_fd_sc_hd__a21oi_1 _23591_ (.A1(_13910_),
    .A2(_09583_),
    .B1(_13909_),
    .Y(_09584_));
 sky130_fd_sc_hd__xnor2_2 _23592_ (.A(_13918_),
    .B(_09584_),
    .Y(\hash.CA1.p3[7] ));
 sky130_fd_sc_hd__nor2_2 _23593_ (.A(_13917_),
    .B(_09478_),
    .Y(_09585_));
 sky130_fd_sc_hd__xnor2_4 _23594_ (.A(_13927_),
    .B(_09585_),
    .Y(\hash.CA1.p3[8] ));
 sky130_fd_sc_hd__nor3_2 _23595_ (.A(_13936_),
    .B(_13926_),
    .C(_09489_),
    .Y(_09586_));
 sky130_fd_sc_hd__nor2_4 _23596_ (.A(_09490_),
    .B(_09586_),
    .Y(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__xor2_1 _23597_ (.A(\hash.CA1.k_i2[31] ),
    .B(_12495_),
    .X(_09587_));
 sky130_fd_sc_hd__xnor2_1 _23598_ (.A(_06418_),
    .B(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__xnor2_1 _23599_ (.A(\hash.CA1.w_i2[31] ),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__o21bai_1 _23600_ (.A1(_08034_),
    .A2(_08038_),
    .B1_N(_13825_),
    .Y(_09590_));
 sky130_fd_sc_hd__a21o_1 _23601_ (.A1(_13833_),
    .A2(_09590_),
    .B1(_13832_),
    .X(_09591_));
 sky130_fd_sc_hd__a21oi_1 _23602_ (.A1(_13839_),
    .A2(_09591_),
    .B1(_13838_),
    .Y(_09592_));
 sky130_fd_sc_hd__o21ai_0 _23603_ (.A1(_08035_),
    .A2(_08051_),
    .B1(_09592_),
    .Y(_09593_));
 sky130_fd_sc_hd__a21oi_2 _23604_ (.A1(_13844_),
    .A2(_09593_),
    .B1(_13843_),
    .Y(_09594_));
 sky130_fd_sc_hd__xnor2_4 _23605_ (.A(_09589_),
    .B(_09594_),
    .Y(\hash.CA1.p4[31] ));
 sky130_fd_sc_hd__clkinv_1 _23606_ (.A(_13723_),
    .Y(_09595_));
 sky130_fd_sc_hd__a21o_4 _23607_ (.A1(_13712_),
    .A2(_13704_),
    .B1(_13711_),
    .X(_09596_));
 sky130_fd_sc_hd__a21oi_4 _23608_ (.A1(_13718_),
    .A2(_09596_),
    .B1(_13717_),
    .Y(_09597_));
 sky130_fd_sc_hd__clkinv_1 _23609_ (.A(_13698_),
    .Y(_09598_));
 sky130_fd_sc_hd__clkinv_1 _23610_ (.A(_13680_),
    .Y(_09599_));
 sky130_fd_sc_hd__nor2b_1 _23611_ (.A(_12896_),
    .B_N(_13675_),
    .Y(_09600_));
 sky130_fd_sc_hd__o21ai_1 _23612_ (.A1(_13674_),
    .A2(_09600_),
    .B1(_13681_),
    .Y(_09601_));
 sky130_fd_sc_hd__a21boi_2 _23613_ (.A1(_09599_),
    .A2(_09601_),
    .B1_N(_13687_),
    .Y(_09602_));
 sky130_fd_sc_hd__o21a_4 _23614_ (.A1(_13686_),
    .A2(_09602_),
    .B1(_13693_),
    .X(_09603_));
 sky130_fd_sc_hd__o21ai_2 _23615_ (.A1(_13692_),
    .A2(_09603_),
    .B1(_13699_),
    .Y(_09604_));
 sky130_fd_sc_hd__and3_4 _23616_ (.A(_13705_),
    .B(_13712_),
    .C(_13718_),
    .X(_09605_));
 sky130_fd_sc_hd__a21bo_4 _23617_ (.A1(_09598_),
    .A2(_09604_),
    .B1_N(_09605_),
    .X(_09606_));
 sky130_fd_sc_hd__nand2_1 _23618_ (.A(_09597_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__xnor2_1 _23619_ (.A(_09595_),
    .B(_09607_),
    .Y(\hash.CA1.p5[10] ));
 sky130_fd_sc_hd__inv_1 _23620_ (.A(_13681_),
    .Y(_09608_));
 sky130_fd_sc_hd__a21o_1 _23621_ (.A1(_12898_),
    .A2(_13670_),
    .B1(_13669_),
    .X(_09609_));
 sky130_fd_sc_hd__a21oi_2 _23622_ (.A1(_13675_),
    .A2(_09609_),
    .B1(_13674_),
    .Y(_09610_));
 sky130_fd_sc_hd__o21ai_2 _23623_ (.A1(_09608_),
    .A2(_09610_),
    .B1(_09599_),
    .Y(_09611_));
 sky130_fd_sc_hd__a21oi_4 _23624_ (.A1(_13687_),
    .A2(_09611_),
    .B1(_13686_),
    .Y(_09612_));
 sky130_fd_sc_hd__nor2_2 _23625_ (.A(_13692_),
    .B(_13698_),
    .Y(_09613_));
 sky130_fd_sc_hd__nand3_1 _23626_ (.A(_13723_),
    .B(_13729_),
    .C(_09605_),
    .Y(_09614_));
 sky130_fd_sc_hd__o21a_1 _23627_ (.A1(_13693_),
    .A2(_13692_),
    .B1(_13699_),
    .X(_09615_));
 sky130_fd_sc_hd__nor2_2 _23628_ (.A(_13698_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__a211oi_2 _23629_ (.A1(_09612_),
    .A2(_09613_),
    .B1(_09614_),
    .C1(_09616_),
    .Y(_09617_));
 sky130_fd_sc_hd__nand2_1 _23630_ (.A(_13723_),
    .B(_13729_),
    .Y(_09618_));
 sky130_fd_sc_hd__nand2_1 _23631_ (.A(_13729_),
    .B(_13722_),
    .Y(_09619_));
 sky130_fd_sc_hd__o21ai_2 _23632_ (.A1(_09597_),
    .A2(_09618_),
    .B1(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__a21oi_2 _23633_ (.A1(_09612_),
    .A2(_09613_),
    .B1(_09616_),
    .Y(_09621_));
 sky130_fd_sc_hd__nand2_1 _23634_ (.A(_09605_),
    .B(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__nand2_1 _23635_ (.A(_09597_),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__a211oi_1 _23636_ (.A1(_13723_),
    .A2(_09623_),
    .B1(_13722_),
    .C1(_13729_),
    .Y(_09624_));
 sky130_fd_sc_hd__nor3_1 _23637_ (.A(_09617_),
    .B(_09620_),
    .C(_09624_),
    .Y(\hash.CA1.p5[11] ));
 sky130_fd_sc_hd__a21o_1 _23638_ (.A1(_13723_),
    .A2(_09607_),
    .B1(_13722_),
    .X(_09625_));
 sky130_fd_sc_hd__a21oi_1 _23639_ (.A1(_13729_),
    .A2(_09625_),
    .B1(_13728_),
    .Y(_09626_));
 sky130_fd_sc_hd__xnor2_1 _23640_ (.A(_13736_),
    .B(_09626_),
    .Y(\hash.CA1.p5[12] ));
 sky130_fd_sc_hd__o31ai_1 _23641_ (.A1(_13728_),
    .A2(_09617_),
    .A3(_09620_),
    .B1(_13736_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand2b_1 _23642_ (.A_N(_13735_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__xor2_1 _23643_ (.A(_13742_),
    .B(_09628_),
    .X(\hash.CA1.p5[13] ));
 sky130_fd_sc_hd__nand2_1 _23644_ (.A(_13729_),
    .B(_13736_),
    .Y(_09629_));
 sky130_fd_sc_hd__a211oi_2 _23645_ (.A1(_09597_),
    .A2(_09606_),
    .B1(_09629_),
    .C1(_09595_),
    .Y(_09630_));
 sky130_fd_sc_hd__nand2b_1 _23646_ (.A_N(_13728_),
    .B(_09619_),
    .Y(_09631_));
 sky130_fd_sc_hd__a21o_4 _23647_ (.A1(_13736_),
    .A2(_09631_),
    .B1(_13735_),
    .X(_09632_));
 sky130_fd_sc_hd__o21ai_2 _23648_ (.A1(_09630_),
    .A2(_09632_),
    .B1(_13742_),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2b_4 _23649_ (.A_N(_13741_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__xor2_1 _23650_ (.A(_13748_),
    .B(_09634_),
    .X(\hash.CA1.p5[14] ));
 sky130_fd_sc_hd__or3_1 _23651_ (.A(_13728_),
    .B(_13735_),
    .C(_13741_),
    .X(_09635_));
 sky130_fd_sc_hd__nor3_1 _23652_ (.A(_13736_),
    .B(_13735_),
    .C(_13741_),
    .Y(_09636_));
 sky130_fd_sc_hd__nor2_1 _23653_ (.A(_13742_),
    .B(_13741_),
    .Y(_09637_));
 sky130_fd_sc_hd__nor2_1 _23654_ (.A(_09636_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__o31ai_2 _23655_ (.A1(_09617_),
    .A2(_09620_),
    .A3(_09635_),
    .B1(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__nor2b_1 _23656_ (.A(_09639_),
    .B_N(_13748_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2_1 _23657_ (.A(_13747_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__xnor2_1 _23658_ (.A(_13755_),
    .B(_09641_),
    .Y(\hash.CA1.p5[15] ));
 sky130_fd_sc_hd__a21o_1 _23659_ (.A1(_13748_),
    .A2(_09634_),
    .B1(_13747_),
    .X(_09642_));
 sky130_fd_sc_hd__a21o_1 _23660_ (.A1(_13755_),
    .A2(_09642_),
    .B1(_13754_),
    .X(_09643_));
 sky130_fd_sc_hd__xor2_1 _23661_ (.A(_13762_),
    .B(_09643_),
    .X(\hash.CA1.p5[16] ));
 sky130_fd_sc_hd__o21ai_0 _23662_ (.A1(_13747_),
    .A2(_09640_),
    .B1(_13755_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand2b_1 _23663_ (.A_N(_13754_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__a21oi_1 _23664_ (.A1(_13762_),
    .A2(_09645_),
    .B1(_13761_),
    .Y(_09646_));
 sky130_fd_sc_hd__xnor2_1 _23665_ (.A(_13769_),
    .B(_09646_),
    .Y(\hash.CA1.p5[17] ));
 sky130_fd_sc_hd__and2_0 _23666_ (.A(_13762_),
    .B(_13769_),
    .X(_09647_));
 sky130_fd_sc_hd__a221oi_1 _23667_ (.A1(_13769_),
    .A2(_13761_),
    .B1(_09643_),
    .B2(_09647_),
    .C1(_13768_),
    .Y(_09648_));
 sky130_fd_sc_hd__xnor2_1 _23668_ (.A(_13775_),
    .B(_09648_),
    .Y(\hash.CA1.p5[18] ));
 sky130_fd_sc_hd__clkinv_1 _23669_ (.A(_13780_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21o_1 _23670_ (.A1(_13755_),
    .A2(_13747_),
    .B1(_13754_),
    .X(_09650_));
 sky130_fd_sc_hd__a21o_1 _23671_ (.A1(_13762_),
    .A2(_09650_),
    .B1(_13761_),
    .X(_09651_));
 sky130_fd_sc_hd__a21o_1 _23672_ (.A1(_13769_),
    .A2(_09651_),
    .B1(_13768_),
    .X(_09652_));
 sky130_fd_sc_hd__a21oi_2 _23673_ (.A1(_13775_),
    .A2(_09652_),
    .B1(_13774_),
    .Y(_09653_));
 sky130_fd_sc_hd__and4_4 _23674_ (.A(_13748_),
    .B(_13755_),
    .C(_13775_),
    .D(_09647_),
    .X(_09654_));
 sky130_fd_sc_hd__nand2b_1 _23675_ (.A_N(_09639_),
    .B(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _23676_ (.A(_09653_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__xnor2_1 _23677_ (.A(_09649_),
    .B(_09656_),
    .Y(\hash.CA1.p5[19] ));
 sky130_fd_sc_hd__o21bai_1 _23678_ (.A1(_09649_),
    .A2(_09653_),
    .B1_N(_13779_),
    .Y(_09657_));
 sky130_fd_sc_hd__a31oi_1 _23679_ (.A1(_13780_),
    .A2(_09634_),
    .A3(_09654_),
    .B1(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__xnor2_1 _23680_ (.A(_13785_),
    .B(_09658_),
    .Y(\hash.CA1.p5[20] ));
 sky130_fd_sc_hd__nand3_1 _23681_ (.A(_13780_),
    .B(_13785_),
    .C(_09654_),
    .Y(_09659_));
 sky130_fd_sc_hd__a21oi_1 _23682_ (.A1(_13785_),
    .A2(_09657_),
    .B1(_13784_),
    .Y(_09660_));
 sky130_fd_sc_hd__o21ai_2 _23683_ (.A1(_09639_),
    .A2(_09659_),
    .B1(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__xor2_1 _23684_ (.A(_13790_),
    .B(_09661_),
    .X(\hash.CA1.p5[21] ));
 sky130_fd_sc_hd__o2111ai_2 _23685_ (.A1(_09630_),
    .A2(_09632_),
    .B1(_09654_),
    .C1(_13780_),
    .D1(_13742_),
    .Y(_09662_));
 sky130_fd_sc_hd__nor2_1 _23686_ (.A(_09649_),
    .B(_09653_),
    .Y(_09663_));
 sky130_fd_sc_hd__a31oi_1 _23687_ (.A1(_13780_),
    .A2(_13741_),
    .A3(_09654_),
    .B1(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__nor3_1 _23688_ (.A(_13779_),
    .B(_13784_),
    .C(_13789_),
    .Y(_09665_));
 sky130_fd_sc_hd__or2_0 _23689_ (.A(_13785_),
    .B(_13784_),
    .X(_09666_));
 sky130_fd_sc_hd__a21oi_1 _23690_ (.A1(_13790_),
    .A2(_09666_),
    .B1(_13789_),
    .Y(_09667_));
 sky130_fd_sc_hd__a31oi_2 _23691_ (.A1(_09662_),
    .A2(_09664_),
    .A3(_09665_),
    .B1(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__xor2_1 _23692_ (.A(_13795_),
    .B(_09668_),
    .X(\hash.CA1.p5[22] ));
 sky130_fd_sc_hd__inv_1 _23693_ (.A(_13801_),
    .Y(_09669_));
 sky130_fd_sc_hd__a21oi_1 _23694_ (.A1(_13795_),
    .A2(_13789_),
    .B1(_13794_),
    .Y(_09670_));
 sky130_fd_sc_hd__nand3_1 _23695_ (.A(_13790_),
    .B(_13795_),
    .C(_09661_),
    .Y(_09671_));
 sky130_fd_sc_hd__nand2_1 _23696_ (.A(_09670_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__xnor2_1 _23697_ (.A(_09669_),
    .B(_09672_),
    .Y(\hash.CA1.p5[23] ));
 sky130_fd_sc_hd__a21o_1 _23698_ (.A1(_13795_),
    .A2(_09668_),
    .B1(_13794_),
    .X(_09673_));
 sky130_fd_sc_hd__a21oi_1 _23699_ (.A1(_13801_),
    .A2(_09673_),
    .B1(_13800_),
    .Y(_09674_));
 sky130_fd_sc_hd__xnor2_1 _23700_ (.A(_13808_),
    .B(_09674_),
    .Y(\hash.CA1.p5[24] ));
 sky130_fd_sc_hd__nand2_1 _23701_ (.A(_13801_),
    .B(_13808_),
    .Y(_09675_));
 sky130_fd_sc_hd__o21bai_1 _23702_ (.A1(_09669_),
    .A2(_09670_),
    .B1_N(_13800_),
    .Y(_09676_));
 sky130_fd_sc_hd__a21oi_1 _23703_ (.A1(_13808_),
    .A2(_09676_),
    .B1(_13807_),
    .Y(_09677_));
 sky130_fd_sc_hd__o21ai_0 _23704_ (.A1(_09671_),
    .A2(_09675_),
    .B1(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__xor2_1 _23705_ (.A(_13815_),
    .B(_09678_),
    .X(\hash.CA1.p5[25] ));
 sky130_fd_sc_hd__and2_4 _23706_ (.A(_13801_),
    .B(_13808_),
    .X(_09679_));
 sky130_fd_sc_hd__nand4_1 _23707_ (.A(_13795_),
    .B(_13815_),
    .C(_09668_),
    .D(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__a21oi_1 _23708_ (.A1(_13808_),
    .A2(_13800_),
    .B1(_13807_),
    .Y(_09681_));
 sky130_fd_sc_hd__nor2b_1 _23709_ (.A(_09681_),
    .B_N(_13815_),
    .Y(_09682_));
 sky130_fd_sc_hd__a31oi_1 _23710_ (.A1(_13815_),
    .A2(_13794_),
    .A3(_09679_),
    .B1(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__nand2_1 _23711_ (.A(_09680_),
    .B(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__nor2_1 _23712_ (.A(_13814_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__xnor2_1 _23713_ (.A(_13822_),
    .B(_09685_),
    .Y(\hash.CA1.p5[26] ));
 sky130_fd_sc_hd__nand2_1 _23714_ (.A(_13790_),
    .B(_13795_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand2_1 _23715_ (.A(_13815_),
    .B(_09679_),
    .Y(_09687_));
 sky130_fd_sc_hd__nor3b_1 _23716_ (.A(_09686_),
    .B(_09687_),
    .C_N(_09661_),
    .Y(_09688_));
 sky130_fd_sc_hd__nor2b_1 _23717_ (.A(_09677_),
    .B_N(_13815_),
    .Y(_09689_));
 sky130_fd_sc_hd__o31ai_1 _23718_ (.A1(_13814_),
    .A2(_09688_),
    .A3(_09689_),
    .B1(_13822_),
    .Y(_09690_));
 sky130_fd_sc_hd__nor2b_1 _23719_ (.A(_13821_),
    .B_N(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__xnor2_1 _23720_ (.A(_13829_),
    .B(_09691_),
    .Y(\hash.CA1.p5[27] ));
 sky130_fd_sc_hd__nor3_1 _23721_ (.A(_13814_),
    .B(_13821_),
    .C(_13828_),
    .Y(_09692_));
 sky130_fd_sc_hd__or2_0 _23722_ (.A(_13829_),
    .B(_13828_),
    .X(_09693_));
 sky130_fd_sc_hd__o31ai_1 _23723_ (.A1(_13822_),
    .A2(_13821_),
    .A3(_13828_),
    .B1(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__a31oi_1 _23724_ (.A1(_09680_),
    .A2(_09683_),
    .A3(_09692_),
    .B1(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__xor2_1 _23725_ (.A(_13836_),
    .B(_09695_),
    .X(\hash.CA1.p5[28] ));
 sky130_fd_sc_hd__inv_1 _23726_ (.A(_13842_),
    .Y(_09696_));
 sky130_fd_sc_hd__nor3_1 _23727_ (.A(_13821_),
    .B(_13828_),
    .C(_13835_),
    .Y(_09697_));
 sky130_fd_sc_hd__a21oi_1 _23728_ (.A1(_13836_),
    .A2(_09693_),
    .B1(_13835_),
    .Y(_09698_));
 sky130_fd_sc_hd__a21oi_1 _23729_ (.A1(_09690_),
    .A2(_09697_),
    .B1(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__xnor2_1 _23730_ (.A(_09696_),
    .B(_09699_),
    .Y(\hash.CA1.p5[29] ));
 sky130_fd_sc_hd__xnor2_1 _23731_ (.A(_12896_),
    .B(_13675_),
    .Y(\hash.CA1.p5[2] ));
 sky130_fd_sc_hd__a21oi_1 _23732_ (.A1(_13836_),
    .A2(_09695_),
    .B1(_13835_),
    .Y(_09700_));
 sky130_fd_sc_hd__o21bai_1 _23733_ (.A1(_09696_),
    .A2(_09700_),
    .B1_N(_13841_),
    .Y(_09701_));
 sky130_fd_sc_hd__xor2_1 _23734_ (.A(_13847_),
    .B(_09701_),
    .X(\hash.CA1.p5[30] ));
 sky130_fd_sc_hd__a21o_1 _23735_ (.A1(_13842_),
    .A2(_09699_),
    .B1(_13841_),
    .X(_09702_));
 sky130_fd_sc_hd__a21oi_1 _23736_ (.A1(_13847_),
    .A2(_09702_),
    .B1(_13846_),
    .Y(_09703_));
 sky130_fd_sc_hd__nand2_1 _23737_ (.A(_06002_),
    .B(\hash.CA2.a_dash[31] ),
    .Y(_09704_));
 sky130_fd_sc_hd__xnor2_1 _23738_ (.A(_09703_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__xnor2_1 _23739_ (.A(\hash.CA1.p4[31] ),
    .B(_09705_),
    .Y(\hash.CA1.p5[31] ));
 sky130_fd_sc_hd__xnor2_1 _23740_ (.A(_13681_),
    .B(_09610_),
    .Y(\hash.CA1.p5[3] ));
 sky130_fd_sc_hd__nand2_1 _23741_ (.A(_09599_),
    .B(_09601_),
    .Y(_09706_));
 sky130_fd_sc_hd__nor2_1 _23742_ (.A(_13687_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__nor2_1 _23743_ (.A(_09602_),
    .B(_09707_),
    .Y(\hash.CA1.p5[4] ));
 sky130_fd_sc_hd__xnor2_1 _23744_ (.A(_13693_),
    .B(_09612_),
    .Y(\hash.CA1.p5[5] ));
 sky130_fd_sc_hd__nor2_1 _23745_ (.A(_13692_),
    .B(_09603_),
    .Y(_09708_));
 sky130_fd_sc_hd__xnor2_1 _23746_ (.A(_13699_),
    .B(_09708_),
    .Y(\hash.CA1.p5[6] ));
 sky130_fd_sc_hd__xor2_1 _23747_ (.A(_13705_),
    .B(_09621_),
    .X(\hash.CA1.p5[7] ));
 sky130_fd_sc_hd__nand2_1 _23748_ (.A(_09598_),
    .B(_09604_),
    .Y(_09709_));
 sky130_fd_sc_hd__a21oi_1 _23749_ (.A1(_13705_),
    .A2(_09709_),
    .B1(_13704_),
    .Y(_09710_));
 sky130_fd_sc_hd__xnor2_1 _23750_ (.A(_13712_),
    .B(_09710_),
    .Y(\hash.CA1.p5[8] ));
 sky130_fd_sc_hd__inv_1 _23751_ (.A(_13712_),
    .Y(_09711_));
 sky130_fd_sc_hd__a21oi_1 _23752_ (.A1(_13705_),
    .A2(_09621_),
    .B1(_13704_),
    .Y(_09712_));
 sky130_fd_sc_hd__o21bai_1 _23753_ (.A1(_09711_),
    .A2(_09712_),
    .B1_N(_13711_),
    .Y(_09713_));
 sky130_fd_sc_hd__xor2_1 _23754_ (.A(_13718_),
    .B(_09713_),
    .X(\hash.CA1.p5[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_637 ();
 sky130_fd_sc_hd__or2_0 _23764_ (.A(\hash.CA2.b_dash[1] ),
    .B(net355),
    .X(_12657_));
 sky130_fd_sc_hd__inv_1 _23765_ (.A(_12657_),
    .Y(_00751_));
 sky130_fd_sc_hd__or2_4 _23766_ (.A(net349),
    .B(\hash.CA2.a_dash[1] ),
    .X(_12899_));
 sky130_fd_sc_hd__clkinv_1 _23767_ (.A(_12899_),
    .Y(_00721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_636 ();
 sky130_fd_sc_hd__or2_4 _23769_ (.A(net349),
    .B(_12922_),
    .X(\hash.CA1.b[0] ));
 sky130_fd_sc_hd__inv_1 _23770_ (.A(\hash.CA1.b[0] ),
    .Y(_00690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_634 ();
 sky130_fd_sc_hd__nand4_1 _23773_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_13541_),
    .D(\count_2[5] ),
    .Y(_09726_));
 sky130_fd_sc_hd__or2_4 _23774_ (.A(\count_2[6] ),
    .B(_09726_),
    .X(_09727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_633 ();
 sky130_fd_sc_hd__clkinv_2 _23776_ (.A(_09727_),
    .Y(_00128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_631 ();
 sky130_fd_sc_hd__clkinv_16 _23779_ (.A(net1044),
    .Y(_09731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_627 ();
 sky130_fd_sc_hd__nor3_4 _23784_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_2 _23785_ (.A(_13528_),
    .B(_09735_),
    .Y(_09736_));
 sky130_fd_sc_hd__nand2_8 _23786_ (.A(_09731_),
    .B(_09736_),
    .Y(_00127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_625 ();
 sky130_fd_sc_hd__nor3b_4 _23789_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C_N(\count_1[3] ),
    .Y(_09739_));
 sky130_fd_sc_hd__nand2_4 _23790_ (.A(_13531_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nand2_8 _23791_ (.A(_09731_),
    .B(_09740_),
    .Y(_00126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_624 ();
 sky130_fd_sc_hd__nand2_2 _23793_ (.A(_13529_),
    .B(_09739_),
    .Y(_09742_));
 sky130_fd_sc_hd__nand2_8 _23794_ (.A(_09731_),
    .B(_09742_),
    .Y(_00125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_623 ();
 sky130_fd_sc_hd__nand2_2 _23796_ (.A(_13533_),
    .B(_09739_),
    .Y(_09744_));
 sky130_fd_sc_hd__nand2_8 _23797_ (.A(_09731_),
    .B(_09744_),
    .Y(_00124_));
 sky130_fd_sc_hd__nor3b_4 _23798_ (.A(\count_1[5] ),
    .B(\count_1[3] ),
    .C_N(\count_1[4] ),
    .Y(_09745_));
 sky130_fd_sc_hd__nand2_2 _23799_ (.A(_13528_),
    .B(_09745_),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_8 _23800_ (.A(_09731_),
    .B(_09746_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_2 _23801_ (.A(_13531_),
    .B(_09745_),
    .Y(_09747_));
 sky130_fd_sc_hd__nand2_8 _23802_ (.A(_09731_),
    .B(_09747_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_4 _23803_ (.A(_13529_),
    .B(_09745_),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_8 _23804_ (.A(_09731_),
    .B(_09748_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_2 _23805_ (.A(_13533_),
    .B(_09745_),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_8 _23806_ (.A(_09731_),
    .B(_09749_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _23807_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .Y(_09750_));
 sky130_fd_sc_hd__nor2_4 _23808_ (.A(\count_1[5] ),
    .B(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__nand2_4 _23809_ (.A(_13528_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__nand2_8 _23810_ (.A(_09731_),
    .B(_09752_),
    .Y(_00119_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_621 ();
 sky130_fd_sc_hd__nand2_4 _23813_ (.A(_13531_),
    .B(_09751_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand2_8 _23814_ (.A(_09731_),
    .B(_09755_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_4 _23815_ (.A(_13529_),
    .B(_09751_),
    .Y(_09756_));
 sky130_fd_sc_hd__nand2_8 _23816_ (.A(_09731_),
    .B(_09756_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_4 _23817_ (.A(_13531_),
    .B(_09735_),
    .Y(_09757_));
 sky130_fd_sc_hd__nand2_8 _23818_ (.A(_09731_),
    .B(_09757_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_4 _23819_ (.A(_13533_),
    .B(_09751_),
    .Y(_09758_));
 sky130_fd_sc_hd__nand2_8 _23820_ (.A(_09731_),
    .B(_09758_),
    .Y(_00115_));
 sky130_fd_sc_hd__nor3b_4 _23821_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C_N(\count_1[5] ),
    .Y(_09759_));
 sky130_fd_sc_hd__nand2_4 _23822_ (.A(_13528_),
    .B(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__nand2_8 _23823_ (.A(_09731_),
    .B(_09760_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_4 _23824_ (.A(_13531_),
    .B(_09759_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_8 _23825_ (.A(_09731_),
    .B(_09761_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_4 _23826_ (.A(_13529_),
    .B(_09759_),
    .Y(_09762_));
 sky130_fd_sc_hd__nand2_8 _23827_ (.A(_09731_),
    .B(_09762_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_2 _23828_ (.A(_13533_),
    .B(_09759_),
    .Y(_09763_));
 sky130_fd_sc_hd__nand2_8 _23829_ (.A(_09731_),
    .B(_09763_),
    .Y(_00111_));
 sky130_fd_sc_hd__and3b_4 _23830_ (.A_N(\count_1[4] ),
    .B(\count_1[3] ),
    .C(\count_1[5] ),
    .X(_09764_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_620 ();
 sky130_fd_sc_hd__nand2_2 _23832_ (.A(_13528_),
    .B(_09764_),
    .Y(_09766_));
 sky130_fd_sc_hd__nand2_8 _23833_ (.A(_09731_),
    .B(_09766_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_4 _23834_ (.A(_13531_),
    .B(_09764_),
    .Y(_09767_));
 sky130_fd_sc_hd__nand2_8 _23835_ (.A(_09731_),
    .B(_09767_),
    .Y(_00109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_619 ();
 sky130_fd_sc_hd__nand2_2 _23837_ (.A(_13529_),
    .B(_09764_),
    .Y(_09769_));
 sky130_fd_sc_hd__nand2_8 _23838_ (.A(_09731_),
    .B(_09769_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_2 _23839_ (.A(_13533_),
    .B(_09764_),
    .Y(_09770_));
 sky130_fd_sc_hd__nand2_8 _23840_ (.A(_09731_),
    .B(_09770_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3b_4 _23841_ (.A_N(\count_1[3] ),
    .B(\count_1[4] ),
    .C(\count_1[5] ),
    .X(_09771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_618 ();
 sky130_fd_sc_hd__nand2_2 _23843_ (.A(_13528_),
    .B(_09771_),
    .Y(_09773_));
 sky130_fd_sc_hd__nand2_8 _23844_ (.A(_09731_),
    .B(_09773_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_2 _23845_ (.A(_13529_),
    .B(_09735_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand2_8 _23846_ (.A(_09731_),
    .B(_09774_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_2 _23847_ (.A(_13531_),
    .B(_09771_),
    .Y(_09775_));
 sky130_fd_sc_hd__nand2_8 _23848_ (.A(_09731_),
    .B(_09775_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_2 _23849_ (.A(_13529_),
    .B(_09771_),
    .Y(_09776_));
 sky130_fd_sc_hd__nand2_8 _23850_ (.A(_09731_),
    .B(_09776_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_4 _23851_ (.A(_13533_),
    .B(_09771_),
    .Y(_09777_));
 sky130_fd_sc_hd__nand2_8 _23852_ (.A(_09731_),
    .B(_09777_),
    .Y(_00102_));
 sky130_fd_sc_hd__and3_4 _23853_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .X(_09778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_617 ();
 sky130_fd_sc_hd__nand2_2 _23855_ (.A(_13528_),
    .B(_09778_),
    .Y(_09780_));
 sky130_fd_sc_hd__nand2_8 _23856_ (.A(_09731_),
    .B(_09780_),
    .Y(_00101_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_614 ();
 sky130_fd_sc_hd__nor3b_4 _23860_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .C_N(\count_2[3] ),
    .Y(_09784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_613 ();
 sky130_fd_sc_hd__nand2_4 _23862_ (.A(_13539_),
    .B(_09784_),
    .Y(_09786_));
 sky130_fd_sc_hd__nand2_8 _23863_ (.A(_09731_),
    .B(_09786_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_4 _23864_ (.A(_13531_),
    .B(_09778_),
    .Y(_09787_));
 sky130_fd_sc_hd__nand2_8 _23865_ (.A(_09731_),
    .B(_09787_),
    .Y(_00100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_611 ();
 sky130_fd_sc_hd__nand2_2 _23868_ (.A(_13537_),
    .B(_09784_),
    .Y(_09790_));
 sky130_fd_sc_hd__nand2_8 _23869_ (.A(_09731_),
    .B(_09790_),
    .Y(_00094_));
 sky130_fd_sc_hd__nand2_2 _23870_ (.A(_13541_),
    .B(_09784_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand2_8 _23871_ (.A(_09731_),
    .B(_09791_),
    .Y(_00093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_610 ();
 sky130_fd_sc_hd__nand2b_4 _23873_ (.A_N(\count_2[3] ),
    .B(\count_2[4] ),
    .Y(_09793_));
 sky130_fd_sc_hd__nor2_4 _23874_ (.A(\count_2[5] ),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__nand2_4 _23875_ (.A(_13536_),
    .B(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__nand2_8 _23876_ (.A(_09731_),
    .B(_09795_),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_2 _23877_ (.A(_13539_),
    .B(_09794_),
    .Y(_09796_));
 sky130_fd_sc_hd__nand2_8 _23878_ (.A(_09731_),
    .B(_09796_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor3_4 _23879_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(\count_2[5] ),
    .Y(_09797_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_609 ();
 sky130_fd_sc_hd__nand2_4 _23881_ (.A(_13536_),
    .B(_09797_),
    .Y(_09799_));
 sky130_fd_sc_hd__nand2_8 _23882_ (.A(_09731_),
    .B(_09799_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_2 _23883_ (.A(_13537_),
    .B(_09794_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_8 _23884_ (.A(_09731_),
    .B(_09800_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_4 _23885_ (.A(_13529_),
    .B(_09778_),
    .Y(_09801_));
 sky130_fd_sc_hd__nand2_8 _23886_ (.A(_09731_),
    .B(_09801_),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_8 _23887_ (.A(\count_2[5] ),
    .Y(_09802_));
 sky130_fd_sc_hd__nand2_4 _23888_ (.A(_13541_),
    .B(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__o21ai_4 _23889_ (.A1(_09793_),
    .A2(_09803_),
    .B1(_09731_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_4 _23890_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .Y(_09804_));
 sky130_fd_sc_hd__nor2_4 _23891_ (.A(\count_2[5] ),
    .B(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__nand2_4 _23892_ (.A(_13536_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_8 _23893_ (.A(_09731_),
    .B(_09806_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand2_4 _23894_ (.A(_13539_),
    .B(_09805_),
    .Y(_09807_));
 sky130_fd_sc_hd__nand2_8 _23895_ (.A(_09731_),
    .B(_09807_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_2 _23896_ (.A(_13537_),
    .B(_09805_),
    .Y(_09808_));
 sky130_fd_sc_hd__nand2_8 _23897_ (.A(_09731_),
    .B(_09808_),
    .Y(_00085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_608 ();
 sky130_fd_sc_hd__nand2_4 _23899_ (.A(_13541_),
    .B(_09805_),
    .Y(_09810_));
 sky130_fd_sc_hd__nand2_8 _23900_ (.A(_09731_),
    .B(_09810_),
    .Y(_00084_));
 sky130_fd_sc_hd__nor3_4 _23901_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_09802_),
    .Y(_09811_));
 sky130_fd_sc_hd__nand2_4 _23902_ (.A(_13536_),
    .B(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__nand2_8 _23903_ (.A(_09731_),
    .B(_09812_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_4 _23904_ (.A(_13533_),
    .B(_09778_),
    .Y(_09813_));
 sky130_fd_sc_hd__nand2_8 _23905_ (.A(_09731_),
    .B(_09813_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_2 _23906_ (.A(_13539_),
    .B(_09811_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2_8 _23907_ (.A(_09731_),
    .B(_09814_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand2_4 _23908_ (.A(_13537_),
    .B(_09811_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand2_8 _23909_ (.A(_09731_),
    .B(_09815_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_4 _23910_ (.A(_13541_),
    .B(\count_2[5] ),
    .Y(_09816_));
 sky130_fd_sc_hd__o31ai_4 _23911_ (.A1(\count_2[4] ),
    .A2(\count_2[3] ),
    .A3(_09816_),
    .B1(_09731_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_2 _23912_ (.A(_13539_),
    .B(_09797_),
    .Y(_09817_));
 sky130_fd_sc_hd__nand2_8 _23913_ (.A(_09731_),
    .B(_09817_),
    .Y(_00079_));
 sky130_fd_sc_hd__nor3b_4 _23914_ (.A(_09802_),
    .B(\count_2[4] ),
    .C_N(\count_2[3] ),
    .Y(_09818_));
 sky130_fd_sc_hd__nand2_4 _23915_ (.A(_13536_),
    .B(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__nand2_8 _23916_ (.A(_09731_),
    .B(_09819_),
    .Y(_00078_));
 sky130_fd_sc_hd__nand2_2 _23917_ (.A(_13539_),
    .B(_09818_),
    .Y(_09820_));
 sky130_fd_sc_hd__nand2_8 _23918_ (.A(_09731_),
    .B(_09820_),
    .Y(_00077_));
 sky130_fd_sc_hd__nand2_4 _23919_ (.A(_13533_),
    .B(_09735_),
    .Y(_09821_));
 sky130_fd_sc_hd__nand2_8 _23920_ (.A(_09731_),
    .B(_09821_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_4 _23921_ (.A(_13537_),
    .B(_09818_),
    .Y(_09822_));
 sky130_fd_sc_hd__nand2_8 _23922_ (.A(_09731_),
    .B(_09822_),
    .Y(_00076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_607 ();
 sky130_fd_sc_hd__nand2_4 _23924_ (.A(_13541_),
    .B(_09818_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_8 _23925_ (.A(_09731_),
    .B(_09824_),
    .Y(_00075_));
 sky130_fd_sc_hd__nor2_4 _23926_ (.A(_09802_),
    .B(_09793_),
    .Y(_09825_));
 sky130_fd_sc_hd__nand2_2 _23927_ (.A(_13536_),
    .B(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__nand2_8 _23928_ (.A(_09731_),
    .B(_09826_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_2 _23929_ (.A(_13539_),
    .B(_09825_),
    .Y(_09827_));
 sky130_fd_sc_hd__nand2_8 _23930_ (.A(_09731_),
    .B(_09827_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_2 _23931_ (.A(_13537_),
    .B(_09825_),
    .Y(_09828_));
 sky130_fd_sc_hd__nand2_8 _23932_ (.A(_09731_),
    .B(_09828_),
    .Y(_00072_));
 sky130_fd_sc_hd__o21ai_4 _23933_ (.A1(_09816_),
    .A2(_09793_),
    .B1(_09731_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand2_2 _23934_ (.A(_13528_),
    .B(_09739_),
    .Y(_09829_));
 sky130_fd_sc_hd__nand2_8 _23935_ (.A(_09731_),
    .B(_09829_),
    .Y(_00096_));
 sky130_fd_sc_hd__nor2_4 _23936_ (.A(_09802_),
    .B(_09804_),
    .Y(_09830_));
 sky130_fd_sc_hd__nand2_4 _23937_ (.A(_13536_),
    .B(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__nand2_8 _23938_ (.A(_09731_),
    .B(_09831_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_4 _23939_ (.A(_13539_),
    .B(_09830_),
    .Y(_09832_));
 sky130_fd_sc_hd__nand2_8 _23940_ (.A(_09731_),
    .B(_09832_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_4 _23941_ (.A(_13537_),
    .B(_09797_),
    .Y(_09833_));
 sky130_fd_sc_hd__nand2_8 _23942_ (.A(_09731_),
    .B(_09833_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_2 _23943_ (.A(_13537_),
    .B(_09830_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_8 _23944_ (.A(_09731_),
    .B(_09834_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_8 _23945_ (.A(_09731_),
    .B(_09726_),
    .Y(_00066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_606 ();
 sky130_fd_sc_hd__nor3_4 _23947_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_09803_),
    .Y(_09836_));
 sky130_fd_sc_hd__or2_4 _23948_ (.A(net1043),
    .B(_09836_),
    .X(_00065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_605 ();
 sky130_fd_sc_hd__nand2_2 _23950_ (.A(_13536_),
    .B(_09784_),
    .Y(_09838_));
 sky130_fd_sc_hd__nand2_8 _23951_ (.A(_09731_),
    .B(_09838_),
    .Y(_00064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_600 ();
 sky130_fd_sc_hd__mux4_2 _23957_ (.A0(\w[19][0] ),
    .A1(\w[17][0] ),
    .A2(\w[23][0] ),
    .A3(\w[21][0] ),
    .S0(net368),
    .S1(net314),
    .X(_09844_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_598 ();
 sky130_fd_sc_hd__mux4_2 _23960_ (.A0(\w[27][0] ),
    .A1(\w[25][0] ),
    .A2(\w[31][0] ),
    .A3(\w[29][0] ),
    .S0(net368),
    .S1(net314),
    .X(_09847_));
 sky130_fd_sc_hd__mux4_2 _23961_ (.A0(\w[3][0] ),
    .A1(\w[1][0] ),
    .A2(\w[7][0] ),
    .A3(\w[5][0] ),
    .S0(net368),
    .S1(net314),
    .X(_09848_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_595 ();
 sky130_fd_sc_hd__mux4_2 _23965_ (.A0(\w[11][0] ),
    .A1(\w[9][0] ),
    .A2(\w[15][0] ),
    .A3(\w[13][0] ),
    .S0(net368),
    .S1(net314),
    .X(_09852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_594 ();
 sky130_fd_sc_hd__xor2_4 _23967_ (.A(\count_hash2[3] ),
    .B(_12908_),
    .X(_09854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_593 ();
 sky130_fd_sc_hd__nand3_4 _23969_ (.A(\count_hash2[3] ),
    .B(\count_hash2[2] ),
    .C(\count_hash2[1] ),
    .Y(_09856_));
 sky130_fd_sc_hd__xor2_4 _23970_ (.A(\count_hash2[4] ),
    .B(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_592 ();
 sky130_fd_sc_hd__mux4_2 _23972_ (.A0(_09844_),
    .A1(_09847_),
    .A2(_09848_),
    .A3(_09852_),
    .S0(net344),
    .S1(net335),
    .X(_09859_));
 sky130_fd_sc_hd__mux4_2 _23973_ (.A0(\w[51][0] ),
    .A1(\w[49][0] ),
    .A2(\w[55][0] ),
    .A3(\w[53][0] ),
    .S0(net369),
    .S1(net315),
    .X(_09860_));
 sky130_fd_sc_hd__mux4_2 _23974_ (.A0(\w[59][0] ),
    .A1(\w[57][0] ),
    .A2(\w[63][0] ),
    .A3(\w[61][0] ),
    .S0(net369),
    .S1(net315),
    .X(_09861_));
 sky130_fd_sc_hd__mux4_2 _23975_ (.A0(\w[35][0] ),
    .A1(\w[33][0] ),
    .A2(\w[39][0] ),
    .A3(\w[37][0] ),
    .S0(net369),
    .S1(net315),
    .X(_09862_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_591 ();
 sky130_fd_sc_hd__mux4_2 _23977_ (.A0(\w[43][0] ),
    .A1(\w[41][0] ),
    .A2(\w[47][0] ),
    .A3(\w[45][0] ),
    .S0(net369),
    .S1(net315),
    .X(_09864_));
 sky130_fd_sc_hd__mux4_2 _23978_ (.A0(_09860_),
    .A1(_09861_),
    .A2(_09862_),
    .A3(_09864_),
    .S0(net343),
    .S1(net337),
    .X(_09865_));
 sky130_fd_sc_hd__nand3_4 _23979_ (.A(\count_hash2[4] ),
    .B(\count_hash2[3] ),
    .C(_12908_),
    .Y(_09866_));
 sky130_fd_sc_hd__xnor2_1 _23980_ (.A(\count_hash2[5] ),
    .B(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_589 ();
 sky130_fd_sc_hd__mux2i_1 _23983_ (.A0(_09859_),
    .A1(_09865_),
    .S(net297),
    .Y(_09870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_587 ();
 sky130_fd_sc_hd__nand4_1 _23986_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(\count_hash1[5] ),
    .D(\count_hash1[2] ),
    .Y(_09873_));
 sky130_fd_sc_hd__nor2_2 _23987_ (.A(_12914_),
    .B(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__or3_4 _23988_ (.A(\count_hash1[6] ),
    .B(net540),
    .C(_09874_),
    .X(_09875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_584 ();
 sky130_fd_sc_hd__nand2_2 _23992_ (.A(net357),
    .B(\w[1][0] ),
    .Y(_09879_));
 sky130_fd_sc_hd__o21ai_4 _23993_ (.A1(_09870_),
    .A2(net292),
    .B1(_09879_),
    .Y(_00032_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_580 ();
 sky130_fd_sc_hd__mux4_2 _23998_ (.A0(\w[19][1] ),
    .A1(\w[17][1] ),
    .A2(\w[23][1] ),
    .A3(\w[21][1] ),
    .S0(net368),
    .S1(net314),
    .X(_09884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_578 ();
 sky130_fd_sc_hd__mux4_2 _24001_ (.A0(\w[27][1] ),
    .A1(\w[25][1] ),
    .A2(\w[31][1] ),
    .A3(\w[29][1] ),
    .S0(net368),
    .S1(net314),
    .X(_09887_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_576 ();
 sky130_fd_sc_hd__mux4_2 _24004_ (.A0(\w[3][1] ),
    .A1(\w[1][1] ),
    .A2(\w[7][1] ),
    .A3(\w[5][1] ),
    .S0(net368),
    .S1(net314),
    .X(_09890_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_574 ();
 sky130_fd_sc_hd__mux4_2 _24007_ (.A0(\w[11][1] ),
    .A1(\w[9][1] ),
    .A2(\w[15][1] ),
    .A3(\w[13][1] ),
    .S0(net368),
    .S1(net314),
    .X(_09893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_572 ();
 sky130_fd_sc_hd__mux4_2 _24010_ (.A0(_09884_),
    .A1(_09887_),
    .A2(_09890_),
    .A3(_09893_),
    .S0(net343),
    .S1(net334),
    .X(_09896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_570 ();
 sky130_fd_sc_hd__mux4_2 _24013_ (.A0(\w[51][1] ),
    .A1(\w[49][1] ),
    .A2(\w[55][1] ),
    .A3(\w[53][1] ),
    .S0(net369),
    .S1(net315),
    .X(_09899_));
 sky130_fd_sc_hd__mux4_2 _24014_ (.A0(\w[59][1] ),
    .A1(\w[57][1] ),
    .A2(\w[63][1] ),
    .A3(\w[61][1] ),
    .S0(net369),
    .S1(net315),
    .X(_09900_));
 sky130_fd_sc_hd__mux4_2 _24015_ (.A0(\w[35][1] ),
    .A1(\w[33][1] ),
    .A2(\w[39][1] ),
    .A3(\w[37][1] ),
    .S0(net369),
    .S1(net315),
    .X(_09901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_568 ();
 sky130_fd_sc_hd__mux4_2 _24018_ (.A0(\w[43][1] ),
    .A1(\w[41][1] ),
    .A2(\w[47][1] ),
    .A3(\w[45][1] ),
    .S0(net369),
    .S1(net315),
    .X(_09904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_565 ();
 sky130_fd_sc_hd__mux4_2 _24022_ (.A0(_09899_),
    .A1(_09900_),
    .A2(_09901_),
    .A3(_09904_),
    .S0(net343),
    .S1(net337),
    .X(_09908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_564 ();
 sky130_fd_sc_hd__mux2i_1 _24024_ (.A0(_09896_),
    .A1(_09908_),
    .S(net297),
    .Y(_09910_));
 sky130_fd_sc_hd__nand2_2 _24025_ (.A(net357),
    .B(\w[1][1] ),
    .Y(_09911_));
 sky130_fd_sc_hd__o21ai_4 _24026_ (.A1(net292),
    .A2(_09910_),
    .B1(_09911_),
    .Y(_00043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_563 ();
 sky130_fd_sc_hd__mux4_2 _24028_ (.A0(\w[19][2] ),
    .A1(\w[17][2] ),
    .A2(\w[23][2] ),
    .A3(\w[21][2] ),
    .S0(net368),
    .S1(net314),
    .X(_09913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_562 ();
 sky130_fd_sc_hd__mux4_2 _24030_ (.A0(\w[27][2] ),
    .A1(\w[25][2] ),
    .A2(\w[31][2] ),
    .A3(\w[29][2] ),
    .S0(net368),
    .S1(net314),
    .X(_09915_));
 sky130_fd_sc_hd__mux4_2 _24031_ (.A0(\w[3][2] ),
    .A1(\w[1][2] ),
    .A2(\w[7][2] ),
    .A3(\w[5][2] ),
    .S0(net368),
    .S1(net314),
    .X(_09916_));
 sky130_fd_sc_hd__mux4_2 _24032_ (.A0(\w[11][2] ),
    .A1(\w[9][2] ),
    .A2(\w[15][2] ),
    .A3(\w[13][2] ),
    .S0(net368),
    .S1(net314),
    .X(_09917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_561 ();
 sky130_fd_sc_hd__mux4_2 _24034_ (.A0(_09913_),
    .A1(_09915_),
    .A2(_09916_),
    .A3(_09917_),
    .S0(net343),
    .S1(net334),
    .X(_09919_));
 sky130_fd_sc_hd__mux4_2 _24035_ (.A0(\w[51][2] ),
    .A1(\w[49][2] ),
    .A2(\w[55][2] ),
    .A3(\w[53][2] ),
    .S0(net369),
    .S1(net315),
    .X(_09920_));
 sky130_fd_sc_hd__mux4_2 _24036_ (.A0(\w[59][2] ),
    .A1(\w[57][2] ),
    .A2(\w[63][2] ),
    .A3(\w[61][2] ),
    .S0(net369),
    .S1(net315),
    .X(_09921_));
 sky130_fd_sc_hd__mux4_2 _24037_ (.A0(\w[35][2] ),
    .A1(\w[33][2] ),
    .A2(\w[39][2] ),
    .A3(\w[37][2] ),
    .S0(net369),
    .S1(net315),
    .X(_09922_));
 sky130_fd_sc_hd__mux4_2 _24038_ (.A0(\w[43][2] ),
    .A1(\w[41][2] ),
    .A2(\w[47][2] ),
    .A3(\w[45][2] ),
    .S0(net369),
    .S1(net315),
    .X(_09923_));
 sky130_fd_sc_hd__mux4_2 _24039_ (.A0(_09920_),
    .A1(_09921_),
    .A2(_09922_),
    .A3(_09923_),
    .S0(net346),
    .S1(net337),
    .X(_09924_));
 sky130_fd_sc_hd__mux2i_1 _24040_ (.A0(_09919_),
    .A1(_09924_),
    .S(net297),
    .Y(_09925_));
 sky130_fd_sc_hd__nand2_2 _24041_ (.A(net357),
    .B(\w[1][2] ),
    .Y(_09926_));
 sky130_fd_sc_hd__o21ai_4 _24042_ (.A1(net292),
    .A2(_09925_),
    .B1(_09926_),
    .Y(_00054_));
 sky130_fd_sc_hd__mux4_2 _24043_ (.A0(\w[19][3] ),
    .A1(\w[17][3] ),
    .A2(\w[23][3] ),
    .A3(\w[21][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09927_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_560 ();
 sky130_fd_sc_hd__mux4_2 _24045_ (.A0(\w[27][3] ),
    .A1(\w[25][3] ),
    .A2(\w[31][3] ),
    .A3(\w[29][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09929_));
 sky130_fd_sc_hd__mux4_2 _24046_ (.A0(\w[3][3] ),
    .A1(\w[1][3] ),
    .A2(\w[7][3] ),
    .A3(\w[5][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09930_));
 sky130_fd_sc_hd__mux4_2 _24047_ (.A0(\w[11][3] ),
    .A1(\w[9][3] ),
    .A2(\w[15][3] ),
    .A3(\w[13][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09931_));
 sky130_fd_sc_hd__mux4_2 _24048_ (.A0(_09927_),
    .A1(_09929_),
    .A2(_09930_),
    .A3(_09931_),
    .S0(net343),
    .S1(net334),
    .X(_09932_));
 sky130_fd_sc_hd__mux4_2 _24049_ (.A0(\w[51][3] ),
    .A1(\w[49][3] ),
    .A2(\w[55][3] ),
    .A3(\w[53][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09933_));
 sky130_fd_sc_hd__mux4_2 _24050_ (.A0(\w[59][3] ),
    .A1(\w[57][3] ),
    .A2(\w[63][3] ),
    .A3(\w[61][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09934_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_559 ();
 sky130_fd_sc_hd__mux4_2 _24052_ (.A0(\w[35][3] ),
    .A1(\w[33][3] ),
    .A2(\w[39][3] ),
    .A3(\w[37][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09936_));
 sky130_fd_sc_hd__mux4_2 _24053_ (.A0(\w[43][3] ),
    .A1(\w[41][3] ),
    .A2(\w[47][3] ),
    .A3(\w[45][3] ),
    .S0(net367),
    .S1(net316),
    .X(_09937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_558 ();
 sky130_fd_sc_hd__mux4_2 _24055_ (.A0(_09933_),
    .A1(_09934_),
    .A2(_09936_),
    .A3(_09937_),
    .S0(net342),
    .S1(net336),
    .X(_09939_));
 sky130_fd_sc_hd__mux2i_1 _24056_ (.A0(_09932_),
    .A1(_09939_),
    .S(net297),
    .Y(_09940_));
 sky130_fd_sc_hd__nand2_2 _24057_ (.A(net357),
    .B(\w[1][3] ),
    .Y(_09941_));
 sky130_fd_sc_hd__o21ai_4 _24058_ (.A1(net292),
    .A2(_09940_),
    .B1(_09941_),
    .Y(_00057_));
 sky130_fd_sc_hd__mux4_2 _24059_ (.A0(\w[19][4] ),
    .A1(\w[17][4] ),
    .A2(\w[23][4] ),
    .A3(\w[21][4] ),
    .S0(net368),
    .S1(net314),
    .X(_09942_));
 sky130_fd_sc_hd__mux4_2 _24060_ (.A0(\w[27][4] ),
    .A1(\w[25][4] ),
    .A2(\w[31][4] ),
    .A3(\w[29][4] ),
    .S0(net368),
    .S1(net314),
    .X(_09943_));
 sky130_fd_sc_hd__mux4_2 _24061_ (.A0(\w[3][4] ),
    .A1(\w[1][4] ),
    .A2(\w[7][4] ),
    .A3(\w[5][4] ),
    .S0(net368),
    .S1(net314),
    .X(_09944_));
 sky130_fd_sc_hd__mux4_2 _24062_ (.A0(\w[11][4] ),
    .A1(\w[9][4] ),
    .A2(\w[15][4] ),
    .A3(\w[13][4] ),
    .S0(net368),
    .S1(net314),
    .X(_09945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_557 ();
 sky130_fd_sc_hd__mux4_2 _24064_ (.A0(_09942_),
    .A1(_09943_),
    .A2(_09944_),
    .A3(_09945_),
    .S0(net343),
    .S1(net334),
    .X(_09947_));
 sky130_fd_sc_hd__mux4_2 _24065_ (.A0(\w[51][4] ),
    .A1(\w[49][4] ),
    .A2(\w[55][4] ),
    .A3(\w[53][4] ),
    .S0(net367),
    .S1(net316),
    .X(_09948_));
 sky130_fd_sc_hd__mux4_2 _24066_ (.A0(\w[59][4] ),
    .A1(\w[57][4] ),
    .A2(\w[63][4] ),
    .A3(\w[61][4] ),
    .S0(net367),
    .S1(net316),
    .X(_09949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_556 ();
 sky130_fd_sc_hd__mux4_2 _24068_ (.A0(\w[35][4] ),
    .A1(\w[33][4] ),
    .A2(\w[39][4] ),
    .A3(\w[37][4] ),
    .S0(net367),
    .S1(net316),
    .X(_09951_));
 sky130_fd_sc_hd__mux4_2 _24069_ (.A0(\w[43][4] ),
    .A1(\w[41][4] ),
    .A2(\w[47][4] ),
    .A3(\w[45][4] ),
    .S0(net367),
    .S1(net316),
    .X(_09952_));
 sky130_fd_sc_hd__mux4_2 _24070_ (.A0(_09948_),
    .A1(_09949_),
    .A2(_09951_),
    .A3(_09952_),
    .S0(net346),
    .S1(net337),
    .X(_09953_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_553 ();
 sky130_fd_sc_hd__mux2i_1 _24074_ (.A0(_09947_),
    .A1(_09953_),
    .S(net297),
    .Y(_09957_));
 sky130_fd_sc_hd__nand2_2 _24075_ (.A(net357),
    .B(\w[1][4] ),
    .Y(_09958_));
 sky130_fd_sc_hd__o21ai_4 _24076_ (.A1(net292),
    .A2(_09957_),
    .B1(_09958_),
    .Y(_00058_));
 sky130_fd_sc_hd__mux4_2 _24077_ (.A0(\w[19][5] ),
    .A1(\w[17][5] ),
    .A2(\w[23][5] ),
    .A3(\w[21][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09959_));
 sky130_fd_sc_hd__mux4_2 _24078_ (.A0(\w[27][5] ),
    .A1(\w[25][5] ),
    .A2(\w[31][5] ),
    .A3(\w[29][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09960_));
 sky130_fd_sc_hd__mux4_2 _24079_ (.A0(\w[3][5] ),
    .A1(\w[1][5] ),
    .A2(\w[7][5] ),
    .A3(\w[5][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09961_));
 sky130_fd_sc_hd__mux4_2 _24080_ (.A0(\w[11][5] ),
    .A1(\w[9][5] ),
    .A2(\w[15][5] ),
    .A3(\w[13][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09962_));
 sky130_fd_sc_hd__mux4_2 _24081_ (.A0(_09959_),
    .A1(_09960_),
    .A2(_09961_),
    .A3(_09962_),
    .S0(net342),
    .S1(net336),
    .X(_09963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_552 ();
 sky130_fd_sc_hd__mux4_2 _24083_ (.A0(\w[51][5] ),
    .A1(\w[49][5] ),
    .A2(\w[55][5] ),
    .A3(\w[53][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09965_));
 sky130_fd_sc_hd__mux4_2 _24084_ (.A0(\w[59][5] ),
    .A1(\w[57][5] ),
    .A2(\w[63][5] ),
    .A3(\w[61][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09966_));
 sky130_fd_sc_hd__mux4_2 _24085_ (.A0(\w[35][5] ),
    .A1(\w[33][5] ),
    .A2(\w[39][5] ),
    .A3(\w[37][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09967_));
 sky130_fd_sc_hd__mux4_2 _24086_ (.A0(\w[43][5] ),
    .A1(\w[41][5] ),
    .A2(\w[47][5] ),
    .A3(\w[45][5] ),
    .S0(net367),
    .S1(net316),
    .X(_09968_));
 sky130_fd_sc_hd__mux4_2 _24087_ (.A0(_09965_),
    .A1(_09966_),
    .A2(_09967_),
    .A3(_09968_),
    .S0(net342),
    .S1(net336),
    .X(_09969_));
 sky130_fd_sc_hd__mux2i_1 _24088_ (.A0(_09963_),
    .A1(_09969_),
    .S(net297),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_2 _24089_ (.A(net357),
    .B(\w[1][5] ),
    .Y(_09971_));
 sky130_fd_sc_hd__o21ai_4 _24090_ (.A1(net292),
    .A2(_09970_),
    .B1(_09971_),
    .Y(_00059_));
 sky130_fd_sc_hd__mux4_2 _24091_ (.A0(\w[19][6] ),
    .A1(\w[17][6] ),
    .A2(\w[23][6] ),
    .A3(\w[21][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09972_));
 sky130_fd_sc_hd__mux4_2 _24092_ (.A0(\w[27][6] ),
    .A1(\w[25][6] ),
    .A2(\w[31][6] ),
    .A3(\w[29][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_551 ();
 sky130_fd_sc_hd__mux4_2 _24094_ (.A0(\w[3][6] ),
    .A1(\w[1][6] ),
    .A2(\w[7][6] ),
    .A3(\w[5][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09975_));
 sky130_fd_sc_hd__mux4_2 _24095_ (.A0(\w[11][6] ),
    .A1(\w[9][6] ),
    .A2(\w[15][6] ),
    .A3(\w[13][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09976_));
 sky130_fd_sc_hd__mux4_2 _24096_ (.A0(_09972_),
    .A1(_09973_),
    .A2(_09975_),
    .A3(_09976_),
    .S0(net341),
    .S1(net340),
    .X(_09977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_550 ();
 sky130_fd_sc_hd__mux4_2 _24098_ (.A0(\w[51][6] ),
    .A1(\w[49][6] ),
    .A2(\w[55][6] ),
    .A3(\w[53][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09979_));
 sky130_fd_sc_hd__mux4_2 _24099_ (.A0(\w[59][6] ),
    .A1(\w[57][6] ),
    .A2(\w[63][6] ),
    .A3(\w[61][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09980_));
 sky130_fd_sc_hd__mux4_2 _24100_ (.A0(\w[35][6] ),
    .A1(\w[33][6] ),
    .A2(\w[39][6] ),
    .A3(\w[37][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09981_));
 sky130_fd_sc_hd__mux4_2 _24101_ (.A0(\w[43][6] ),
    .A1(\w[41][6] ),
    .A2(\w[47][6] ),
    .A3(\w[45][6] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09982_));
 sky130_fd_sc_hd__mux4_2 _24102_ (.A0(_09979_),
    .A1(_09980_),
    .A2(_09981_),
    .A3(_09982_),
    .S0(net341),
    .S1(net340),
    .X(_09983_));
 sky130_fd_sc_hd__mux2i_1 _24103_ (.A0(_09977_),
    .A1(_09983_),
    .S(net299),
    .Y(_09984_));
 sky130_fd_sc_hd__nand2_2 _24104_ (.A(net357),
    .B(\w[1][6] ),
    .Y(_09985_));
 sky130_fd_sc_hd__o21ai_4 _24105_ (.A1(net291),
    .A2(_09984_),
    .B1(_09985_),
    .Y(_00060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_549 ();
 sky130_fd_sc_hd__mux4_2 _24107_ (.A0(\w[19][7] ),
    .A1(\w[17][7] ),
    .A2(\w[23][7] ),
    .A3(\w[21][7] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09987_));
 sky130_fd_sc_hd__mux4_2 _24108_ (.A0(\w[27][7] ),
    .A1(\w[25][7] ),
    .A2(\w[31][7] ),
    .A3(\w[29][7] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09988_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_548 ();
 sky130_fd_sc_hd__mux4_2 _24110_ (.A0(\w[3][7] ),
    .A1(\w[1][7] ),
    .A2(\w[7][7] ),
    .A3(\w[5][7] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09990_));
 sky130_fd_sc_hd__mux4_2 _24111_ (.A0(\w[11][7] ),
    .A1(\w[9][7] ),
    .A2(\w[15][7] ),
    .A3(\w[13][7] ),
    .S0(net366),
    .S1(_00657_),
    .X(_09991_));
 sky130_fd_sc_hd__mux4_2 _24112_ (.A0(_09987_),
    .A1(_09988_),
    .A2(_09990_),
    .A3(_09991_),
    .S0(net341),
    .S1(net340),
    .X(_09992_));
 sky130_fd_sc_hd__mux4_2 _24113_ (.A0(\w[51][7] ),
    .A1(\w[49][7] ),
    .A2(\w[55][7] ),
    .A3(\w[53][7] ),
    .S0(net366),
    .S1(net313),
    .X(_09993_));
 sky130_fd_sc_hd__mux4_2 _24114_ (.A0(\w[59][7] ),
    .A1(\w[57][7] ),
    .A2(\w[63][7] ),
    .A3(\w[61][7] ),
    .S0(net366),
    .S1(net313),
    .X(_09994_));
 sky130_fd_sc_hd__mux4_2 _24115_ (.A0(\w[35][7] ),
    .A1(\w[33][7] ),
    .A2(\w[39][7] ),
    .A3(\w[37][7] ),
    .S0(net366),
    .S1(net313),
    .X(_09995_));
 sky130_fd_sc_hd__mux4_2 _24116_ (.A0(\w[43][7] ),
    .A1(\w[41][7] ),
    .A2(\w[47][7] ),
    .A3(\w[45][7] ),
    .S0(net366),
    .S1(net313),
    .X(_09996_));
 sky130_fd_sc_hd__mux4_2 _24117_ (.A0(_09993_),
    .A1(_09994_),
    .A2(_09995_),
    .A3(_09996_),
    .S0(net341),
    .S1(net338),
    .X(_09997_));
 sky130_fd_sc_hd__mux2i_1 _24118_ (.A0(_09992_),
    .A1(_09997_),
    .S(net299),
    .Y(_09998_));
 sky130_fd_sc_hd__nand2_2 _24119_ (.A(net357),
    .B(\w[1][7] ),
    .Y(_09999_));
 sky130_fd_sc_hd__o21ai_4 _24120_ (.A1(net291),
    .A2(_09998_),
    .B1(_09999_),
    .Y(_00061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_547 ();
 sky130_fd_sc_hd__mux4_2 _24122_ (.A0(\w[19][8] ),
    .A1(\w[17][8] ),
    .A2(\w[23][8] ),
    .A3(\w[21][8] ),
    .S0(net368),
    .S1(net314),
    .X(_10001_));
 sky130_fd_sc_hd__mux4_2 _24123_ (.A0(\w[27][8] ),
    .A1(\w[25][8] ),
    .A2(\w[31][8] ),
    .A3(\w[29][8] ),
    .S0(net368),
    .S1(net314),
    .X(_10002_));
 sky130_fd_sc_hd__mux4_2 _24124_ (.A0(\w[3][8] ),
    .A1(\w[1][8] ),
    .A2(\w[7][8] ),
    .A3(\w[5][8] ),
    .S0(net368),
    .S1(net314),
    .X(_10003_));
 sky130_fd_sc_hd__mux4_2 _24125_ (.A0(\w[11][8] ),
    .A1(\w[9][8] ),
    .A2(\w[15][8] ),
    .A3(\w[13][8] ),
    .S0(net368),
    .S1(net314),
    .X(_10004_));
 sky130_fd_sc_hd__mux4_2 _24126_ (.A0(_10001_),
    .A1(_10002_),
    .A2(_10003_),
    .A3(_10004_),
    .S0(net343),
    .S1(net334),
    .X(_10005_));
 sky130_fd_sc_hd__mux4_2 _24127_ (.A0(\w[51][8] ),
    .A1(\w[49][8] ),
    .A2(\w[55][8] ),
    .A3(\w[53][8] ),
    .S0(net372),
    .S1(net316),
    .X(_10006_));
 sky130_fd_sc_hd__mux4_2 _24128_ (.A0(\w[59][8] ),
    .A1(\w[57][8] ),
    .A2(\w[63][8] ),
    .A3(\w[61][8] ),
    .S0(net372),
    .S1(net316),
    .X(_10007_));
 sky130_fd_sc_hd__mux4_2 _24129_ (.A0(\w[35][8] ),
    .A1(\w[33][8] ),
    .A2(\w[39][8] ),
    .A3(\w[37][8] ),
    .S0(net372),
    .S1(net316),
    .X(_10008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_546 ();
 sky130_fd_sc_hd__mux4_2 _24131_ (.A0(\w[43][8] ),
    .A1(\w[41][8] ),
    .A2(\w[47][8] ),
    .A3(\w[45][8] ),
    .S0(net372),
    .S1(net316),
    .X(_10010_));
 sky130_fd_sc_hd__mux4_2 _24132_ (.A0(_10006_),
    .A1(_10007_),
    .A2(_10008_),
    .A3(_10010_),
    .S0(net346),
    .S1(net338),
    .X(_10011_));
 sky130_fd_sc_hd__mux2i_1 _24133_ (.A0(_10005_),
    .A1(_10011_),
    .S(net297),
    .Y(_10012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_544 ();
 sky130_fd_sc_hd__nand2_2 _24136_ (.A(net357),
    .B(\w[1][8] ),
    .Y(_10015_));
 sky130_fd_sc_hd__o21ai_4 _24137_ (.A1(net292),
    .A2(_10012_),
    .B1(_10015_),
    .Y(_00062_));
 sky130_fd_sc_hd__mux4_2 _24138_ (.A0(\w[19][9] ),
    .A1(\w[17][9] ),
    .A2(\w[23][9] ),
    .A3(\w[21][9] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10016_));
 sky130_fd_sc_hd__mux4_2 _24139_ (.A0(\w[27][9] ),
    .A1(\w[25][9] ),
    .A2(\w[31][9] ),
    .A3(\w[29][9] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10017_));
 sky130_fd_sc_hd__mux4_2 _24140_ (.A0(\w[3][9] ),
    .A1(\w[1][9] ),
    .A2(\w[7][9] ),
    .A3(\w[5][9] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10018_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_543 ();
 sky130_fd_sc_hd__mux4_2 _24142_ (.A0(\w[11][9] ),
    .A1(\w[9][9] ),
    .A2(\w[15][9] ),
    .A3(\w[13][9] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10020_));
 sky130_fd_sc_hd__mux4_2 _24143_ (.A0(_10016_),
    .A1(_10017_),
    .A2(_10018_),
    .A3(_10020_),
    .S0(net347),
    .S1(net340),
    .X(_10021_));
 sky130_fd_sc_hd__mux4_2 _24144_ (.A0(\w[51][9] ),
    .A1(\w[49][9] ),
    .A2(\w[55][9] ),
    .A3(\w[53][9] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_542 ();
 sky130_fd_sc_hd__mux4_2 _24146_ (.A0(\w[59][9] ),
    .A1(\w[57][9] ),
    .A2(\w[63][9] ),
    .A3(\w[61][9] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10024_));
 sky130_fd_sc_hd__mux4_2 _24147_ (.A0(\w[35][9] ),
    .A1(\w[33][9] ),
    .A2(\w[39][9] ),
    .A3(\w[37][9] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_541 ();
 sky130_fd_sc_hd__mux4_2 _24149_ (.A0(\w[43][9] ),
    .A1(\w[41][9] ),
    .A2(\w[47][9] ),
    .A3(\w[45][9] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10027_));
 sky130_fd_sc_hd__mux4_2 _24150_ (.A0(_10022_),
    .A1(_10024_),
    .A2(_10025_),
    .A3(_10027_),
    .S0(_09854_),
    .S1(net340),
    .X(_10028_));
 sky130_fd_sc_hd__mux2i_1 _24151_ (.A0(_10021_),
    .A1(_10028_),
    .S(net299),
    .Y(_10029_));
 sky130_fd_sc_hd__nand2_1 _24152_ (.A(net540),
    .B(\w[1][9] ),
    .Y(_10030_));
 sky130_fd_sc_hd__o21ai_1 _24153_ (.A1(net292),
    .A2(_10029_),
    .B1(_10030_),
    .Y(_00063_));
 sky130_fd_sc_hd__mux4_2 _24154_ (.A0(\w[19][10] ),
    .A1(\w[17][10] ),
    .A2(\w[23][10] ),
    .A3(\w[21][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10031_));
 sky130_fd_sc_hd__mux4_2 _24155_ (.A0(\w[27][10] ),
    .A1(\w[25][10] ),
    .A2(\w[31][10] ),
    .A3(\w[29][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10032_));
 sky130_fd_sc_hd__mux4_2 _24156_ (.A0(\w[3][10] ),
    .A1(\w[1][10] ),
    .A2(\w[7][10] ),
    .A3(\w[5][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10033_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_540 ();
 sky130_fd_sc_hd__mux4_2 _24158_ (.A0(\w[11][10] ),
    .A1(\w[9][10] ),
    .A2(\w[15][10] ),
    .A3(\w[13][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10035_));
 sky130_fd_sc_hd__mux4_2 _24159_ (.A0(_10031_),
    .A1(_10032_),
    .A2(_10033_),
    .A3(_10035_),
    .S0(net345),
    .S1(net335),
    .X(_10036_));
 sky130_fd_sc_hd__mux4_2 _24160_ (.A0(\w[51][10] ),
    .A1(\w[49][10] ),
    .A2(\w[55][10] ),
    .A3(\w[53][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_539 ();
 sky130_fd_sc_hd__mux4_2 _24162_ (.A0(\w[59][10] ),
    .A1(\w[57][10] ),
    .A2(\w[63][10] ),
    .A3(\w[61][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10039_));
 sky130_fd_sc_hd__mux4_2 _24163_ (.A0(\w[35][10] ),
    .A1(\w[33][10] ),
    .A2(\w[39][10] ),
    .A3(\w[37][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10040_));
 sky130_fd_sc_hd__mux4_2 _24164_ (.A0(\w[43][10] ),
    .A1(\w[41][10] ),
    .A2(\w[47][10] ),
    .A3(\w[45][10] ),
    .S0(net371),
    .S1(net318),
    .X(_10041_));
 sky130_fd_sc_hd__mux4_2 _24165_ (.A0(_10037_),
    .A1(_10039_),
    .A2(_10040_),
    .A3(_10041_),
    .S0(net346),
    .S1(_09857_),
    .X(_10042_));
 sky130_fd_sc_hd__mux2i_1 _24166_ (.A0(_10036_),
    .A1(_10042_),
    .S(net298),
    .Y(_10043_));
 sky130_fd_sc_hd__nand2_1 _24167_ (.A(net357),
    .B(\w[1][10] ),
    .Y(_10044_));
 sky130_fd_sc_hd__o21ai_0 _24168_ (.A1(net292),
    .A2(_10043_),
    .B1(_10044_),
    .Y(_00033_));
 sky130_fd_sc_hd__mux4_2 _24169_ (.A0(\w[19][11] ),
    .A1(\w[17][11] ),
    .A2(\w[23][11] ),
    .A3(\w[21][11] ),
    .S0(net370),
    .S1(net317),
    .X(_10045_));
 sky130_fd_sc_hd__mux4_2 _24170_ (.A0(\w[27][11] ),
    .A1(\w[25][11] ),
    .A2(\w[31][11] ),
    .A3(\w[29][11] ),
    .S0(net370),
    .S1(net317),
    .X(_10046_));
 sky130_fd_sc_hd__mux4_2 _24171_ (.A0(\w[3][11] ),
    .A1(\w[1][11] ),
    .A2(\w[7][11] ),
    .A3(\w[5][11] ),
    .S0(net370),
    .S1(net317),
    .X(_10047_));
 sky130_fd_sc_hd__mux4_2 _24172_ (.A0(\w[11][11] ),
    .A1(\w[9][11] ),
    .A2(\w[15][11] ),
    .A3(\w[13][11] ),
    .S0(net370),
    .S1(net317),
    .X(_10048_));
 sky130_fd_sc_hd__mux4_2 _24173_ (.A0(_10045_),
    .A1(_10046_),
    .A2(_10047_),
    .A3(_10048_),
    .S0(net344),
    .S1(net335),
    .X(_10049_));
 sky130_fd_sc_hd__mux4_2 _24174_ (.A0(\w[51][11] ),
    .A1(\w[49][11] ),
    .A2(\w[55][11] ),
    .A3(\w[53][11] ),
    .S0(net372),
    .S1(net318),
    .X(_10050_));
 sky130_fd_sc_hd__mux4_2 _24175_ (.A0(\w[59][11] ),
    .A1(\w[57][11] ),
    .A2(\w[63][11] ),
    .A3(\w[61][11] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10051_));
 sky130_fd_sc_hd__mux4_2 _24176_ (.A0(\w[35][11] ),
    .A1(\w[33][11] ),
    .A2(\w[39][11] ),
    .A3(\w[37][11] ),
    .S0(net372),
    .S1(net318),
    .X(_10052_));
 sky130_fd_sc_hd__mux4_2 _24177_ (.A0(\w[43][11] ),
    .A1(\w[41][11] ),
    .A2(\w[47][11] ),
    .A3(\w[45][11] ),
    .S0(net372),
    .S1(net318),
    .X(_10053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_538 ();
 sky130_fd_sc_hd__mux4_2 _24179_ (.A0(_10050_),
    .A1(_10051_),
    .A2(_10052_),
    .A3(_10053_),
    .S0(net347),
    .S1(net338),
    .X(_10055_));
 sky130_fd_sc_hd__mux2i_1 _24180_ (.A0(_10049_),
    .A1(_10055_),
    .S(net297),
    .Y(_10056_));
 sky130_fd_sc_hd__nand2_1 _24181_ (.A(net357),
    .B(\w[1][11] ),
    .Y(_10057_));
 sky130_fd_sc_hd__o21ai_2 _24182_ (.A1(net292),
    .A2(_10056_),
    .B1(_10057_),
    .Y(_00034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_537 ();
 sky130_fd_sc_hd__mux4_2 _24184_ (.A0(\w[19][12] ),
    .A1(\w[17][12] ),
    .A2(\w[23][12] ),
    .A3(\w[21][12] ),
    .S0(net370),
    .S1(net317),
    .X(_10059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_536 ();
 sky130_fd_sc_hd__mux4_2 _24186_ (.A0(\w[27][12] ),
    .A1(\w[25][12] ),
    .A2(\w[31][12] ),
    .A3(\w[29][12] ),
    .S0(net370),
    .S1(net317),
    .X(_10061_));
 sky130_fd_sc_hd__mux4_2 _24187_ (.A0(\w[3][12] ),
    .A1(\w[1][12] ),
    .A2(\w[7][12] ),
    .A3(\w[5][12] ),
    .S0(net370),
    .S1(net317),
    .X(_10062_));
 sky130_fd_sc_hd__mux4_2 _24188_ (.A0(\w[11][12] ),
    .A1(\w[9][12] ),
    .A2(\w[15][12] ),
    .A3(\w[13][12] ),
    .S0(net370),
    .S1(net317),
    .X(_10063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_535 ();
 sky130_fd_sc_hd__mux4_2 _24190_ (.A0(_10059_),
    .A1(_10061_),
    .A2(_10062_),
    .A3(_10063_),
    .S0(net344),
    .S1(net334),
    .X(_10065_));
 sky130_fd_sc_hd__mux4_2 _24191_ (.A0(\w[51][12] ),
    .A1(\w[49][12] ),
    .A2(\w[55][12] ),
    .A3(\w[53][12] ),
    .S0(net372),
    .S1(net316),
    .X(_10066_));
 sky130_fd_sc_hd__mux4_2 _24192_ (.A0(\w[59][12] ),
    .A1(\w[57][12] ),
    .A2(\w[63][12] ),
    .A3(\w[61][12] ),
    .S0(net372),
    .S1(net316),
    .X(_10067_));
 sky130_fd_sc_hd__mux4_2 _24193_ (.A0(\w[35][12] ),
    .A1(\w[33][12] ),
    .A2(\w[39][12] ),
    .A3(\w[37][12] ),
    .S0(net372),
    .S1(net316),
    .X(_10068_));
 sky130_fd_sc_hd__mux4_2 _24194_ (.A0(\w[43][12] ),
    .A1(\w[41][12] ),
    .A2(\w[47][12] ),
    .A3(\w[45][12] ),
    .S0(net372),
    .S1(net316),
    .X(_10069_));
 sky130_fd_sc_hd__mux4_2 _24195_ (.A0(_10066_),
    .A1(_10067_),
    .A2(_10068_),
    .A3(_10069_),
    .S0(net346),
    .S1(net338),
    .X(_10070_));
 sky130_fd_sc_hd__mux2i_1 _24196_ (.A0(_10065_),
    .A1(_10070_),
    .S(net297),
    .Y(_10071_));
 sky130_fd_sc_hd__nand2_2 _24197_ (.A(net357),
    .B(\w[1][12] ),
    .Y(_10072_));
 sky130_fd_sc_hd__o21ai_4 _24198_ (.A1(net292),
    .A2(_10071_),
    .B1(_10072_),
    .Y(_00035_));
 sky130_fd_sc_hd__mux4_2 _24199_ (.A0(\w[19][13] ),
    .A1(\w[17][13] ),
    .A2(\w[23][13] ),
    .A3(\w[21][13] ),
    .S0(net371),
    .S1(net318),
    .X(_10073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_534 ();
 sky130_fd_sc_hd__mux4_2 _24201_ (.A0(\w[27][13] ),
    .A1(\w[25][13] ),
    .A2(\w[31][13] ),
    .A3(\w[29][13] ),
    .S0(net371),
    .S1(net318),
    .X(_10075_));
 sky130_fd_sc_hd__mux4_2 _24202_ (.A0(\w[3][13] ),
    .A1(\w[1][13] ),
    .A2(\w[7][13] ),
    .A3(\w[5][13] ),
    .S0(net371),
    .S1(net318),
    .X(_10076_));
 sky130_fd_sc_hd__mux4_2 _24203_ (.A0(\w[11][13] ),
    .A1(\w[9][13] ),
    .A2(\w[15][13] ),
    .A3(\w[13][13] ),
    .S0(net371),
    .S1(net318),
    .X(_10077_));
 sky130_fd_sc_hd__mux4_2 _24204_ (.A0(_10073_),
    .A1(_10075_),
    .A2(_10076_),
    .A3(_10077_),
    .S0(net345),
    .S1(net335),
    .X(_10078_));
 sky130_fd_sc_hd__mux4_2 _24205_ (.A0(\w[51][13] ),
    .A1(\w[49][13] ),
    .A2(\w[55][13] ),
    .A3(\w[53][13] ),
    .S0(net372),
    .S1(net317),
    .X(_10079_));
 sky130_fd_sc_hd__mux4_2 _24206_ (.A0(\w[59][13] ),
    .A1(\w[57][13] ),
    .A2(\w[63][13] ),
    .A3(\w[61][13] ),
    .S0(net372),
    .S1(net318),
    .X(_10080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_533 ();
 sky130_fd_sc_hd__mux4_2 _24208_ (.A0(\w[35][13] ),
    .A1(\w[33][13] ),
    .A2(\w[39][13] ),
    .A3(\w[37][13] ),
    .S0(net371),
    .S1(net318),
    .X(_10082_));
 sky130_fd_sc_hd__mux4_2 _24209_ (.A0(\w[43][13] ),
    .A1(\w[41][13] ),
    .A2(\w[47][13] ),
    .A3(\w[45][13] ),
    .S0(net372),
    .S1(net317),
    .X(_10083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_532 ();
 sky130_fd_sc_hd__mux4_2 _24211_ (.A0(_10079_),
    .A1(_10080_),
    .A2(_10082_),
    .A3(_10083_),
    .S0(net347),
    .S1(net338),
    .X(_10085_));
 sky130_fd_sc_hd__mux2i_1 _24212_ (.A0(_10078_),
    .A1(_10085_),
    .S(net298),
    .Y(_10086_));
 sky130_fd_sc_hd__nand2_1 _24213_ (.A(net357),
    .B(\w[1][13] ),
    .Y(_10087_));
 sky130_fd_sc_hd__o21ai_0 _24214_ (.A1(net292),
    .A2(_10086_),
    .B1(_10087_),
    .Y(_00036_));
 sky130_fd_sc_hd__mux4_2 _24215_ (.A0(\w[19][14] ),
    .A1(\w[17][14] ),
    .A2(\w[23][14] ),
    .A3(\w[21][14] ),
    .S0(net370),
    .S1(net317),
    .X(_10088_));
 sky130_fd_sc_hd__mux4_2 _24216_ (.A0(\w[27][14] ),
    .A1(\w[25][14] ),
    .A2(\w[31][14] ),
    .A3(\w[29][14] ),
    .S0(net370),
    .S1(net317),
    .X(_10089_));
 sky130_fd_sc_hd__mux4_2 _24217_ (.A0(\w[3][14] ),
    .A1(\w[1][14] ),
    .A2(\w[7][14] ),
    .A3(\w[5][14] ),
    .S0(net370),
    .S1(net317),
    .X(_10090_));
 sky130_fd_sc_hd__mux4_2 _24218_ (.A0(\w[11][14] ),
    .A1(\w[9][14] ),
    .A2(\w[15][14] ),
    .A3(\w[13][14] ),
    .S0(net370),
    .S1(net317),
    .X(_10091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_531 ();
 sky130_fd_sc_hd__mux4_2 _24220_ (.A0(_10088_),
    .A1(_10089_),
    .A2(_10090_),
    .A3(_10091_),
    .S0(net344),
    .S1(net335),
    .X(_10093_));
 sky130_fd_sc_hd__mux4_2 _24221_ (.A0(\w[51][14] ),
    .A1(\w[49][14] ),
    .A2(\w[55][14] ),
    .A3(\w[53][14] ),
    .S0(net368),
    .S1(net314),
    .X(_10094_));
 sky130_fd_sc_hd__mux4_2 _24222_ (.A0(\w[59][14] ),
    .A1(\w[57][14] ),
    .A2(\w[63][14] ),
    .A3(\w[61][14] ),
    .S0(net368),
    .S1(net314),
    .X(_10095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_530 ();
 sky130_fd_sc_hd__mux4_2 _24224_ (.A0(\w[35][14] ),
    .A1(\w[33][14] ),
    .A2(\w[39][14] ),
    .A3(\w[37][14] ),
    .S0(net368),
    .S1(net314),
    .X(_10097_));
 sky130_fd_sc_hd__mux4_2 _24225_ (.A0(\w[43][14] ),
    .A1(\w[41][14] ),
    .A2(\w[47][14] ),
    .A3(\w[45][14] ),
    .S0(net368),
    .S1(net314),
    .X(_10098_));
 sky130_fd_sc_hd__mux4_2 _24226_ (.A0(_10094_),
    .A1(_10095_),
    .A2(_10097_),
    .A3(_10098_),
    .S0(net343),
    .S1(net334),
    .X(_10099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_529 ();
 sky130_fd_sc_hd__mux2i_1 _24228_ (.A0(_10093_),
    .A1(_10099_),
    .S(net297),
    .Y(_10101_));
 sky130_fd_sc_hd__nand2_2 _24229_ (.A(net357),
    .B(\w[1][14] ),
    .Y(_10102_));
 sky130_fd_sc_hd__o21ai_4 _24230_ (.A1(net292),
    .A2(_10101_),
    .B1(_10102_),
    .Y(_00037_));
 sky130_fd_sc_hd__mux4_2 _24231_ (.A0(\w[19][15] ),
    .A1(\w[17][15] ),
    .A2(\w[23][15] ),
    .A3(\w[21][15] ),
    .S0(net365),
    .S1(net313),
    .X(_10103_));
 sky130_fd_sc_hd__mux4_2 _24232_ (.A0(\w[27][15] ),
    .A1(\w[25][15] ),
    .A2(\w[31][15] ),
    .A3(\w[29][15] ),
    .S0(net365),
    .S1(net313),
    .X(_10104_));
 sky130_fd_sc_hd__mux4_2 _24233_ (.A0(\w[3][15] ),
    .A1(\w[1][15] ),
    .A2(\w[7][15] ),
    .A3(\w[5][15] ),
    .S0(net365),
    .S1(net313),
    .X(_10105_));
 sky130_fd_sc_hd__mux4_2 _24234_ (.A0(\w[11][15] ),
    .A1(\w[9][15] ),
    .A2(\w[15][15] ),
    .A3(\w[13][15] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10106_));
 sky130_fd_sc_hd__mux4_2 _24235_ (.A0(_10103_),
    .A1(_10104_),
    .A2(_10105_),
    .A3(_10106_),
    .S0(net341),
    .S1(net338),
    .X(_10107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_528 ();
 sky130_fd_sc_hd__mux4_2 _24237_ (.A0(\w[51][15] ),
    .A1(\w[49][15] ),
    .A2(\w[55][15] ),
    .A3(\w[53][15] ),
    .S0(net365),
    .S1(net313),
    .X(_10109_));
 sky130_fd_sc_hd__mux4_2 _24238_ (.A0(\w[59][15] ),
    .A1(\w[57][15] ),
    .A2(\w[63][15] ),
    .A3(\w[61][15] ),
    .S0(net365),
    .S1(net313),
    .X(_10110_));
 sky130_fd_sc_hd__mux4_2 _24239_ (.A0(\w[35][15] ),
    .A1(\w[33][15] ),
    .A2(\w[39][15] ),
    .A3(\w[37][15] ),
    .S0(net365),
    .S1(net313),
    .X(_10111_));
 sky130_fd_sc_hd__mux4_2 _24240_ (.A0(\w[43][15] ),
    .A1(\w[41][15] ),
    .A2(\w[47][15] ),
    .A3(\w[45][15] ),
    .S0(net365),
    .S1(net313),
    .X(_10112_));
 sky130_fd_sc_hd__mux4_2 _24241_ (.A0(_10109_),
    .A1(_10110_),
    .A2(_10111_),
    .A3(_10112_),
    .S0(net341),
    .S1(net338),
    .X(_10113_));
 sky130_fd_sc_hd__mux2i_1 _24242_ (.A0(_10107_),
    .A1(_10113_),
    .S(net299),
    .Y(_10114_));
 sky130_fd_sc_hd__nand2_2 _24243_ (.A(net357),
    .B(\w[1][15] ),
    .Y(_10115_));
 sky130_fd_sc_hd__o21ai_4 _24244_ (.A1(net291),
    .A2(_10114_),
    .B1(_10115_),
    .Y(_00038_));
 sky130_fd_sc_hd__mux4_2 _24245_ (.A0(\w[19][16] ),
    .A1(\w[17][16] ),
    .A2(\w[23][16] ),
    .A3(\w[21][16] ),
    .S0(net368),
    .S1(net314),
    .X(_10116_));
 sky130_fd_sc_hd__mux4_2 _24246_ (.A0(\w[27][16] ),
    .A1(\w[25][16] ),
    .A2(\w[31][16] ),
    .A3(\w[29][16] ),
    .S0(net368),
    .S1(net314),
    .X(_10117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_527 ();
 sky130_fd_sc_hd__mux4_2 _24248_ (.A0(\w[3][16] ),
    .A1(\w[1][16] ),
    .A2(\w[7][16] ),
    .A3(\w[5][16] ),
    .S0(net368),
    .S1(net314),
    .X(_10119_));
 sky130_fd_sc_hd__mux4_2 _24249_ (.A0(\w[11][16] ),
    .A1(\w[9][16] ),
    .A2(\w[15][16] ),
    .A3(\w[13][16] ),
    .S0(net368),
    .S1(net314),
    .X(_10120_));
 sky130_fd_sc_hd__mux4_2 _24250_ (.A0(_10116_),
    .A1(_10117_),
    .A2(_10119_),
    .A3(_10120_),
    .S0(net344),
    .S1(net335),
    .X(_10121_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_526 ();
 sky130_fd_sc_hd__mux4_2 _24252_ (.A0(\w[51][16] ),
    .A1(\w[49][16] ),
    .A2(\w[55][16] ),
    .A3(\w[53][16] ),
    .S0(net367),
    .S1(net316),
    .X(_10123_));
 sky130_fd_sc_hd__mux4_2 _24253_ (.A0(\w[59][16] ),
    .A1(\w[57][16] ),
    .A2(\w[63][16] ),
    .A3(\w[61][16] ),
    .S0(net367),
    .S1(net316),
    .X(_10124_));
 sky130_fd_sc_hd__mux4_2 _24254_ (.A0(\w[35][16] ),
    .A1(\w[33][16] ),
    .A2(\w[39][16] ),
    .A3(\w[37][16] ),
    .S0(net367),
    .S1(net316),
    .X(_10125_));
 sky130_fd_sc_hd__mux4_2 _24255_ (.A0(\w[43][16] ),
    .A1(\w[41][16] ),
    .A2(\w[47][16] ),
    .A3(\w[45][16] ),
    .S0(net367),
    .S1(net316),
    .X(_10126_));
 sky130_fd_sc_hd__mux4_2 _24256_ (.A0(_10123_),
    .A1(_10124_),
    .A2(_10125_),
    .A3(_10126_),
    .S0(net346),
    .S1(net337),
    .X(_10127_));
 sky130_fd_sc_hd__mux2i_1 _24257_ (.A0(_10121_),
    .A1(_10127_),
    .S(net297),
    .Y(_10128_));
 sky130_fd_sc_hd__nand2_2 _24258_ (.A(net357),
    .B(\w[1][16] ),
    .Y(_10129_));
 sky130_fd_sc_hd__o21ai_4 _24259_ (.A1(net292),
    .A2(_10128_),
    .B1(_10129_),
    .Y(_00039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_525 ();
 sky130_fd_sc_hd__mux4_2 _24261_ (.A0(\w[19][17] ),
    .A1(\w[17][17] ),
    .A2(\w[23][17] ),
    .A3(\w[21][17] ),
    .S0(net369),
    .S1(net315),
    .X(_10131_));
 sky130_fd_sc_hd__mux4_2 _24262_ (.A0(\w[27][17] ),
    .A1(\w[25][17] ),
    .A2(\w[31][17] ),
    .A3(\w[29][17] ),
    .S0(net369),
    .S1(net315),
    .X(_10132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_524 ();
 sky130_fd_sc_hd__mux4_2 _24264_ (.A0(\w[3][17] ),
    .A1(\w[1][17] ),
    .A2(\w[7][17] ),
    .A3(\w[5][17] ),
    .S0(net369),
    .S1(net315),
    .X(_10134_));
 sky130_fd_sc_hd__mux4_2 _24265_ (.A0(\w[11][17] ),
    .A1(\w[9][17] ),
    .A2(\w[15][17] ),
    .A3(\w[13][17] ),
    .S0(net368),
    .S1(net314),
    .X(_10135_));
 sky130_fd_sc_hd__mux4_2 _24266_ (.A0(_10131_),
    .A1(_10132_),
    .A2(_10134_),
    .A3(_10135_),
    .S0(net343),
    .S1(net337),
    .X(_10136_));
 sky130_fd_sc_hd__mux4_2 _24267_ (.A0(\w[51][17] ),
    .A1(\w[49][17] ),
    .A2(\w[55][17] ),
    .A3(\w[53][17] ),
    .S0(net367),
    .S1(net316),
    .X(_10137_));
 sky130_fd_sc_hd__mux4_2 _24268_ (.A0(\w[59][17] ),
    .A1(\w[57][17] ),
    .A2(\w[63][17] ),
    .A3(\w[61][17] ),
    .S0(net367),
    .S1(net316),
    .X(_10138_));
 sky130_fd_sc_hd__mux4_2 _24269_ (.A0(\w[35][17] ),
    .A1(\w[33][17] ),
    .A2(\w[39][17] ),
    .A3(\w[37][17] ),
    .S0(net367),
    .S1(net316),
    .X(_10139_));
 sky130_fd_sc_hd__mux4_2 _24270_ (.A0(\w[43][17] ),
    .A1(\w[41][17] ),
    .A2(\w[47][17] ),
    .A3(\w[45][17] ),
    .S0(net367),
    .S1(net316),
    .X(_10140_));
 sky130_fd_sc_hd__mux4_2 _24271_ (.A0(_10137_),
    .A1(_10138_),
    .A2(_10139_),
    .A3(_10140_),
    .S0(net346),
    .S1(net337),
    .X(_10141_));
 sky130_fd_sc_hd__mux2i_1 _24272_ (.A0(_10136_),
    .A1(_10141_),
    .S(net297),
    .Y(_10142_));
 sky130_fd_sc_hd__nand2_2 _24273_ (.A(net357),
    .B(\w[1][17] ),
    .Y(_10143_));
 sky130_fd_sc_hd__o21ai_4 _24274_ (.A1(net292),
    .A2(_10142_),
    .B1(_10143_),
    .Y(_00040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_523 ();
 sky130_fd_sc_hd__mux4_2 _24276_ (.A0(\w[19][18] ),
    .A1(\w[17][18] ),
    .A2(\w[23][18] ),
    .A3(\w[21][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10145_));
 sky130_fd_sc_hd__mux4_2 _24277_ (.A0(\w[27][18] ),
    .A1(\w[25][18] ),
    .A2(\w[31][18] ),
    .A3(\w[29][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10146_));
 sky130_fd_sc_hd__mux4_2 _24278_ (.A0(\w[3][18] ),
    .A1(\w[1][18] ),
    .A2(\w[7][18] ),
    .A3(\w[5][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10147_));
 sky130_fd_sc_hd__mux4_2 _24279_ (.A0(\w[11][18] ),
    .A1(\w[9][18] ),
    .A2(\w[15][18] ),
    .A3(\w[13][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10148_));
 sky130_fd_sc_hd__mux4_2 _24280_ (.A0(_10145_),
    .A1(_10146_),
    .A2(_10147_),
    .A3(_10148_),
    .S0(net345),
    .S1(net335),
    .X(_10149_));
 sky130_fd_sc_hd__mux4_2 _24281_ (.A0(\w[51][18] ),
    .A1(\w[49][18] ),
    .A2(\w[55][18] ),
    .A3(\w[53][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10150_));
 sky130_fd_sc_hd__mux4_2 _24282_ (.A0(\w[59][18] ),
    .A1(\w[57][18] ),
    .A2(\w[63][18] ),
    .A3(\w[61][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10151_));
 sky130_fd_sc_hd__mux4_2 _24283_ (.A0(\w[35][18] ),
    .A1(\w[33][18] ),
    .A2(\w[39][18] ),
    .A3(\w[37][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_522 ();
 sky130_fd_sc_hd__mux4_2 _24285_ (.A0(\w[43][18] ),
    .A1(\w[41][18] ),
    .A2(\w[47][18] ),
    .A3(\w[45][18] ),
    .S0(net371),
    .S1(net318),
    .X(_10154_));
 sky130_fd_sc_hd__mux4_2 _24286_ (.A0(_10150_),
    .A1(_10151_),
    .A2(_10152_),
    .A3(_10154_),
    .S0(net344),
    .S1(net334),
    .X(_10155_));
 sky130_fd_sc_hd__mux2i_1 _24287_ (.A0(_10149_),
    .A1(_10155_),
    .S(net297),
    .Y(_10156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_521 ();
 sky130_fd_sc_hd__nand2_1 _24289_ (.A(net357),
    .B(\w[1][18] ),
    .Y(_10158_));
 sky130_fd_sc_hd__o21ai_0 _24290_ (.A1(net292),
    .A2(_10156_),
    .B1(_10158_),
    .Y(_00041_));
 sky130_fd_sc_hd__mux4_2 _24291_ (.A0(\w[19][19] ),
    .A1(\w[17][19] ),
    .A2(\w[23][19] ),
    .A3(\w[21][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10159_));
 sky130_fd_sc_hd__mux4_2 _24292_ (.A0(\w[27][19] ),
    .A1(\w[25][19] ),
    .A2(\w[31][19] ),
    .A3(\w[29][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10160_));
 sky130_fd_sc_hd__mux4_2 _24293_ (.A0(\w[3][19] ),
    .A1(\w[1][19] ),
    .A2(\w[7][19] ),
    .A3(\w[5][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_520 ();
 sky130_fd_sc_hd__mux4_2 _24295_ (.A0(\w[11][19] ),
    .A1(\w[9][19] ),
    .A2(\w[15][19] ),
    .A3(\w[13][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10163_));
 sky130_fd_sc_hd__mux4_2 _24296_ (.A0(_10159_),
    .A1(_10160_),
    .A2(_10161_),
    .A3(_10163_),
    .S0(net344),
    .S1(net335),
    .X(_10164_));
 sky130_fd_sc_hd__mux4_2 _24297_ (.A0(\w[51][19] ),
    .A1(\w[49][19] ),
    .A2(\w[55][19] ),
    .A3(\w[53][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_519 ();
 sky130_fd_sc_hd__mux4_2 _24299_ (.A0(\w[59][19] ),
    .A1(\w[57][19] ),
    .A2(\w[63][19] ),
    .A3(\w[61][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10167_));
 sky130_fd_sc_hd__mux4_2 _24300_ (.A0(\w[35][19] ),
    .A1(\w[33][19] ),
    .A2(\w[39][19] ),
    .A3(\w[37][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_518 ();
 sky130_fd_sc_hd__mux4_2 _24302_ (.A0(\w[43][19] ),
    .A1(\w[41][19] ),
    .A2(\w[47][19] ),
    .A3(\w[45][19] ),
    .S0(net370),
    .S1(net317),
    .X(_10170_));
 sky130_fd_sc_hd__mux4_2 _24303_ (.A0(_10165_),
    .A1(_10167_),
    .A2(_10168_),
    .A3(_10170_),
    .S0(net344),
    .S1(net335),
    .X(_10171_));
 sky130_fd_sc_hd__mux2i_1 _24304_ (.A0(_10164_),
    .A1(_10171_),
    .S(net297),
    .Y(_10172_));
 sky130_fd_sc_hd__nand2_2 _24305_ (.A(net357),
    .B(\w[1][19] ),
    .Y(_10173_));
 sky130_fd_sc_hd__o21ai_4 _24306_ (.A1(net292),
    .A2(_10172_),
    .B1(_10173_),
    .Y(_00042_));
 sky130_fd_sc_hd__mux4_2 _24307_ (.A0(\w[19][20] ),
    .A1(\w[17][20] ),
    .A2(\w[23][20] ),
    .A3(\w[21][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10174_));
 sky130_fd_sc_hd__mux4_2 _24308_ (.A0(\w[27][20] ),
    .A1(\w[25][20] ),
    .A2(\w[31][20] ),
    .A3(\w[29][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10175_));
 sky130_fd_sc_hd__mux4_2 _24309_ (.A0(\w[3][20] ),
    .A1(\w[1][20] ),
    .A2(\w[7][20] ),
    .A3(\w[5][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_517 ();
 sky130_fd_sc_hd__mux4_2 _24311_ (.A0(\w[11][20] ),
    .A1(\w[9][20] ),
    .A2(\w[15][20] ),
    .A3(\w[13][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10178_));
 sky130_fd_sc_hd__mux4_2 _24312_ (.A0(_10174_),
    .A1(_10175_),
    .A2(_10176_),
    .A3(_10178_),
    .S0(_09854_),
    .S1(net340),
    .X(_10179_));
 sky130_fd_sc_hd__mux4_2 _24313_ (.A0(\w[51][20] ),
    .A1(\w[49][20] ),
    .A2(\w[55][20] ),
    .A3(\w[53][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_516 ();
 sky130_fd_sc_hd__mux4_2 _24315_ (.A0(\w[59][20] ),
    .A1(\w[57][20] ),
    .A2(\w[63][20] ),
    .A3(\w[61][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10182_));
 sky130_fd_sc_hd__mux4_2 _24316_ (.A0(\w[35][20] ),
    .A1(\w[33][20] ),
    .A2(\w[39][20] ),
    .A3(\w[37][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10183_));
 sky130_fd_sc_hd__mux4_2 _24317_ (.A0(\w[43][20] ),
    .A1(\w[41][20] ),
    .A2(\w[47][20] ),
    .A3(\w[45][20] ),
    .S0(net372),
    .S1(_00657_),
    .X(_10184_));
 sky130_fd_sc_hd__mux4_2 _24318_ (.A0(_10180_),
    .A1(_10182_),
    .A2(_10183_),
    .A3(_10184_),
    .S0(_09854_),
    .S1(net340),
    .X(_10185_));
 sky130_fd_sc_hd__mux2i_1 _24319_ (.A0(_10179_),
    .A1(_10185_),
    .S(net300),
    .Y(_10186_));
 sky130_fd_sc_hd__nand2_1 _24320_ (.A(net540),
    .B(\w[1][20] ),
    .Y(_10187_));
 sky130_fd_sc_hd__o21ai_2 _24321_ (.A1(net292),
    .A2(_10186_),
    .B1(_10187_),
    .Y(_00044_));
 sky130_fd_sc_hd__mux4_2 _24322_ (.A0(\w[19][21] ),
    .A1(\w[17][21] ),
    .A2(\w[23][21] ),
    .A3(\w[21][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10188_));
 sky130_fd_sc_hd__mux4_2 _24323_ (.A0(\w[27][21] ),
    .A1(\w[25][21] ),
    .A2(\w[31][21] ),
    .A3(\w[29][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10189_));
 sky130_fd_sc_hd__mux4_2 _24324_ (.A0(\w[3][21] ),
    .A1(\w[1][21] ),
    .A2(\w[7][21] ),
    .A3(\w[5][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10190_));
 sky130_fd_sc_hd__mux4_2 _24325_ (.A0(\w[11][21] ),
    .A1(\w[9][21] ),
    .A2(\w[15][21] ),
    .A3(\w[13][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10191_));
 sky130_fd_sc_hd__mux4_2 _24326_ (.A0(_10188_),
    .A1(_10189_),
    .A2(_10190_),
    .A3(_10191_),
    .S0(net345),
    .S1(net335),
    .X(_10192_));
 sky130_fd_sc_hd__mux4_2 _24327_ (.A0(\w[51][21] ),
    .A1(\w[49][21] ),
    .A2(\w[55][21] ),
    .A3(\w[53][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10193_));
 sky130_fd_sc_hd__mux4_2 _24328_ (.A0(\w[59][21] ),
    .A1(\w[57][21] ),
    .A2(\w[63][21] ),
    .A3(\w[61][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10194_));
 sky130_fd_sc_hd__mux4_2 _24329_ (.A0(\w[35][21] ),
    .A1(\w[33][21] ),
    .A2(\w[39][21] ),
    .A3(\w[37][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10195_));
 sky130_fd_sc_hd__mux4_2 _24330_ (.A0(\w[43][21] ),
    .A1(\w[41][21] ),
    .A2(\w[47][21] ),
    .A3(\w[45][21] ),
    .S0(net371),
    .S1(net318),
    .X(_10196_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_515 ();
 sky130_fd_sc_hd__mux4_2 _24332_ (.A0(_10193_),
    .A1(_10194_),
    .A2(_10195_),
    .A3(_10196_),
    .S0(net344),
    .S1(net335),
    .X(_10198_));
 sky130_fd_sc_hd__mux2i_1 _24333_ (.A0(_10192_),
    .A1(_10198_),
    .S(net298),
    .Y(_10199_));
 sky130_fd_sc_hd__nand2_1 _24334_ (.A(net357),
    .B(\w[1][21] ),
    .Y(_10200_));
 sky130_fd_sc_hd__o21ai_0 _24335_ (.A1(net292),
    .A2(_10199_),
    .B1(_10200_),
    .Y(_00045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_514 ();
 sky130_fd_sc_hd__mux4_2 _24337_ (.A0(\w[19][22] ),
    .A1(\w[17][22] ),
    .A2(\w[23][22] ),
    .A3(\w[21][22] ),
    .S0(net371),
    .S1(net318),
    .X(_10202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_513 ();
 sky130_fd_sc_hd__mux4_2 _24339_ (.A0(\w[27][22] ),
    .A1(\w[25][22] ),
    .A2(\w[31][22] ),
    .A3(\w[29][22] ),
    .S0(net371),
    .S1(net318),
    .X(_10204_));
 sky130_fd_sc_hd__mux4_2 _24340_ (.A0(\w[3][22] ),
    .A1(\w[1][22] ),
    .A2(\w[7][22] ),
    .A3(\w[5][22] ),
    .S0(net371),
    .S1(net318),
    .X(_10205_));
 sky130_fd_sc_hd__mux4_2 _24341_ (.A0(\w[11][22] ),
    .A1(\w[9][22] ),
    .A2(\w[15][22] ),
    .A3(\w[13][22] ),
    .S0(net371),
    .S1(net318),
    .X(_10206_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_512 ();
 sky130_fd_sc_hd__mux4_2 _24343_ (.A0(_10202_),
    .A1(_10204_),
    .A2(_10205_),
    .A3(_10206_),
    .S0(net345),
    .S1(net335),
    .X(_10208_));
 sky130_fd_sc_hd__mux4_2 _24344_ (.A0(\w[51][22] ),
    .A1(\w[49][22] ),
    .A2(\w[55][22] ),
    .A3(\w[53][22] ),
    .S0(net370),
    .S1(net317),
    .X(_10209_));
 sky130_fd_sc_hd__mux4_2 _24345_ (.A0(\w[59][22] ),
    .A1(\w[57][22] ),
    .A2(\w[63][22] ),
    .A3(\w[61][22] ),
    .S0(net370),
    .S1(net317),
    .X(_10210_));
 sky130_fd_sc_hd__mux4_2 _24346_ (.A0(\w[35][22] ),
    .A1(\w[33][22] ),
    .A2(\w[39][22] ),
    .A3(\w[37][22] ),
    .S0(net370),
    .S1(net317),
    .X(_10211_));
 sky130_fd_sc_hd__mux4_2 _24347_ (.A0(\w[43][22] ),
    .A1(\w[41][22] ),
    .A2(\w[47][22] ),
    .A3(\w[45][22] ),
    .S0(net370),
    .S1(net317),
    .X(_10212_));
 sky130_fd_sc_hd__mux4_2 _24348_ (.A0(_10209_),
    .A1(_10210_),
    .A2(_10211_),
    .A3(_10212_),
    .S0(net343),
    .S1(net334),
    .X(_10213_));
 sky130_fd_sc_hd__mux2i_1 _24349_ (.A0(_10208_),
    .A1(_10213_),
    .S(net297),
    .Y(_10214_));
 sky130_fd_sc_hd__nand2_1 _24350_ (.A(net357),
    .B(\w[1][22] ),
    .Y(_10215_));
 sky130_fd_sc_hd__o21ai_0 _24351_ (.A1(net292),
    .A2(_10214_),
    .B1(_10215_),
    .Y(_00046_));
 sky130_fd_sc_hd__mux4_2 _24352_ (.A0(\w[19][23] ),
    .A1(\w[17][23] ),
    .A2(\w[23][23] ),
    .A3(\w[21][23] ),
    .S0(net365),
    .S1(net313),
    .X(_10216_));
 sky130_fd_sc_hd__mux4_2 _24353_ (.A0(\w[27][23] ),
    .A1(\w[25][23] ),
    .A2(\w[31][23] ),
    .A3(\w[29][23] ),
    .S0(net365),
    .S1(net313),
    .X(_10217_));
 sky130_fd_sc_hd__mux4_2 _24354_ (.A0(\w[3][23] ),
    .A1(\w[1][23] ),
    .A2(\w[7][23] ),
    .A3(\w[5][23] ),
    .S0(net365),
    .S1(net313),
    .X(_10218_));
 sky130_fd_sc_hd__mux4_2 _24355_ (.A0(\w[11][23] ),
    .A1(\w[9][23] ),
    .A2(\w[15][23] ),
    .A3(\w[13][23] ),
    .S0(net365),
    .S1(net313),
    .X(_10219_));
 sky130_fd_sc_hd__mux4_2 _24356_ (.A0(_10216_),
    .A1(_10217_),
    .A2(_10218_),
    .A3(_10219_),
    .S0(net342),
    .S1(net336),
    .X(_10220_));
 sky130_fd_sc_hd__mux4_2 _24357_ (.A0(\w[51][23] ),
    .A1(\w[49][23] ),
    .A2(\w[55][23] ),
    .A3(\w[53][23] ),
    .S0(net367),
    .S1(net313),
    .X(_10221_));
 sky130_fd_sc_hd__mux4_2 _24358_ (.A0(\w[59][23] ),
    .A1(\w[57][23] ),
    .A2(\w[63][23] ),
    .A3(\w[61][23] ),
    .S0(net367),
    .S1(net313),
    .X(_10222_));
 sky130_fd_sc_hd__mux4_2 _24359_ (.A0(\w[35][23] ),
    .A1(\w[33][23] ),
    .A2(\w[39][23] ),
    .A3(\w[37][23] ),
    .S0(net367),
    .S1(net313),
    .X(_10223_));
 sky130_fd_sc_hd__mux4_2 _24360_ (.A0(\w[43][23] ),
    .A1(\w[41][23] ),
    .A2(\w[47][23] ),
    .A3(\w[45][23] ),
    .S0(net367),
    .S1(net313),
    .X(_10224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_511 ();
 sky130_fd_sc_hd__mux4_2 _24362_ (.A0(_10221_),
    .A1(_10222_),
    .A2(_10223_),
    .A3(_10224_),
    .S0(net342),
    .S1(net338),
    .X(_10226_));
 sky130_fd_sc_hd__mux2i_1 _24363_ (.A0(_10220_),
    .A1(_10226_),
    .S(net299),
    .Y(_10227_));
 sky130_fd_sc_hd__nand2_2 _24364_ (.A(net357),
    .B(\w[1][23] ),
    .Y(_10228_));
 sky130_fd_sc_hd__o21ai_4 _24365_ (.A1(net291),
    .A2(_10227_),
    .B1(_10228_),
    .Y(_00047_));
 sky130_fd_sc_hd__mux4_2 _24366_ (.A0(\w[19][24] ),
    .A1(\w[17][24] ),
    .A2(\w[23][24] ),
    .A3(\w[21][24] ),
    .S0(net365),
    .S1(net316),
    .X(_10229_));
 sky130_fd_sc_hd__mux4_2 _24367_ (.A0(\w[27][24] ),
    .A1(\w[25][24] ),
    .A2(\w[31][24] ),
    .A3(\w[29][24] ),
    .S0(net365),
    .S1(net316),
    .X(_10230_));
 sky130_fd_sc_hd__mux4_2 _24368_ (.A0(\w[3][24] ),
    .A1(\w[1][24] ),
    .A2(\w[7][24] ),
    .A3(\w[5][24] ),
    .S0(net365),
    .S1(net316),
    .X(_10231_));
 sky130_fd_sc_hd__mux4_2 _24369_ (.A0(\w[11][24] ),
    .A1(\w[9][24] ),
    .A2(\w[15][24] ),
    .A3(\w[13][24] ),
    .S0(net365),
    .S1(net316),
    .X(_10232_));
 sky130_fd_sc_hd__mux4_2 _24370_ (.A0(_10229_),
    .A1(_10230_),
    .A2(_10231_),
    .A3(_10232_),
    .S0(net342),
    .S1(net336),
    .X(_10233_));
 sky130_fd_sc_hd__mux4_2 _24371_ (.A0(\w[51][24] ),
    .A1(\w[49][24] ),
    .A2(\w[55][24] ),
    .A3(\w[53][24] ),
    .S0(net365),
    .S1(net313),
    .X(_10234_));
 sky130_fd_sc_hd__mux4_2 _24372_ (.A0(\w[59][24] ),
    .A1(\w[57][24] ),
    .A2(\w[63][24] ),
    .A3(\w[61][24] ),
    .S0(net367),
    .S1(net313),
    .X(_10235_));
 sky130_fd_sc_hd__mux4_2 _24373_ (.A0(\w[35][24] ),
    .A1(\w[33][24] ),
    .A2(\w[39][24] ),
    .A3(\w[37][24] ),
    .S0(net367),
    .S1(net313),
    .X(_10236_));
 sky130_fd_sc_hd__mux4_2 _24374_ (.A0(\w[43][24] ),
    .A1(\w[41][24] ),
    .A2(\w[47][24] ),
    .A3(\w[45][24] ),
    .S0(net365),
    .S1(net313),
    .X(_10237_));
 sky130_fd_sc_hd__mux4_2 _24375_ (.A0(_10234_),
    .A1(_10235_),
    .A2(_10236_),
    .A3(_10237_),
    .S0(net342),
    .S1(net336),
    .X(_10238_));
 sky130_fd_sc_hd__mux2i_1 _24376_ (.A0(_10233_),
    .A1(_10238_),
    .S(net299),
    .Y(_10239_));
 sky130_fd_sc_hd__nand2_2 _24377_ (.A(net357),
    .B(\w[1][24] ),
    .Y(_10240_));
 sky130_fd_sc_hd__o21ai_4 _24378_ (.A1(net291),
    .A2(_10239_),
    .B1(_10240_),
    .Y(_00048_));
 sky130_fd_sc_hd__mux4_2 _24379_ (.A0(\w[19][25] ),
    .A1(\w[17][25] ),
    .A2(\w[23][25] ),
    .A3(\w[21][25] ),
    .S0(net370),
    .S1(net317),
    .X(_10241_));
 sky130_fd_sc_hd__mux4_2 _24380_ (.A0(\w[27][25] ),
    .A1(\w[25][25] ),
    .A2(\w[31][25] ),
    .A3(\w[29][25] ),
    .S0(net370),
    .S1(net317),
    .X(_10242_));
 sky130_fd_sc_hd__mux4_2 _24381_ (.A0(\w[3][25] ),
    .A1(\w[1][25] ),
    .A2(\w[7][25] ),
    .A3(\w[5][25] ),
    .S0(net370),
    .S1(net317),
    .X(_10243_));
 sky130_fd_sc_hd__mux4_2 _24382_ (.A0(\w[11][25] ),
    .A1(\w[9][25] ),
    .A2(\w[15][25] ),
    .A3(\w[13][25] ),
    .S0(net370),
    .S1(net317),
    .X(_10244_));
 sky130_fd_sc_hd__mux4_2 _24383_ (.A0(_10241_),
    .A1(_10242_),
    .A2(_10243_),
    .A3(_10244_),
    .S0(net344),
    .S1(net335),
    .X(_10245_));
 sky130_fd_sc_hd__mux4_2 _24384_ (.A0(\w[51][25] ),
    .A1(\w[49][25] ),
    .A2(\w[55][25] ),
    .A3(\w[53][25] ),
    .S0(net369),
    .S1(net315),
    .X(_10246_));
 sky130_fd_sc_hd__mux4_2 _24385_ (.A0(\w[59][25] ),
    .A1(\w[57][25] ),
    .A2(\w[63][25] ),
    .A3(\w[61][25] ),
    .S0(net369),
    .S1(net315),
    .X(_10247_));
 sky130_fd_sc_hd__mux4_2 _24386_ (.A0(\w[35][25] ),
    .A1(\w[33][25] ),
    .A2(\w[39][25] ),
    .A3(\w[37][25] ),
    .S0(net369),
    .S1(net315),
    .X(_10248_));
 sky130_fd_sc_hd__mux4_2 _24387_ (.A0(\w[43][25] ),
    .A1(\w[41][25] ),
    .A2(\w[47][25] ),
    .A3(\w[45][25] ),
    .S0(net369),
    .S1(net315),
    .X(_10249_));
 sky130_fd_sc_hd__mux4_2 _24388_ (.A0(_10246_),
    .A1(_10247_),
    .A2(_10248_),
    .A3(_10249_),
    .S0(net344),
    .S1(net335),
    .X(_10250_));
 sky130_fd_sc_hd__mux2i_1 _24389_ (.A0(_10245_),
    .A1(_10250_),
    .S(net297),
    .Y(_10251_));
 sky130_fd_sc_hd__nand2_2 _24390_ (.A(net357),
    .B(\w[1][25] ),
    .Y(_10252_));
 sky130_fd_sc_hd__o21ai_4 _24391_ (.A1(net292),
    .A2(_10251_),
    .B1(_10252_),
    .Y(_00049_));
 sky130_fd_sc_hd__mux4_2 _24392_ (.A0(\w[19][26] ),
    .A1(\w[17][26] ),
    .A2(\w[23][26] ),
    .A3(\w[21][26] ),
    .S0(net365),
    .S1(_00657_),
    .X(_10253_));
 sky130_fd_sc_hd__mux4_2 _24393_ (.A0(\w[27][26] ),
    .A1(\w[25][26] ),
    .A2(\w[31][26] ),
    .A3(\w[29][26] ),
    .S0(net365),
    .S1(net313),
    .X(_10254_));
 sky130_fd_sc_hd__mux4_2 _24394_ (.A0(\w[3][26] ),
    .A1(\w[1][26] ),
    .A2(\w[7][26] ),
    .A3(\w[5][26] ),
    .S0(net365),
    .S1(_00657_),
    .X(_10255_));
 sky130_fd_sc_hd__mux4_2 _24395_ (.A0(\w[11][26] ),
    .A1(\w[9][26] ),
    .A2(\w[15][26] ),
    .A3(\w[13][26] ),
    .S0(net365),
    .S1(_00657_),
    .X(_10256_));
 sky130_fd_sc_hd__mux4_2 _24396_ (.A0(_10253_),
    .A1(_10254_),
    .A2(_10255_),
    .A3(_10256_),
    .S0(net342),
    .S1(net336),
    .X(_10257_));
 sky130_fd_sc_hd__mux4_2 _24397_ (.A0(\w[51][26] ),
    .A1(\w[49][26] ),
    .A2(\w[55][26] ),
    .A3(\w[53][26] ),
    .S0(net366),
    .S1(net313),
    .X(_10258_));
 sky130_fd_sc_hd__mux4_2 _24398_ (.A0(\w[59][26] ),
    .A1(\w[57][26] ),
    .A2(\w[63][26] ),
    .A3(\w[61][26] ),
    .S0(net366),
    .S1(net313),
    .X(_10259_));
 sky130_fd_sc_hd__mux4_2 _24399_ (.A0(\w[35][26] ),
    .A1(\w[33][26] ),
    .A2(\w[39][26] ),
    .A3(\w[37][26] ),
    .S0(net366),
    .S1(net313),
    .X(_10260_));
 sky130_fd_sc_hd__mux4_2 _24400_ (.A0(\w[43][26] ),
    .A1(\w[41][26] ),
    .A2(\w[47][26] ),
    .A3(\w[45][26] ),
    .S0(net366),
    .S1(net313),
    .X(_10261_));
 sky130_fd_sc_hd__mux4_2 _24401_ (.A0(_10258_),
    .A1(_10259_),
    .A2(_10260_),
    .A3(_10261_),
    .S0(net341),
    .S1(net338),
    .X(_10262_));
 sky130_fd_sc_hd__mux2i_1 _24402_ (.A0(_10257_),
    .A1(_10262_),
    .S(net299),
    .Y(_10263_));
 sky130_fd_sc_hd__nand2_2 _24403_ (.A(net357),
    .B(\w[1][26] ),
    .Y(_10264_));
 sky130_fd_sc_hd__o21ai_4 _24404_ (.A1(net291),
    .A2(_10263_),
    .B1(_10264_),
    .Y(_00050_));
 sky130_fd_sc_hd__mux4_2 _24405_ (.A0(\w[19][27] ),
    .A1(\w[17][27] ),
    .A2(\w[23][27] ),
    .A3(\w[21][27] ),
    .S0(net368),
    .S1(net314),
    .X(_10265_));
 sky130_fd_sc_hd__mux4_2 _24406_ (.A0(\w[27][27] ),
    .A1(\w[25][27] ),
    .A2(\w[31][27] ),
    .A3(\w[29][27] ),
    .S0(net368),
    .S1(net314),
    .X(_10266_));
 sky130_fd_sc_hd__mux4_2 _24407_ (.A0(\w[3][27] ),
    .A1(\w[1][27] ),
    .A2(\w[7][27] ),
    .A3(\w[5][27] ),
    .S0(net368),
    .S1(net314),
    .X(_10267_));
 sky130_fd_sc_hd__mux4_2 _24408_ (.A0(\w[11][27] ),
    .A1(\w[9][27] ),
    .A2(\w[15][27] ),
    .A3(\w[13][27] ),
    .S0(net368),
    .S1(net314),
    .X(_10268_));
 sky130_fd_sc_hd__mux4_2 _24409_ (.A0(_10265_),
    .A1(_10266_),
    .A2(_10267_),
    .A3(_10268_),
    .S0(net343),
    .S1(net334),
    .X(_10269_));
 sky130_fd_sc_hd__mux4_2 _24410_ (.A0(\w[51][27] ),
    .A1(\w[49][27] ),
    .A2(\w[55][27] ),
    .A3(\w[53][27] ),
    .S0(net367),
    .S1(net313),
    .X(_10270_));
 sky130_fd_sc_hd__mux4_2 _24411_ (.A0(\w[59][27] ),
    .A1(\w[57][27] ),
    .A2(\w[63][27] ),
    .A3(\w[61][27] ),
    .S0(net367),
    .S1(net313),
    .X(_10271_));
 sky130_fd_sc_hd__mux4_2 _24412_ (.A0(\w[35][27] ),
    .A1(\w[33][27] ),
    .A2(\w[39][27] ),
    .A3(\w[37][27] ),
    .S0(net367),
    .S1(net313),
    .X(_10272_));
 sky130_fd_sc_hd__mux4_2 _24413_ (.A0(\w[43][27] ),
    .A1(\w[41][27] ),
    .A2(\w[47][27] ),
    .A3(\w[45][27] ),
    .S0(net367),
    .S1(net313),
    .X(_10273_));
 sky130_fd_sc_hd__mux4_2 _24414_ (.A0(_10270_),
    .A1(_10271_),
    .A2(_10272_),
    .A3(_10273_),
    .S0(net342),
    .S1(net336),
    .X(_10274_));
 sky130_fd_sc_hd__mux2i_1 _24415_ (.A0(_10269_),
    .A1(_10274_),
    .S(net297),
    .Y(_10275_));
 sky130_fd_sc_hd__nand2_1 _24416_ (.A(net357),
    .B(\w[1][27] ),
    .Y(_10276_));
 sky130_fd_sc_hd__o21ai_4 _24417_ (.A1(net292),
    .A2(_10275_),
    .B1(_10276_),
    .Y(_00051_));
 sky130_fd_sc_hd__mux4_2 _24418_ (.A0(\w[19][28] ),
    .A1(\w[17][28] ),
    .A2(\w[23][28] ),
    .A3(\w[21][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10277_));
 sky130_fd_sc_hd__mux4_2 _24419_ (.A0(\w[27][28] ),
    .A1(\w[25][28] ),
    .A2(\w[31][28] ),
    .A3(\w[29][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10278_));
 sky130_fd_sc_hd__mux4_2 _24420_ (.A0(\w[3][28] ),
    .A1(\w[1][28] ),
    .A2(\w[7][28] ),
    .A3(\w[5][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10279_));
 sky130_fd_sc_hd__mux4_2 _24421_ (.A0(\w[11][28] ),
    .A1(\w[9][28] ),
    .A2(\w[15][28] ),
    .A3(\w[13][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10280_));
 sky130_fd_sc_hd__mux4_2 _24422_ (.A0(_10277_),
    .A1(_10278_),
    .A2(_10279_),
    .A3(_10280_),
    .S0(net342),
    .S1(net336),
    .X(_10281_));
 sky130_fd_sc_hd__mux4_2 _24423_ (.A0(\w[51][28] ),
    .A1(\w[49][28] ),
    .A2(\w[55][28] ),
    .A3(\w[53][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10282_));
 sky130_fd_sc_hd__mux4_2 _24424_ (.A0(\w[59][28] ),
    .A1(\w[57][28] ),
    .A2(\w[63][28] ),
    .A3(\w[61][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10283_));
 sky130_fd_sc_hd__mux4_2 _24425_ (.A0(\w[35][28] ),
    .A1(\w[33][28] ),
    .A2(\w[39][28] ),
    .A3(\w[37][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10284_));
 sky130_fd_sc_hd__mux4_2 _24426_ (.A0(\w[43][28] ),
    .A1(\w[41][28] ),
    .A2(\w[47][28] ),
    .A3(\w[45][28] ),
    .S0(net365),
    .S1(net313),
    .X(_10285_));
 sky130_fd_sc_hd__mux4_2 _24427_ (.A0(_10282_),
    .A1(_10283_),
    .A2(_10284_),
    .A3(_10285_),
    .S0(net342),
    .S1(net336),
    .X(_10286_));
 sky130_fd_sc_hd__mux2i_1 _24428_ (.A0(_10281_),
    .A1(_10286_),
    .S(net299),
    .Y(_10287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_510 ();
 sky130_fd_sc_hd__nand2_2 _24430_ (.A(net357),
    .B(\w[1][28] ),
    .Y(_10289_));
 sky130_fd_sc_hd__o21ai_4 _24431_ (.A1(net291),
    .A2(_10287_),
    .B1(_10289_),
    .Y(_00052_));
 sky130_fd_sc_hd__mux4_2 _24432_ (.A0(\w[19][29] ),
    .A1(\w[17][29] ),
    .A2(\w[23][29] ),
    .A3(\w[21][29] ),
    .S0(net365),
    .S1(net313),
    .X(_10290_));
 sky130_fd_sc_hd__mux4_2 _24433_ (.A0(\w[27][29] ),
    .A1(\w[25][29] ),
    .A2(\w[31][29] ),
    .A3(\w[29][29] ),
    .S0(net365),
    .S1(net313),
    .X(_10291_));
 sky130_fd_sc_hd__mux4_2 _24434_ (.A0(\w[3][29] ),
    .A1(\w[1][29] ),
    .A2(\w[7][29] ),
    .A3(\w[5][29] ),
    .S0(net365),
    .S1(net313),
    .X(_10292_));
 sky130_fd_sc_hd__mux4_2 _24435_ (.A0(\w[11][29] ),
    .A1(\w[9][29] ),
    .A2(\w[15][29] ),
    .A3(\w[13][29] ),
    .S0(net365),
    .S1(net313),
    .X(_10293_));
 sky130_fd_sc_hd__mux4_2 _24436_ (.A0(_10290_),
    .A1(_10291_),
    .A2(_10292_),
    .A3(_10293_),
    .S0(net342),
    .S1(net336),
    .X(_10294_));
 sky130_fd_sc_hd__mux4_2 _24437_ (.A0(\w[51][29] ),
    .A1(\w[49][29] ),
    .A2(\w[55][29] ),
    .A3(\w[53][29] ),
    .S0(net365),
    .S1(net313),
    .X(_10295_));
 sky130_fd_sc_hd__mux4_2 _24438_ (.A0(\w[59][29] ),
    .A1(\w[57][29] ),
    .A2(\w[63][29] ),
    .A3(\w[61][29] ),
    .S0(net365),
    .S1(net313),
    .X(_10296_));
 sky130_fd_sc_hd__mux4_2 _24439_ (.A0(\w[35][29] ),
    .A1(\w[33][29] ),
    .A2(\w[39][29] ),
    .A3(\w[37][29] ),
    .S0(net366),
    .S1(net313),
    .X(_10297_));
 sky130_fd_sc_hd__mux4_2 _24440_ (.A0(\w[43][29] ),
    .A1(\w[41][29] ),
    .A2(\w[47][29] ),
    .A3(\w[45][29] ),
    .S0(net365),
    .S1(net313),
    .X(_10298_));
 sky130_fd_sc_hd__mux4_2 _24441_ (.A0(_10295_),
    .A1(_10296_),
    .A2(_10297_),
    .A3(_10298_),
    .S0(net341),
    .S1(net338),
    .X(_10299_));
 sky130_fd_sc_hd__mux2i_1 _24442_ (.A0(_10294_),
    .A1(_10299_),
    .S(net299),
    .Y(_10300_));
 sky130_fd_sc_hd__nand2_2 _24443_ (.A(net357),
    .B(\w[1][29] ),
    .Y(_10301_));
 sky130_fd_sc_hd__o21ai_4 _24444_ (.A1(net291),
    .A2(_10300_),
    .B1(_10301_),
    .Y(_00053_));
 sky130_fd_sc_hd__mux4_2 _24445_ (.A0(\w[19][30] ),
    .A1(\w[17][30] ),
    .A2(\w[23][30] ),
    .A3(\w[21][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10302_));
 sky130_fd_sc_hd__mux4_2 _24446_ (.A0(\w[27][30] ),
    .A1(\w[25][30] ),
    .A2(\w[31][30] ),
    .A3(\w[29][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10303_));
 sky130_fd_sc_hd__mux4_2 _24447_ (.A0(\w[3][30] ),
    .A1(\w[1][30] ),
    .A2(\w[7][30] ),
    .A3(\w[5][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10304_));
 sky130_fd_sc_hd__mux4_2 _24448_ (.A0(\w[11][30] ),
    .A1(\w[9][30] ),
    .A2(\w[15][30] ),
    .A3(\w[13][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10305_));
 sky130_fd_sc_hd__mux4_2 _24449_ (.A0(_10302_),
    .A1(_10303_),
    .A2(_10304_),
    .A3(_10305_),
    .S0(net341),
    .S1(net340),
    .X(_10306_));
 sky130_fd_sc_hd__mux4_2 _24450_ (.A0(\w[51][30] ),
    .A1(\w[49][30] ),
    .A2(\w[55][30] ),
    .A3(\w[53][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10307_));
 sky130_fd_sc_hd__mux4_2 _24451_ (.A0(\w[59][30] ),
    .A1(\w[57][30] ),
    .A2(\w[63][30] ),
    .A3(\w[61][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10308_));
 sky130_fd_sc_hd__mux4_2 _24452_ (.A0(\w[35][30] ),
    .A1(\w[33][30] ),
    .A2(\w[39][30] ),
    .A3(\w[37][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10309_));
 sky130_fd_sc_hd__mux4_2 _24453_ (.A0(\w[43][30] ),
    .A1(\w[41][30] ),
    .A2(\w[47][30] ),
    .A3(\w[45][30] ),
    .S0(net366),
    .S1(_00657_),
    .X(_10310_));
 sky130_fd_sc_hd__mux4_2 _24454_ (.A0(_10307_),
    .A1(_10308_),
    .A2(_10309_),
    .A3(_10310_),
    .S0(net341),
    .S1(net340),
    .X(_10311_));
 sky130_fd_sc_hd__mux2i_1 _24455_ (.A0(_10306_),
    .A1(_10311_),
    .S(net299),
    .Y(_10312_));
 sky130_fd_sc_hd__nand2_2 _24456_ (.A(net357),
    .B(\w[1][30] ),
    .Y(_10313_));
 sky130_fd_sc_hd__o21ai_4 _24457_ (.A1(net291),
    .A2(_10312_),
    .B1(_10313_),
    .Y(_00055_));
 sky130_fd_sc_hd__mux4_2 _24458_ (.A0(\w[19][31] ),
    .A1(\w[17][31] ),
    .A2(\w[23][31] ),
    .A3(\w[21][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10314_));
 sky130_fd_sc_hd__mux4_2 _24459_ (.A0(\w[27][31] ),
    .A1(\w[25][31] ),
    .A2(\w[31][31] ),
    .A3(\w[29][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10315_));
 sky130_fd_sc_hd__mux4_2 _24460_ (.A0(\w[3][31] ),
    .A1(\w[1][31] ),
    .A2(\w[7][31] ),
    .A3(\w[5][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10316_));
 sky130_fd_sc_hd__mux4_2 _24461_ (.A0(\w[11][31] ),
    .A1(\w[9][31] ),
    .A2(\w[15][31] ),
    .A3(\w[13][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10317_));
 sky130_fd_sc_hd__mux4_2 _24462_ (.A0(_10314_),
    .A1(_10315_),
    .A2(_10316_),
    .A3(_10317_),
    .S0(net343),
    .S1(net334),
    .X(_10318_));
 sky130_fd_sc_hd__mux4_2 _24463_ (.A0(\w[51][31] ),
    .A1(\w[49][31] ),
    .A2(\w[55][31] ),
    .A3(\w[53][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10319_));
 sky130_fd_sc_hd__mux4_2 _24464_ (.A0(\w[59][31] ),
    .A1(\w[57][31] ),
    .A2(\w[63][31] ),
    .A3(\w[61][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10320_));
 sky130_fd_sc_hd__mux4_2 _24465_ (.A0(\w[35][31] ),
    .A1(\w[33][31] ),
    .A2(\w[39][31] ),
    .A3(\w[37][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10321_));
 sky130_fd_sc_hd__mux4_2 _24466_ (.A0(\w[43][31] ),
    .A1(\w[41][31] ),
    .A2(\w[47][31] ),
    .A3(\w[45][31] ),
    .S0(net369),
    .S1(net315),
    .X(_10322_));
 sky130_fd_sc_hd__mux4_2 _24467_ (.A0(_10319_),
    .A1(_10320_),
    .A2(_10321_),
    .A3(_10322_),
    .S0(net343),
    .S1(net337),
    .X(_10323_));
 sky130_fd_sc_hd__mux2i_1 _24468_ (.A0(_10318_),
    .A1(_10323_),
    .S(net297),
    .Y(_10324_));
 sky130_fd_sc_hd__nand2_2 _24469_ (.A(net357),
    .B(\w[1][31] ),
    .Y(_10325_));
 sky130_fd_sc_hd__o21ai_4 _24470_ (.A1(net292),
    .A2(_10324_),
    .B1(_10325_),
    .Y(_00056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_503 ();
 sky130_fd_sc_hd__mux4_2 _24478_ (.A0(\w[18][0] ),
    .A1(\w[16][0] ),
    .A2(\w[22][0] ),
    .A3(\w[20][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_499 ();
 sky130_fd_sc_hd__mux4_2 _24483_ (.A0(\w[26][0] ),
    .A1(\w[24][0] ),
    .A2(\w[30][0] ),
    .A3(\w[28][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_497 ();
 sky130_fd_sc_hd__mux4_2 _24486_ (.A0(\w[2][0] ),
    .A1(\w[0][0] ),
    .A2(\w[6][0] ),
    .A3(\w[4][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10341_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_493 ();
 sky130_fd_sc_hd__mux4_2 _24491_ (.A0(\w[10][0] ),
    .A1(\w[8][0] ),
    .A2(\w[14][0] ),
    .A3(\w[12][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10346_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_492 ();
 sky130_fd_sc_hd__xor2_4 _24493_ (.A(\count_hash1[3] ),
    .B(_12920_),
    .X(_10348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_490 ();
 sky130_fd_sc_hd__nand3_4 _24496_ (.A(\count_hash1[3] ),
    .B(\count_hash1[2] ),
    .C(\count_hash1[1] ),
    .Y(_10351_));
 sky130_fd_sc_hd__xor2_4 _24497_ (.A(\count_hash1[4] ),
    .B(_10351_),
    .X(_10352_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_488 ();
 sky130_fd_sc_hd__mux4_2 _24500_ (.A0(_10333_),
    .A1(_10338_),
    .A2(_10341_),
    .A3(_10346_),
    .S0(net333),
    .S1(net322),
    .X(_10355_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_486 ();
 sky130_fd_sc_hd__mux4_2 _24503_ (.A0(\w[50][0] ),
    .A1(\w[48][0] ),
    .A2(\w[54][0] ),
    .A3(\w[52][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10358_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_484 ();
 sky130_fd_sc_hd__mux4_2 _24506_ (.A0(\w[58][0] ),
    .A1(\w[56][0] ),
    .A2(\w[62][0] ),
    .A3(\w[60][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10361_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_482 ();
 sky130_fd_sc_hd__mux4_2 _24509_ (.A0(\w[34][0] ),
    .A1(\w[32][0] ),
    .A2(\w[38][0] ),
    .A3(\w[36][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_480 ();
 sky130_fd_sc_hd__mux4_2 _24512_ (.A0(\w[42][0] ),
    .A1(\w[40][0] ),
    .A2(\w[46][0] ),
    .A3(\w[44][0] ),
    .S0(net377),
    .S1(net312),
    .X(_10367_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_477 ();
 sky130_fd_sc_hd__mux4_2 _24516_ (.A0(_10358_),
    .A1(_10361_),
    .A2(_10364_),
    .A3(_10367_),
    .S0(net331),
    .S1(net322),
    .X(_10371_));
 sky130_fd_sc_hd__nand3_4 _24517_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(_12920_),
    .Y(_10372_));
 sky130_fd_sc_hd__xnor2_4 _24518_ (.A(\count_hash1[5] ),
    .B(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_474 ();
 sky130_fd_sc_hd__mux2i_1 _24522_ (.A0(_10355_),
    .A1(_10371_),
    .S(net296),
    .Y(_10377_));
 sky130_fd_sc_hd__nand2_1 _24523_ (.A(net356),
    .B(\w[0][0] ),
    .Y(_10378_));
 sky130_fd_sc_hd__o21ai_0 _24524_ (.A1(_09875_),
    .A2(_10377_),
    .B1(_10378_),
    .Y(_00000_));
 sky130_fd_sc_hd__mux4_2 _24525_ (.A0(\w[18][1] ),
    .A1(\w[16][1] ),
    .A2(\w[22][1] ),
    .A3(\w[20][1] ),
    .S0(net376),
    .S1(net311),
    .X(_10379_));
 sky130_fd_sc_hd__mux4_2 _24526_ (.A0(\w[26][1] ),
    .A1(\w[24][1] ),
    .A2(\w[30][1] ),
    .A3(\w[28][1] ),
    .S0(net376),
    .S1(net311),
    .X(_10380_));
 sky130_fd_sc_hd__mux4_2 _24527_ (.A0(\w[2][1] ),
    .A1(\w[0][1] ),
    .A2(\w[6][1] ),
    .A3(\w[4][1] ),
    .S0(net376),
    .S1(net311),
    .X(_10381_));
 sky130_fd_sc_hd__mux4_2 _24528_ (.A0(\w[10][1] ),
    .A1(\w[8][1] ),
    .A2(\w[14][1] ),
    .A3(\w[12][1] ),
    .S0(net376),
    .S1(net311),
    .X(_10382_));
 sky130_fd_sc_hd__mux4_2 _24529_ (.A0(_10379_),
    .A1(_10380_),
    .A2(_10381_),
    .A3(_10382_),
    .S0(net329),
    .S1(net323),
    .X(_10383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_473 ();
 sky130_fd_sc_hd__mux4_2 _24531_ (.A0(\w[50][1] ),
    .A1(\w[48][1] ),
    .A2(\w[54][1] ),
    .A3(\w[52][1] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10385_));
 sky130_fd_sc_hd__mux4_2 _24532_ (.A0(\w[58][1] ),
    .A1(\w[56][1] ),
    .A2(\w[62][1] ),
    .A3(\w[60][1] ),
    .S0(net541),
    .S1(net312),
    .X(_10386_));
 sky130_fd_sc_hd__mux4_2 _24533_ (.A0(\w[34][1] ),
    .A1(\w[32][1] ),
    .A2(\w[38][1] ),
    .A3(\w[36][1] ),
    .S0(net376),
    .S1(net311),
    .X(_10387_));
 sky130_fd_sc_hd__mux4_2 _24534_ (.A0(\w[42][1] ),
    .A1(\w[40][1] ),
    .A2(\w[46][1] ),
    .A3(\w[44][1] ),
    .S0(net376),
    .S1(net311),
    .X(_10388_));
 sky130_fd_sc_hd__mux4_2 _24535_ (.A0(_10385_),
    .A1(_10386_),
    .A2(_10387_),
    .A3(_10388_),
    .S0(net330),
    .S1(net323),
    .X(_10389_));
 sky130_fd_sc_hd__mux2i_1 _24536_ (.A0(_10383_),
    .A1(_10389_),
    .S(net295),
    .Y(_10390_));
 sky130_fd_sc_hd__nand2_2 _24537_ (.A(net356),
    .B(\w[0][1] ),
    .Y(_10391_));
 sky130_fd_sc_hd__o21ai_0 _24538_ (.A1(_09875_),
    .A2(_10390_),
    .B1(_10391_),
    .Y(_00011_));
 sky130_fd_sc_hd__mux4_2 _24539_ (.A0(\w[18][2] ),
    .A1(\w[16][2] ),
    .A2(\w[22][2] ),
    .A3(\w[20][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10392_));
 sky130_fd_sc_hd__mux4_2 _24540_ (.A0(\w[26][2] ),
    .A1(\w[24][2] ),
    .A2(\w[30][2] ),
    .A3(\w[28][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10393_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_472 ();
 sky130_fd_sc_hd__mux4_2 _24542_ (.A0(\w[2][2] ),
    .A1(\w[0][2] ),
    .A2(\w[6][2] ),
    .A3(\w[4][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10395_));
 sky130_fd_sc_hd__mux4_2 _24543_ (.A0(\w[10][2] ),
    .A1(\w[8][2] ),
    .A2(\w[14][2] ),
    .A3(\w[12][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10396_));
 sky130_fd_sc_hd__mux4_2 _24544_ (.A0(_10392_),
    .A1(_10393_),
    .A2(_10395_),
    .A3(_10396_),
    .S0(net327),
    .S1(net320),
    .X(_10397_));
 sky130_fd_sc_hd__mux4_2 _24545_ (.A0(\w[50][2] ),
    .A1(\w[48][2] ),
    .A2(\w[54][2] ),
    .A3(\w[52][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10398_));
 sky130_fd_sc_hd__mux4_2 _24546_ (.A0(\w[58][2] ),
    .A1(\w[56][2] ),
    .A2(\w[62][2] ),
    .A3(\w[60][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10399_));
 sky130_fd_sc_hd__mux4_2 _24547_ (.A0(\w[34][2] ),
    .A1(\w[32][2] ),
    .A2(\w[38][2] ),
    .A3(\w[36][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10400_));
 sky130_fd_sc_hd__mux4_2 _24548_ (.A0(\w[42][2] ),
    .A1(\w[40][2] ),
    .A2(\w[46][2] ),
    .A3(\w[44][2] ),
    .S0(net374),
    .S1(net308),
    .X(_10401_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_471 ();
 sky130_fd_sc_hd__mux4_2 _24550_ (.A0(_10398_),
    .A1(_10399_),
    .A2(_10400_),
    .A3(_10401_),
    .S0(net327),
    .S1(net320),
    .X(_10403_));
 sky130_fd_sc_hd__mux2i_1 _24551_ (.A0(_10397_),
    .A1(_10403_),
    .S(net293),
    .Y(_10404_));
 sky130_fd_sc_hd__nand2_2 _24552_ (.A(net356),
    .B(\w[0][2] ),
    .Y(_10405_));
 sky130_fd_sc_hd__o21ai_4 _24553_ (.A1(net290),
    .A2(_10404_),
    .B1(_10405_),
    .Y(_00022_));
 sky130_fd_sc_hd__mux4_2 _24554_ (.A0(\w[18][3] ),
    .A1(\w[16][3] ),
    .A2(\w[22][3] ),
    .A3(\w[20][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10406_));
 sky130_fd_sc_hd__mux4_2 _24555_ (.A0(\w[26][3] ),
    .A1(\w[24][3] ),
    .A2(\w[30][3] ),
    .A3(\w[28][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10407_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_470 ();
 sky130_fd_sc_hd__mux4_2 _24557_ (.A0(\w[2][3] ),
    .A1(\w[0][3] ),
    .A2(\w[6][3] ),
    .A3(\w[4][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10409_));
 sky130_fd_sc_hd__mux4_2 _24558_ (.A0(\w[10][3] ),
    .A1(\w[8][3] ),
    .A2(\w[14][3] ),
    .A3(\w[12][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10410_));
 sky130_fd_sc_hd__mux4_2 _24559_ (.A0(_10406_),
    .A1(_10407_),
    .A2(_10409_),
    .A3(_10410_),
    .S0(net326),
    .S1(net319),
    .X(_10411_));
 sky130_fd_sc_hd__mux4_2 _24560_ (.A0(\w[50][3] ),
    .A1(\w[48][3] ),
    .A2(\w[54][3] ),
    .A3(\w[52][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10412_));
 sky130_fd_sc_hd__mux4_2 _24561_ (.A0(\w[58][3] ),
    .A1(\w[56][3] ),
    .A2(\w[62][3] ),
    .A3(\w[60][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10413_));
 sky130_fd_sc_hd__mux4_2 _24562_ (.A0(\w[34][3] ),
    .A1(\w[32][3] ),
    .A2(\w[38][3] ),
    .A3(\w[36][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10414_));
 sky130_fd_sc_hd__mux4_2 _24563_ (.A0(\w[42][3] ),
    .A1(\w[40][3] ),
    .A2(\w[46][3] ),
    .A3(\w[44][3] ),
    .S0(net373),
    .S1(net309),
    .X(_10415_));
 sky130_fd_sc_hd__mux4_2 _24564_ (.A0(_10412_),
    .A1(_10413_),
    .A2(_10414_),
    .A3(_10415_),
    .S0(net326),
    .S1(net319),
    .X(_10416_));
 sky130_fd_sc_hd__mux2i_1 _24565_ (.A0(_10411_),
    .A1(_10416_),
    .S(net294),
    .Y(_10417_));
 sky130_fd_sc_hd__nand2_2 _24566_ (.A(reset_hash),
    .B(\w[0][3] ),
    .Y(_10418_));
 sky130_fd_sc_hd__o21ai_4 _24567_ (.A1(net291),
    .A2(_10417_),
    .B1(_10418_),
    .Y(_00025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_469 ();
 sky130_fd_sc_hd__mux4_2 _24569_ (.A0(\w[18][4] ),
    .A1(\w[16][4] ),
    .A2(\w[22][4] ),
    .A3(\w[20][4] ),
    .S0(net374),
    .S1(net308),
    .X(_10420_));
 sky130_fd_sc_hd__mux4_2 _24570_ (.A0(\w[26][4] ),
    .A1(\w[24][4] ),
    .A2(\w[30][4] ),
    .A3(\w[28][4] ),
    .S0(net374),
    .S1(net308),
    .X(_10421_));
 sky130_fd_sc_hd__mux4_2 _24571_ (.A0(\w[2][4] ),
    .A1(\w[0][4] ),
    .A2(\w[6][4] ),
    .A3(\w[4][4] ),
    .S0(net374),
    .S1(net308),
    .X(_10422_));
 sky130_fd_sc_hd__mux4_2 _24572_ (.A0(\w[10][4] ),
    .A1(\w[8][4] ),
    .A2(\w[14][4] ),
    .A3(\w[12][4] ),
    .S0(net374),
    .S1(net308),
    .X(_10423_));
 sky130_fd_sc_hd__mux4_2 _24573_ (.A0(_10420_),
    .A1(_10421_),
    .A2(_10422_),
    .A3(_10423_),
    .S0(net326),
    .S1(net319),
    .X(_10424_));
 sky130_fd_sc_hd__mux4_2 _24574_ (.A0(\w[50][4] ),
    .A1(\w[48][4] ),
    .A2(\w[54][4] ),
    .A3(\w[52][4] ),
    .S0(net373),
    .S1(net309),
    .X(_10425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_468 ();
 sky130_fd_sc_hd__mux4_2 _24576_ (.A0(\w[58][4] ),
    .A1(\w[56][4] ),
    .A2(\w[62][4] ),
    .A3(\w[60][4] ),
    .S0(net373),
    .S1(net309),
    .X(_10427_));
 sky130_fd_sc_hd__mux4_2 _24577_ (.A0(\w[34][4] ),
    .A1(\w[32][4] ),
    .A2(\w[38][4] ),
    .A3(\w[36][4] ),
    .S0(net374),
    .S1(net308),
    .X(_10428_));
 sky130_fd_sc_hd__mux4_2 _24578_ (.A0(\w[42][4] ),
    .A1(\w[40][4] ),
    .A2(\w[46][4] ),
    .A3(\w[44][4] ),
    .S0(net373),
    .S1(net309),
    .X(_10429_));
 sky130_fd_sc_hd__mux4_2 _24579_ (.A0(_10425_),
    .A1(_10427_),
    .A2(_10428_),
    .A3(_10429_),
    .S0(net326),
    .S1(net319),
    .X(_10430_));
 sky130_fd_sc_hd__mux2i_1 _24580_ (.A0(_10424_),
    .A1(_10430_),
    .S(net294),
    .Y(_10431_));
 sky130_fd_sc_hd__nand2_2 _24581_ (.A(net356),
    .B(\w[0][4] ),
    .Y(_10432_));
 sky130_fd_sc_hd__o21ai_4 _24582_ (.A1(net290),
    .A2(_10431_),
    .B1(_10432_),
    .Y(_00026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_467 ();
 sky130_fd_sc_hd__mux4_2 _24584_ (.A0(\w[18][5] ),
    .A1(\w[16][5] ),
    .A2(\w[22][5] ),
    .A3(\w[20][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10434_));
 sky130_fd_sc_hd__mux4_2 _24585_ (.A0(\w[26][5] ),
    .A1(\w[24][5] ),
    .A2(\w[30][5] ),
    .A3(\w[28][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10435_));
 sky130_fd_sc_hd__mux4_2 _24586_ (.A0(\w[2][5] ),
    .A1(\w[0][5] ),
    .A2(\w[6][5] ),
    .A3(\w[4][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10436_));
 sky130_fd_sc_hd__mux4_2 _24587_ (.A0(\w[10][5] ),
    .A1(\w[8][5] ),
    .A2(\w[14][5] ),
    .A3(\w[12][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_466 ();
 sky130_fd_sc_hd__mux4_2 _24589_ (.A0(_10434_),
    .A1(_10435_),
    .A2(_10436_),
    .A3(_10437_),
    .S0(net326),
    .S1(net319),
    .X(_10439_));
 sky130_fd_sc_hd__mux4_2 _24590_ (.A0(\w[50][5] ),
    .A1(\w[48][5] ),
    .A2(\w[54][5] ),
    .A3(\w[52][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10440_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_465 ();
 sky130_fd_sc_hd__mux4_2 _24592_ (.A0(\w[58][5] ),
    .A1(\w[56][5] ),
    .A2(\w[62][5] ),
    .A3(\w[60][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10442_));
 sky130_fd_sc_hd__mux4_2 _24593_ (.A0(\w[34][5] ),
    .A1(\w[32][5] ),
    .A2(\w[38][5] ),
    .A3(\w[36][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10443_));
 sky130_fd_sc_hd__mux4_2 _24594_ (.A0(\w[42][5] ),
    .A1(\w[40][5] ),
    .A2(\w[46][5] ),
    .A3(\w[44][5] ),
    .S0(net373),
    .S1(net309),
    .X(_10444_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_464 ();
 sky130_fd_sc_hd__mux4_2 _24596_ (.A0(_10440_),
    .A1(_10442_),
    .A2(_10443_),
    .A3(_10444_),
    .S0(net326),
    .S1(net319),
    .X(_10446_));
 sky130_fd_sc_hd__mux2i_1 _24597_ (.A0(_10439_),
    .A1(_10446_),
    .S(net294),
    .Y(_10447_));
 sky130_fd_sc_hd__nand2_2 _24598_ (.A(net356),
    .B(\w[0][5] ),
    .Y(_10448_));
 sky130_fd_sc_hd__o21ai_4 _24599_ (.A1(net290),
    .A2(_10447_),
    .B1(_10448_),
    .Y(_00027_));
 sky130_fd_sc_hd__mux4_2 _24600_ (.A0(\w[18][6] ),
    .A1(\w[16][6] ),
    .A2(\w[22][6] ),
    .A3(\w[20][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10449_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_463 ();
 sky130_fd_sc_hd__mux4_2 _24602_ (.A0(\w[26][6] ),
    .A1(\w[24][6] ),
    .A2(\w[30][6] ),
    .A3(\w[28][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10451_));
 sky130_fd_sc_hd__mux4_2 _24603_ (.A0(\w[2][6] ),
    .A1(\w[0][6] ),
    .A2(\w[6][6] ),
    .A3(\w[4][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10452_));
 sky130_fd_sc_hd__mux4_2 _24604_ (.A0(\w[10][6] ),
    .A1(\w[8][6] ),
    .A2(\w[14][6] ),
    .A3(\w[12][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10453_));
 sky130_fd_sc_hd__mux4_2 _24605_ (.A0(_10449_),
    .A1(_10451_),
    .A2(_10452_),
    .A3(_10453_),
    .S0(net326),
    .S1(net319),
    .X(_10454_));
 sky130_fd_sc_hd__mux4_2 _24606_ (.A0(\w[50][6] ),
    .A1(\w[48][6] ),
    .A2(\w[54][6] ),
    .A3(\w[52][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10455_));
 sky130_fd_sc_hd__mux4_2 _24607_ (.A0(\w[58][6] ),
    .A1(\w[56][6] ),
    .A2(\w[62][6] ),
    .A3(\w[60][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10456_));
 sky130_fd_sc_hd__mux4_2 _24608_ (.A0(\w[34][6] ),
    .A1(\w[32][6] ),
    .A2(\w[38][6] ),
    .A3(\w[36][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_462 ();
 sky130_fd_sc_hd__mux4_2 _24610_ (.A0(\w[42][6] ),
    .A1(\w[40][6] ),
    .A2(\w[46][6] ),
    .A3(\w[44][6] ),
    .S0(net373),
    .S1(net309),
    .X(_10459_));
 sky130_fd_sc_hd__mux4_2 _24611_ (.A0(_10455_),
    .A1(_10456_),
    .A2(_10457_),
    .A3(_10459_),
    .S0(net326),
    .S1(net319),
    .X(_10460_));
 sky130_fd_sc_hd__mux2i_1 _24612_ (.A0(_10454_),
    .A1(_10460_),
    .S(net294),
    .Y(_10461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_461 ();
 sky130_fd_sc_hd__nand2_2 _24614_ (.A(net356),
    .B(\w[0][6] ),
    .Y(_10463_));
 sky130_fd_sc_hd__o21ai_4 _24615_ (.A1(net290),
    .A2(_10461_),
    .B1(_10463_),
    .Y(_00028_));
 sky130_fd_sc_hd__mux4_2 _24616_ (.A0(\w[18][7] ),
    .A1(\w[16][7] ),
    .A2(\w[22][7] ),
    .A3(\w[20][7] ),
    .S0(net375),
    .S1(net310),
    .X(_10464_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_460 ();
 sky130_fd_sc_hd__mux4_2 _24618_ (.A0(\w[26][7] ),
    .A1(\w[24][7] ),
    .A2(\w[30][7] ),
    .A3(\w[28][7] ),
    .S0(net375),
    .S1(net310),
    .X(_10466_));
 sky130_fd_sc_hd__mux4_2 _24619_ (.A0(\w[2][7] ),
    .A1(\w[0][7] ),
    .A2(\w[6][7] ),
    .A3(\w[4][7] ),
    .S0(net375),
    .S1(net310),
    .X(_10467_));
 sky130_fd_sc_hd__mux4_2 _24620_ (.A0(\w[10][7] ),
    .A1(\w[8][7] ),
    .A2(\w[14][7] ),
    .A3(\w[12][7] ),
    .S0(net375),
    .S1(net310),
    .X(_10468_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_459 ();
 sky130_fd_sc_hd__mux4_2 _24622_ (.A0(_10464_),
    .A1(_10466_),
    .A2(_10467_),
    .A3(_10468_),
    .S0(net328),
    .S1(net324),
    .X(_10470_));
 sky130_fd_sc_hd__mux4_2 _24623_ (.A0(\w[50][7] ),
    .A1(\w[48][7] ),
    .A2(\w[54][7] ),
    .A3(\w[52][7] ),
    .S0(net375),
    .S1(net309),
    .X(_10471_));
 sky130_fd_sc_hd__mux4_2 _24624_ (.A0(\w[58][7] ),
    .A1(\w[56][7] ),
    .A2(\w[62][7] ),
    .A3(\w[60][7] ),
    .S0(net375),
    .S1(net309),
    .X(_10472_));
 sky130_fd_sc_hd__mux4_2 _24625_ (.A0(\w[34][7] ),
    .A1(\w[32][7] ),
    .A2(\w[38][7] ),
    .A3(\w[36][7] ),
    .S0(net375),
    .S1(net309),
    .X(_10473_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_458 ();
 sky130_fd_sc_hd__mux4_2 _24627_ (.A0(\w[42][7] ),
    .A1(\w[40][7] ),
    .A2(\w[46][7] ),
    .A3(\w[44][7] ),
    .S0(net375),
    .S1(net309),
    .X(_10475_));
 sky130_fd_sc_hd__mux4_2 _24628_ (.A0(_10471_),
    .A1(_10472_),
    .A2(_10473_),
    .A3(_10475_),
    .S0(net327),
    .S1(net324),
    .X(_10476_));
 sky130_fd_sc_hd__mux2i_1 _24629_ (.A0(_10470_),
    .A1(_10476_),
    .S(net294),
    .Y(_10477_));
 sky130_fd_sc_hd__nand2_4 _24630_ (.A(net356),
    .B(\w[0][7] ),
    .Y(_10478_));
 sky130_fd_sc_hd__o21ai_4 _24631_ (.A1(net291),
    .A2(_10477_),
    .B1(_10478_),
    .Y(_00029_));
 sky130_fd_sc_hd__mux4_2 _24632_ (.A0(\w[18][8] ),
    .A1(\w[16][8] ),
    .A2(\w[22][8] ),
    .A3(\w[20][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10479_));
 sky130_fd_sc_hd__mux4_2 _24633_ (.A0(\w[26][8] ),
    .A1(\w[24][8] ),
    .A2(\w[30][8] ),
    .A3(\w[28][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10480_));
 sky130_fd_sc_hd__mux4_2 _24634_ (.A0(\w[2][8] ),
    .A1(\w[0][8] ),
    .A2(\w[6][8] ),
    .A3(\w[4][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10481_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_457 ();
 sky130_fd_sc_hd__mux4_2 _24636_ (.A0(\w[10][8] ),
    .A1(\w[8][8] ),
    .A2(\w[14][8] ),
    .A3(\w[12][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10483_));
 sky130_fd_sc_hd__mux4_2 _24637_ (.A0(_10479_),
    .A1(_10480_),
    .A2(_10481_),
    .A3(_10483_),
    .S0(net333),
    .S1(net322),
    .X(_10484_));
 sky130_fd_sc_hd__mux4_2 _24638_ (.A0(\w[50][8] ),
    .A1(\w[48][8] ),
    .A2(\w[54][8] ),
    .A3(\w[52][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10485_));
 sky130_fd_sc_hd__mux4_2 _24639_ (.A0(\w[58][8] ),
    .A1(\w[56][8] ),
    .A2(\w[62][8] ),
    .A3(\w[60][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10486_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_456 ();
 sky130_fd_sc_hd__mux4_2 _24641_ (.A0(\w[34][8] ),
    .A1(\w[32][8] ),
    .A2(\w[38][8] ),
    .A3(\w[36][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10488_));
 sky130_fd_sc_hd__mux4_2 _24642_ (.A0(\w[42][8] ),
    .A1(\w[40][8] ),
    .A2(\w[46][8] ),
    .A3(\w[44][8] ),
    .S0(net377),
    .S1(net312),
    .X(_10489_));
 sky130_fd_sc_hd__mux4_2 _24643_ (.A0(_10485_),
    .A1(_10486_),
    .A2(_10488_),
    .A3(_10489_),
    .S0(net329),
    .S1(net323),
    .X(_10490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_454 ();
 sky130_fd_sc_hd__mux2i_1 _24646_ (.A0(_10484_),
    .A1(_10490_),
    .S(net296),
    .Y(_10493_));
 sky130_fd_sc_hd__nand2_1 _24647_ (.A(net356),
    .B(\w[0][8] ),
    .Y(_10494_));
 sky130_fd_sc_hd__o21ai_0 _24648_ (.A1(_09875_),
    .A2(_10493_),
    .B1(_10494_),
    .Y(_00030_));
 sky130_fd_sc_hd__mux4_2 _24649_ (.A0(\w[18][9] ),
    .A1(\w[16][9] ),
    .A2(\w[22][9] ),
    .A3(\w[20][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10495_));
 sky130_fd_sc_hd__mux4_2 _24650_ (.A0(\w[26][9] ),
    .A1(\w[24][9] ),
    .A2(\w[30][9] ),
    .A3(\w[28][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10496_));
 sky130_fd_sc_hd__mux4_2 _24651_ (.A0(\w[2][9] ),
    .A1(\w[0][9] ),
    .A2(\w[6][9] ),
    .A3(\w[4][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10497_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_453 ();
 sky130_fd_sc_hd__mux4_2 _24653_ (.A0(\w[10][9] ),
    .A1(\w[8][9] ),
    .A2(\w[14][9] ),
    .A3(\w[12][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10499_));
 sky130_fd_sc_hd__mux4_2 _24654_ (.A0(_10495_),
    .A1(_10496_),
    .A2(_10497_),
    .A3(_10499_),
    .S0(net333),
    .S1(net322),
    .X(_10500_));
 sky130_fd_sc_hd__mux4_2 _24655_ (.A0(\w[50][9] ),
    .A1(\w[48][9] ),
    .A2(\w[54][9] ),
    .A3(\w[52][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10501_));
 sky130_fd_sc_hd__mux4_2 _24656_ (.A0(\w[58][9] ),
    .A1(\w[56][9] ),
    .A2(\w[62][9] ),
    .A3(\w[60][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10502_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_452 ();
 sky130_fd_sc_hd__mux4_2 _24658_ (.A0(\w[34][9] ),
    .A1(\w[32][9] ),
    .A2(\w[38][9] ),
    .A3(\w[36][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10504_));
 sky130_fd_sc_hd__mux4_2 _24659_ (.A0(\w[42][9] ),
    .A1(\w[40][9] ),
    .A2(\w[46][9] ),
    .A3(\w[44][9] ),
    .S0(net377),
    .S1(net312),
    .X(_10505_));
 sky130_fd_sc_hd__mux4_2 _24660_ (.A0(_10501_),
    .A1(_10502_),
    .A2(_10504_),
    .A3(_10505_),
    .S0(net331),
    .S1(net322),
    .X(_10506_));
 sky130_fd_sc_hd__mux2i_1 _24661_ (.A0(_10500_),
    .A1(_10506_),
    .S(net296),
    .Y(_10507_));
 sky130_fd_sc_hd__nand2_1 _24662_ (.A(net356),
    .B(\w[0][9] ),
    .Y(_10508_));
 sky130_fd_sc_hd__o21ai_0 _24663_ (.A1(_09875_),
    .A2(_10507_),
    .B1(_10508_),
    .Y(_00031_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_451 ();
 sky130_fd_sc_hd__mux4_2 _24665_ (.A0(\w[18][10] ),
    .A1(\w[16][10] ),
    .A2(\w[22][10] ),
    .A3(\w[20][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10510_));
 sky130_fd_sc_hd__mux4_2 _24666_ (.A0(\w[26][10] ),
    .A1(\w[24][10] ),
    .A2(\w[30][10] ),
    .A3(\w[28][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10511_));
 sky130_fd_sc_hd__mux4_2 _24667_ (.A0(\w[2][10] ),
    .A1(\w[0][10] ),
    .A2(\w[6][10] ),
    .A3(\w[4][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10512_));
 sky130_fd_sc_hd__mux4_2 _24668_ (.A0(\w[10][10] ),
    .A1(\w[8][10] ),
    .A2(\w[14][10] ),
    .A3(\w[12][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10513_));
 sky130_fd_sc_hd__mux4_2 _24669_ (.A0(_10510_),
    .A1(_10511_),
    .A2(_10512_),
    .A3(_10513_),
    .S0(net333),
    .S1(net322),
    .X(_10514_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_450 ();
 sky130_fd_sc_hd__mux4_2 _24671_ (.A0(\w[50][10] ),
    .A1(\w[48][10] ),
    .A2(\w[54][10] ),
    .A3(\w[52][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10516_));
 sky130_fd_sc_hd__mux4_2 _24672_ (.A0(\w[58][10] ),
    .A1(\w[56][10] ),
    .A2(\w[62][10] ),
    .A3(\w[60][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10517_));
 sky130_fd_sc_hd__mux4_2 _24673_ (.A0(\w[34][10] ),
    .A1(\w[32][10] ),
    .A2(\w[38][10] ),
    .A3(\w[36][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10518_));
 sky130_fd_sc_hd__mux4_2 _24674_ (.A0(\w[42][10] ),
    .A1(\w[40][10] ),
    .A2(\w[46][10] ),
    .A3(\w[44][10] ),
    .S0(net377),
    .S1(net312),
    .X(_10519_));
 sky130_fd_sc_hd__mux4_2 _24675_ (.A0(_10516_),
    .A1(_10517_),
    .A2(_10518_),
    .A3(_10519_),
    .S0(net331),
    .S1(net322),
    .X(_10520_));
 sky130_fd_sc_hd__mux2i_1 _24676_ (.A0(_10514_),
    .A1(_10520_),
    .S(net296),
    .Y(_10521_));
 sky130_fd_sc_hd__nand2_1 _24677_ (.A(net356),
    .B(\w[0][10] ),
    .Y(_10522_));
 sky130_fd_sc_hd__o21ai_2 _24678_ (.A1(_09875_),
    .A2(_10521_),
    .B1(_10522_),
    .Y(_00001_));
 sky130_fd_sc_hd__mux4_2 _24679_ (.A0(\w[18][11] ),
    .A1(\w[16][11] ),
    .A2(\w[22][11] ),
    .A3(\w[20][11] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10523_));
 sky130_fd_sc_hd__mux4_2 _24680_ (.A0(\w[26][11] ),
    .A1(\w[24][11] ),
    .A2(\w[30][11] ),
    .A3(\w[28][11] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10524_));
 sky130_fd_sc_hd__mux4_2 _24681_ (.A0(\w[2][11] ),
    .A1(\w[0][11] ),
    .A2(\w[6][11] ),
    .A3(\w[4][11] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10525_));
 sky130_fd_sc_hd__mux4_2 _24682_ (.A0(\w[10][11] ),
    .A1(\w[8][11] ),
    .A2(\w[14][11] ),
    .A3(\w[12][11] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10526_));
 sky130_fd_sc_hd__mux4_2 _24683_ (.A0(_10523_),
    .A1(_10524_),
    .A2(_10525_),
    .A3(_10526_),
    .S0(net330),
    .S1(net321),
    .X(_10527_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_449 ();
 sky130_fd_sc_hd__mux4_2 _24685_ (.A0(\w[50][11] ),
    .A1(\w[48][11] ),
    .A2(\w[54][11] ),
    .A3(\w[52][11] ),
    .S0(net379),
    .S1(net310),
    .X(_10529_));
 sky130_fd_sc_hd__mux4_2 _24686_ (.A0(\w[58][11] ),
    .A1(\w[56][11] ),
    .A2(\w[62][11] ),
    .A3(\w[60][11] ),
    .S0(net379),
    .S1(net310),
    .X(_10530_));
 sky130_fd_sc_hd__mux4_2 _24687_ (.A0(\w[34][11] ),
    .A1(\w[32][11] ),
    .A2(\w[38][11] ),
    .A3(\w[36][11] ),
    .S0(net379),
    .S1(net310),
    .X(_10531_));
 sky130_fd_sc_hd__mux4_2 _24688_ (.A0(\w[42][11] ),
    .A1(\w[40][11] ),
    .A2(\w[46][11] ),
    .A3(\w[44][11] ),
    .S0(net379),
    .S1(net310),
    .X(_10532_));
 sky130_fd_sc_hd__mux4_2 _24689_ (.A0(_10529_),
    .A1(_10530_),
    .A2(_10531_),
    .A3(_10532_),
    .S0(net332),
    .S1(net324),
    .X(_10533_));
 sky130_fd_sc_hd__mux2i_1 _24690_ (.A0(_10527_),
    .A1(_10533_),
    .S(net294),
    .Y(_10534_));
 sky130_fd_sc_hd__nand2_4 _24691_ (.A(net356),
    .B(\w[0][11] ),
    .Y(_10535_));
 sky130_fd_sc_hd__o21ai_4 _24692_ (.A1(net291),
    .A2(_10534_),
    .B1(_10535_),
    .Y(_00002_));
 sky130_fd_sc_hd__mux4_2 _24693_ (.A0(\w[18][12] ),
    .A1(\w[16][12] ),
    .A2(\w[22][12] ),
    .A3(\w[20][12] ),
    .S0(net375),
    .S1(net310),
    .X(_10536_));
 sky130_fd_sc_hd__mux4_2 _24694_ (.A0(\w[26][12] ),
    .A1(\w[24][12] ),
    .A2(\w[30][12] ),
    .A3(\w[28][12] ),
    .S0(net375),
    .S1(net310),
    .X(_10537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_448 ();
 sky130_fd_sc_hd__mux4_2 _24696_ (.A0(\w[2][12] ),
    .A1(\w[0][12] ),
    .A2(\w[6][12] ),
    .A3(\w[4][12] ),
    .S0(net375),
    .S1(net310),
    .X(_10539_));
 sky130_fd_sc_hd__mux4_2 _24697_ (.A0(\w[10][12] ),
    .A1(\w[8][12] ),
    .A2(\w[14][12] ),
    .A3(\w[12][12] ),
    .S0(net375),
    .S1(net310),
    .X(_10540_));
 sky130_fd_sc_hd__mux4_2 _24698_ (.A0(_10536_),
    .A1(_10537_),
    .A2(_10539_),
    .A3(_10540_),
    .S0(net328),
    .S1(net324),
    .X(_10541_));
 sky130_fd_sc_hd__mux4_2 _24699_ (.A0(\w[50][12] ),
    .A1(\w[48][12] ),
    .A2(\w[54][12] ),
    .A3(\w[52][12] ),
    .S0(net373),
    .S1(net309),
    .X(_10542_));
 sky130_fd_sc_hd__mux4_2 _24700_ (.A0(\w[58][12] ),
    .A1(\w[56][12] ),
    .A2(\w[62][12] ),
    .A3(\w[60][12] ),
    .S0(net373),
    .S1(net309),
    .X(_10543_));
 sky130_fd_sc_hd__mux4_2 _24701_ (.A0(\w[34][12] ),
    .A1(\w[32][12] ),
    .A2(\w[38][12] ),
    .A3(\w[36][12] ),
    .S0(net373),
    .S1(net309),
    .X(_10544_));
 sky130_fd_sc_hd__mux4_2 _24702_ (.A0(\w[42][12] ),
    .A1(\w[40][12] ),
    .A2(\w[46][12] ),
    .A3(\w[44][12] ),
    .S0(net373),
    .S1(net309),
    .X(_10545_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_447 ();
 sky130_fd_sc_hd__mux4_2 _24704_ (.A0(_10542_),
    .A1(_10543_),
    .A2(_10544_),
    .A3(_10545_),
    .S0(net326),
    .S1(net319),
    .X(_10547_));
 sky130_fd_sc_hd__mux2i_1 _24705_ (.A0(_10541_),
    .A1(_10547_),
    .S(net293),
    .Y(_10548_));
 sky130_fd_sc_hd__nand2_2 _24706_ (.A(net356),
    .B(\w[0][12] ),
    .Y(_10549_));
 sky130_fd_sc_hd__o21ai_4 _24707_ (.A1(net290),
    .A2(_10548_),
    .B1(_10549_),
    .Y(_00003_));
 sky130_fd_sc_hd__mux4_2 _24708_ (.A0(\w[18][13] ),
    .A1(\w[16][13] ),
    .A2(\w[22][13] ),
    .A3(\w[20][13] ),
    .S0(net375),
    .S1(net310),
    .X(_10550_));
 sky130_fd_sc_hd__mux4_2 _24709_ (.A0(\w[26][13] ),
    .A1(\w[24][13] ),
    .A2(\w[30][13] ),
    .A3(\w[28][13] ),
    .S0(net375),
    .S1(net310),
    .X(_10551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_446 ();
 sky130_fd_sc_hd__mux4_2 _24711_ (.A0(\w[2][13] ),
    .A1(\w[0][13] ),
    .A2(\w[6][13] ),
    .A3(\w[4][13] ),
    .S0(net375),
    .S1(net310),
    .X(_10553_));
 sky130_fd_sc_hd__mux4_2 _24712_ (.A0(\w[10][13] ),
    .A1(\w[8][13] ),
    .A2(\w[14][13] ),
    .A3(\w[12][13] ),
    .S0(net375),
    .S1(net310),
    .X(_10554_));
 sky130_fd_sc_hd__mux4_2 _24713_ (.A0(_10550_),
    .A1(_10551_),
    .A2(_10553_),
    .A3(_10554_),
    .S0(net328),
    .S1(net324),
    .X(_10555_));
 sky130_fd_sc_hd__mux4_2 _24714_ (.A0(\w[50][13] ),
    .A1(\w[48][13] ),
    .A2(\w[54][13] ),
    .A3(\w[52][13] ),
    .S0(net375),
    .S1(net309),
    .X(_10556_));
 sky130_fd_sc_hd__mux4_2 _24715_ (.A0(\w[58][13] ),
    .A1(\w[56][13] ),
    .A2(\w[62][13] ),
    .A3(\w[60][13] ),
    .S0(net375),
    .S1(net309),
    .X(_10557_));
 sky130_fd_sc_hd__mux4_2 _24716_ (.A0(\w[34][13] ),
    .A1(\w[32][13] ),
    .A2(\w[38][13] ),
    .A3(\w[36][13] ),
    .S0(net375),
    .S1(net309),
    .X(_10558_));
 sky130_fd_sc_hd__mux4_2 _24717_ (.A0(\w[42][13] ),
    .A1(\w[40][13] ),
    .A2(\w[46][13] ),
    .A3(\w[44][13] ),
    .S0(net375),
    .S1(net309),
    .X(_10559_));
 sky130_fd_sc_hd__mux4_2 _24718_ (.A0(_10556_),
    .A1(_10557_),
    .A2(_10558_),
    .A3(_10559_),
    .S0(net327),
    .S1(net320),
    .X(_10560_));
 sky130_fd_sc_hd__mux2i_1 _24719_ (.A0(_10555_),
    .A1(_10560_),
    .S(net293),
    .Y(_10561_));
 sky130_fd_sc_hd__nand2_2 _24720_ (.A(net356),
    .B(\w[0][13] ),
    .Y(_10562_));
 sky130_fd_sc_hd__o21ai_4 _24721_ (.A1(net290),
    .A2(_10561_),
    .B1(_10562_),
    .Y(_00004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_445 ();
 sky130_fd_sc_hd__mux4_2 _24723_ (.A0(\w[18][14] ),
    .A1(\w[16][14] ),
    .A2(\w[22][14] ),
    .A3(\w[20][14] ),
    .S0(net379),
    .S1(net310),
    .X(_10564_));
 sky130_fd_sc_hd__mux4_2 _24724_ (.A0(\w[26][14] ),
    .A1(\w[24][14] ),
    .A2(\w[30][14] ),
    .A3(\w[28][14] ),
    .S0(net379),
    .S1(net310),
    .X(_10565_));
 sky130_fd_sc_hd__mux4_2 _24725_ (.A0(\w[2][14] ),
    .A1(\w[0][14] ),
    .A2(\w[6][14] ),
    .A3(\w[4][14] ),
    .S0(net379),
    .S1(net310),
    .X(_10566_));
 sky130_fd_sc_hd__mux4_2 _24726_ (.A0(\w[10][14] ),
    .A1(\w[8][14] ),
    .A2(\w[14][14] ),
    .A3(\w[12][14] ),
    .S0(net379),
    .S1(net310),
    .X(_10567_));
 sky130_fd_sc_hd__mux4_2 _24727_ (.A0(_10564_),
    .A1(_10565_),
    .A2(_10566_),
    .A3(_10567_),
    .S0(net330),
    .S1(net321),
    .X(_10568_));
 sky130_fd_sc_hd__mux4_2 _24728_ (.A0(\w[50][14] ),
    .A1(\w[48][14] ),
    .A2(\w[54][14] ),
    .A3(\w[52][14] ),
    .S0(net375),
    .S1(net310),
    .X(_10569_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_444 ();
 sky130_fd_sc_hd__mux4_2 _24730_ (.A0(\w[58][14] ),
    .A1(\w[56][14] ),
    .A2(\w[62][14] ),
    .A3(\w[60][14] ),
    .S0(net375),
    .S1(net310),
    .X(_10571_));
 sky130_fd_sc_hd__mux4_2 _24731_ (.A0(\w[34][14] ),
    .A1(\w[32][14] ),
    .A2(\w[38][14] ),
    .A3(\w[36][14] ),
    .S0(net375),
    .S1(net310),
    .X(_10572_));
 sky130_fd_sc_hd__mux4_2 _24732_ (.A0(\w[42][14] ),
    .A1(\w[40][14] ),
    .A2(\w[46][14] ),
    .A3(\w[44][14] ),
    .S0(net375),
    .S1(net310),
    .X(_10573_));
 sky130_fd_sc_hd__mux4_2 _24733_ (.A0(_10569_),
    .A1(_10571_),
    .A2(_10572_),
    .A3(_10573_),
    .S0(net328),
    .S1(net321),
    .X(_10574_));
 sky130_fd_sc_hd__mux2i_1 _24734_ (.A0(_10568_),
    .A1(_10574_),
    .S(net293),
    .Y(_10575_));
 sky130_fd_sc_hd__nand2_2 _24735_ (.A(net356),
    .B(\w[0][14] ),
    .Y(_10576_));
 sky130_fd_sc_hd__o21ai_2 _24736_ (.A1(net290),
    .A2(_10575_),
    .B1(_10576_),
    .Y(_00005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_443 ();
 sky130_fd_sc_hd__mux4_2 _24738_ (.A0(\w[18][15] ),
    .A1(\w[16][15] ),
    .A2(\w[22][15] ),
    .A3(\w[20][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10578_));
 sky130_fd_sc_hd__mux4_2 _24739_ (.A0(\w[26][15] ),
    .A1(\w[24][15] ),
    .A2(\w[30][15] ),
    .A3(\w[28][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10579_));
 sky130_fd_sc_hd__mux4_2 _24740_ (.A0(\w[2][15] ),
    .A1(\w[0][15] ),
    .A2(\w[6][15] ),
    .A3(\w[4][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10580_));
 sky130_fd_sc_hd__mux4_2 _24741_ (.A0(\w[10][15] ),
    .A1(\w[8][15] ),
    .A2(\w[14][15] ),
    .A3(\w[12][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_442 ();
 sky130_fd_sc_hd__mux4_2 _24743_ (.A0(_10578_),
    .A1(_10579_),
    .A2(_10580_),
    .A3(_10581_),
    .S0(net327),
    .S1(net320),
    .X(_10583_));
 sky130_fd_sc_hd__mux4_2 _24744_ (.A0(\w[50][15] ),
    .A1(\w[48][15] ),
    .A2(\w[54][15] ),
    .A3(\w[52][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_441 ();
 sky130_fd_sc_hd__mux4_2 _24746_ (.A0(\w[58][15] ),
    .A1(\w[56][15] ),
    .A2(\w[62][15] ),
    .A3(\w[60][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10586_));
 sky130_fd_sc_hd__mux4_2 _24747_ (.A0(\w[34][15] ),
    .A1(\w[32][15] ),
    .A2(\w[38][15] ),
    .A3(\w[36][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10587_));
 sky130_fd_sc_hd__mux4_2 _24748_ (.A0(\w[42][15] ),
    .A1(\w[40][15] ),
    .A2(\w[46][15] ),
    .A3(\w[44][15] ),
    .S0(net374),
    .S1(net308),
    .X(_10588_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_440 ();
 sky130_fd_sc_hd__mux4_2 _24750_ (.A0(_10584_),
    .A1(_10586_),
    .A2(_10587_),
    .A3(_10588_),
    .S0(net327),
    .S1(net320),
    .X(_10590_));
 sky130_fd_sc_hd__mux2i_1 _24751_ (.A0(_10583_),
    .A1(_10590_),
    .S(net293),
    .Y(_10591_));
 sky130_fd_sc_hd__nand2_2 _24752_ (.A(net356),
    .B(\w[0][15] ),
    .Y(_10592_));
 sky130_fd_sc_hd__o21ai_4 _24753_ (.A1(net290),
    .A2(_10591_),
    .B1(_10592_),
    .Y(_00006_));
 sky130_fd_sc_hd__mux4_2 _24754_ (.A0(\w[18][16] ),
    .A1(\w[16][16] ),
    .A2(\w[22][16] ),
    .A3(\w[20][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_439 ();
 sky130_fd_sc_hd__mux4_2 _24756_ (.A0(\w[26][16] ),
    .A1(\w[24][16] ),
    .A2(\w[30][16] ),
    .A3(\w[28][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10595_));
 sky130_fd_sc_hd__mux4_2 _24757_ (.A0(\w[2][16] ),
    .A1(\w[0][16] ),
    .A2(\w[6][16] ),
    .A3(\w[4][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10596_));
 sky130_fd_sc_hd__mux4_2 _24758_ (.A0(\w[10][16] ),
    .A1(\w[8][16] ),
    .A2(\w[14][16] ),
    .A3(\w[12][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10597_));
 sky130_fd_sc_hd__mux4_2 _24759_ (.A0(_10593_),
    .A1(_10595_),
    .A2(_10596_),
    .A3(_10597_),
    .S0(net326),
    .S1(net319),
    .X(_10598_));
 sky130_fd_sc_hd__mux4_2 _24760_ (.A0(\w[50][16] ),
    .A1(\w[48][16] ),
    .A2(\w[54][16] ),
    .A3(\w[52][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10599_));
 sky130_fd_sc_hd__mux4_2 _24761_ (.A0(\w[58][16] ),
    .A1(\w[56][16] ),
    .A2(\w[62][16] ),
    .A3(\w[60][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10600_));
 sky130_fd_sc_hd__mux4_2 _24762_ (.A0(\w[34][16] ),
    .A1(\w[32][16] ),
    .A2(\w[38][16] ),
    .A3(\w[36][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10601_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_438 ();
 sky130_fd_sc_hd__mux4_2 _24764_ (.A0(\w[42][16] ),
    .A1(\w[40][16] ),
    .A2(\w[46][16] ),
    .A3(\w[44][16] ),
    .S0(net373),
    .S1(net309),
    .X(_10603_));
 sky130_fd_sc_hd__mux4_2 _24765_ (.A0(_10599_),
    .A1(_10600_),
    .A2(_10601_),
    .A3(_10603_),
    .S0(net326),
    .S1(net319),
    .X(_10604_));
 sky130_fd_sc_hd__mux2i_1 _24766_ (.A0(_10598_),
    .A1(_10604_),
    .S(net294),
    .Y(_10605_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_437 ();
 sky130_fd_sc_hd__nand2_2 _24768_ (.A(reset_hash),
    .B(\w[0][16] ),
    .Y(_10607_));
 sky130_fd_sc_hd__o21ai_4 _24769_ (.A1(net291),
    .A2(_10605_),
    .B1(_10607_),
    .Y(_00007_));
 sky130_fd_sc_hd__mux4_2 _24770_ (.A0(\w[18][17] ),
    .A1(\w[16][17] ),
    .A2(\w[22][17] ),
    .A3(\w[20][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10608_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_436 ();
 sky130_fd_sc_hd__mux4_2 _24772_ (.A0(\w[26][17] ),
    .A1(\w[24][17] ),
    .A2(\w[30][17] ),
    .A3(\w[28][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10610_));
 sky130_fd_sc_hd__mux4_2 _24773_ (.A0(\w[2][17] ),
    .A1(\w[0][17] ),
    .A2(\w[6][17] ),
    .A3(\w[4][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10611_));
 sky130_fd_sc_hd__mux4_2 _24774_ (.A0(\w[10][17] ),
    .A1(\w[8][17] ),
    .A2(\w[14][17] ),
    .A3(\w[12][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10612_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_435 ();
 sky130_fd_sc_hd__mux4_2 _24776_ (.A0(_10608_),
    .A1(_10610_),
    .A2(_10611_),
    .A3(_10612_),
    .S0(net328),
    .S1(net321),
    .X(_10614_));
 sky130_fd_sc_hd__mux4_2 _24777_ (.A0(\w[50][17] ),
    .A1(\w[48][17] ),
    .A2(\w[54][17] ),
    .A3(\w[52][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10615_));
 sky130_fd_sc_hd__mux4_2 _24778_ (.A0(\w[58][17] ),
    .A1(\w[56][17] ),
    .A2(\w[62][17] ),
    .A3(\w[60][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10616_));
 sky130_fd_sc_hd__mux4_2 _24779_ (.A0(\w[34][17] ),
    .A1(\w[32][17] ),
    .A2(\w[38][17] ),
    .A3(\w[36][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10617_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_434 ();
 sky130_fd_sc_hd__mux4_2 _24781_ (.A0(\w[42][17] ),
    .A1(\w[40][17] ),
    .A2(\w[46][17] ),
    .A3(\w[44][17] ),
    .S0(net379),
    .S1(net310),
    .X(_10619_));
 sky130_fd_sc_hd__mux4_2 _24782_ (.A0(_10615_),
    .A1(_10616_),
    .A2(_10617_),
    .A3(_10619_),
    .S0(net328),
    .S1(net321),
    .X(_10620_));
 sky130_fd_sc_hd__mux2i_1 _24783_ (.A0(_10614_),
    .A1(_10620_),
    .S(net293),
    .Y(_10621_));
 sky130_fd_sc_hd__nand2_1 _24784_ (.A(net356),
    .B(\w[0][17] ),
    .Y(_10622_));
 sky130_fd_sc_hd__o21ai_2 _24785_ (.A1(net290),
    .A2(_10621_),
    .B1(_10622_),
    .Y(_00008_));
 sky130_fd_sc_hd__mux4_2 _24786_ (.A0(\w[18][18] ),
    .A1(\w[16][18] ),
    .A2(\w[22][18] ),
    .A3(\w[20][18] ),
    .S0(net541),
    .S1(net312),
    .X(_10623_));
 sky130_fd_sc_hd__mux4_2 _24787_ (.A0(\w[26][18] ),
    .A1(\w[24][18] ),
    .A2(\w[30][18] ),
    .A3(\w[28][18] ),
    .S0(net541),
    .S1(net312),
    .X(_10624_));
 sky130_fd_sc_hd__mux4_2 _24788_ (.A0(\w[2][18] ),
    .A1(\w[0][18] ),
    .A2(\w[6][18] ),
    .A3(\w[4][18] ),
    .S0(net541),
    .S1(net312),
    .X(_10625_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_433 ();
 sky130_fd_sc_hd__mux4_2 _24790_ (.A0(\w[10][18] ),
    .A1(\w[8][18] ),
    .A2(\w[14][18] ),
    .A3(\w[12][18] ),
    .S0(net541),
    .S1(net312),
    .X(_10627_));
 sky130_fd_sc_hd__mux4_2 _24791_ (.A0(_10623_),
    .A1(_10624_),
    .A2(_10625_),
    .A3(_10627_),
    .S0(net333),
    .S1(net325),
    .X(_10628_));
 sky130_fd_sc_hd__mux4_2 _24792_ (.A0(\w[50][18] ),
    .A1(\w[48][18] ),
    .A2(\w[54][18] ),
    .A3(\w[52][18] ),
    .S0(net379),
    .S1(_00655_),
    .X(_10629_));
 sky130_fd_sc_hd__mux4_2 _24793_ (.A0(\w[58][18] ),
    .A1(\w[56][18] ),
    .A2(\w[62][18] ),
    .A3(\w[60][18] ),
    .S0(net379),
    .S1(_00655_),
    .X(_10630_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_432 ();
 sky130_fd_sc_hd__mux4_2 _24795_ (.A0(\w[34][18] ),
    .A1(\w[32][18] ),
    .A2(\w[38][18] ),
    .A3(\w[36][18] ),
    .S0(net379),
    .S1(_00655_),
    .X(_10632_));
 sky130_fd_sc_hd__mux4_2 _24796_ (.A0(\w[42][18] ),
    .A1(\w[40][18] ),
    .A2(\w[46][18] ),
    .A3(\w[44][18] ),
    .S0(net379),
    .S1(_00655_),
    .X(_10633_));
 sky130_fd_sc_hd__mux4_2 _24797_ (.A0(_10629_),
    .A1(_10630_),
    .A2(_10632_),
    .A3(_10633_),
    .S0(net332),
    .S1(net324),
    .X(_10634_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_431 ();
 sky130_fd_sc_hd__mux2i_1 _24799_ (.A0(_10628_),
    .A1(_10634_),
    .S(net296),
    .Y(_10636_));
 sky130_fd_sc_hd__nand2_1 _24800_ (.A(net540),
    .B(\w[0][18] ),
    .Y(_10637_));
 sky130_fd_sc_hd__o21ai_0 _24801_ (.A1(_09875_),
    .A2(_10636_),
    .B1(_10637_),
    .Y(_00009_));
 sky130_fd_sc_hd__mux4_2 _24802_ (.A0(\w[18][19] ),
    .A1(\w[16][19] ),
    .A2(\w[22][19] ),
    .A3(\w[20][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10638_));
 sky130_fd_sc_hd__mux4_2 _24803_ (.A0(\w[26][19] ),
    .A1(\w[24][19] ),
    .A2(\w[30][19] ),
    .A3(\w[28][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10639_));
 sky130_fd_sc_hd__mux4_2 _24804_ (.A0(\w[2][19] ),
    .A1(\w[0][19] ),
    .A2(\w[6][19] ),
    .A3(\w[4][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_430 ();
 sky130_fd_sc_hd__mux4_2 _24806_ (.A0(\w[10][19] ),
    .A1(\w[8][19] ),
    .A2(\w[14][19] ),
    .A3(\w[12][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10642_));
 sky130_fd_sc_hd__mux4_2 _24807_ (.A0(_10638_),
    .A1(_10639_),
    .A2(_10640_),
    .A3(_10642_),
    .S0(net329),
    .S1(net323),
    .X(_10643_));
 sky130_fd_sc_hd__mux4_2 _24808_ (.A0(\w[50][19] ),
    .A1(\w[48][19] ),
    .A2(\w[54][19] ),
    .A3(\w[52][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10644_));
 sky130_fd_sc_hd__mux4_2 _24809_ (.A0(\w[58][19] ),
    .A1(\w[56][19] ),
    .A2(\w[62][19] ),
    .A3(\w[60][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10645_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_429 ();
 sky130_fd_sc_hd__mux4_2 _24811_ (.A0(\w[34][19] ),
    .A1(\w[32][19] ),
    .A2(\w[38][19] ),
    .A3(\w[36][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10647_));
 sky130_fd_sc_hd__mux4_2 _24812_ (.A0(\w[42][19] ),
    .A1(\w[40][19] ),
    .A2(\w[46][19] ),
    .A3(\w[44][19] ),
    .S0(net376),
    .S1(net311),
    .X(_10648_));
 sky130_fd_sc_hd__mux4_2 _24813_ (.A0(_10644_),
    .A1(_10645_),
    .A2(_10647_),
    .A3(_10648_),
    .S0(net329),
    .S1(net323),
    .X(_10649_));
 sky130_fd_sc_hd__mux2i_1 _24814_ (.A0(_10643_),
    .A1(_10649_),
    .S(net296),
    .Y(_10650_));
 sky130_fd_sc_hd__nand2_1 _24815_ (.A(net356),
    .B(\w[0][19] ),
    .Y(_10651_));
 sky130_fd_sc_hd__o21ai_0 _24816_ (.A1(_09875_),
    .A2(_10650_),
    .B1(_10651_),
    .Y(_00010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_428 ();
 sky130_fd_sc_hd__mux4_2 _24818_ (.A0(\w[18][20] ),
    .A1(\w[16][20] ),
    .A2(\w[22][20] ),
    .A3(\w[20][20] ),
    .S0(net541),
    .S1(net312),
    .X(_10653_));
 sky130_fd_sc_hd__mux4_2 _24819_ (.A0(\w[26][20] ),
    .A1(\w[24][20] ),
    .A2(\w[30][20] ),
    .A3(\w[28][20] ),
    .S0(net541),
    .S1(net312),
    .X(_10654_));
 sky130_fd_sc_hd__mux4_2 _24820_ (.A0(\w[2][20] ),
    .A1(\w[0][20] ),
    .A2(\w[6][20] ),
    .A3(\w[4][20] ),
    .S0(net541),
    .S1(net312),
    .X(_10655_));
 sky130_fd_sc_hd__mux4_2 _24821_ (.A0(\w[10][20] ),
    .A1(\w[8][20] ),
    .A2(\w[14][20] ),
    .A3(\w[12][20] ),
    .S0(net541),
    .S1(net312),
    .X(_10656_));
 sky130_fd_sc_hd__mux4_2 _24822_ (.A0(_10653_),
    .A1(_10654_),
    .A2(_10655_),
    .A3(_10656_),
    .S0(net333),
    .S1(net322),
    .X(_10657_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_427 ();
 sky130_fd_sc_hd__mux4_2 _24824_ (.A0(\w[50][20] ),
    .A1(\w[48][20] ),
    .A2(\w[54][20] ),
    .A3(\w[52][20] ),
    .S0(net541),
    .S1(_00655_),
    .X(_10659_));
 sky130_fd_sc_hd__mux4_2 _24825_ (.A0(\w[58][20] ),
    .A1(\w[56][20] ),
    .A2(\w[62][20] ),
    .A3(\w[60][20] ),
    .S0(net541),
    .S1(_00655_),
    .X(_10660_));
 sky130_fd_sc_hd__mux4_2 _24826_ (.A0(\w[34][20] ),
    .A1(\w[32][20] ),
    .A2(\w[38][20] ),
    .A3(\w[36][20] ),
    .S0(net541),
    .S1(_00655_),
    .X(_10661_));
 sky130_fd_sc_hd__mux4_2 _24827_ (.A0(\w[42][20] ),
    .A1(\w[40][20] ),
    .A2(\w[46][20] ),
    .A3(\w[44][20] ),
    .S0(net541),
    .S1(_00655_),
    .X(_10662_));
 sky130_fd_sc_hd__mux4_2 _24828_ (.A0(_10659_),
    .A1(_10660_),
    .A2(_10661_),
    .A3(_10662_),
    .S0(net330),
    .S1(net323),
    .X(_10663_));
 sky130_fd_sc_hd__mux2i_1 _24829_ (.A0(_10657_),
    .A1(_10663_),
    .S(net296),
    .Y(_10664_));
 sky130_fd_sc_hd__nand2_1 _24830_ (.A(net356),
    .B(\w[0][20] ),
    .Y(_10665_));
 sky130_fd_sc_hd__o21ai_1 _24831_ (.A1(_09875_),
    .A2(_10664_),
    .B1(_10665_),
    .Y(_00012_));
 sky130_fd_sc_hd__mux4_2 _24832_ (.A0(\w[18][21] ),
    .A1(\w[16][21] ),
    .A2(\w[22][21] ),
    .A3(\w[20][21] ),
    .S0(net376),
    .S1(net311),
    .X(_10666_));
 sky130_fd_sc_hd__mux4_2 _24833_ (.A0(\w[26][21] ),
    .A1(\w[24][21] ),
    .A2(\w[30][21] ),
    .A3(\w[28][21] ),
    .S0(net376),
    .S1(net311),
    .X(_10667_));
 sky130_fd_sc_hd__mux4_2 _24834_ (.A0(\w[2][21] ),
    .A1(\w[0][21] ),
    .A2(\w[6][21] ),
    .A3(\w[4][21] ),
    .S0(net376),
    .S1(net311),
    .X(_10668_));
 sky130_fd_sc_hd__mux4_2 _24835_ (.A0(\w[10][21] ),
    .A1(\w[8][21] ),
    .A2(\w[14][21] ),
    .A3(\w[12][21] ),
    .S0(net376),
    .S1(net311),
    .X(_10669_));
 sky130_fd_sc_hd__mux4_2 _24836_ (.A0(_10666_),
    .A1(_10667_),
    .A2(_10668_),
    .A3(_10669_),
    .S0(net329),
    .S1(net323),
    .X(_10670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_426 ();
 sky130_fd_sc_hd__mux4_2 _24838_ (.A0(\w[50][21] ),
    .A1(\w[48][21] ),
    .A2(\w[54][21] ),
    .A3(\w[52][21] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10672_));
 sky130_fd_sc_hd__mux4_2 _24839_ (.A0(\w[58][21] ),
    .A1(\w[56][21] ),
    .A2(\w[62][21] ),
    .A3(\w[60][21] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10673_));
 sky130_fd_sc_hd__mux4_2 _24840_ (.A0(\w[34][21] ),
    .A1(\w[32][21] ),
    .A2(\w[38][21] ),
    .A3(\w[36][21] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10674_));
 sky130_fd_sc_hd__mux4_2 _24841_ (.A0(\w[42][21] ),
    .A1(\w[40][21] ),
    .A2(\w[46][21] ),
    .A3(\w[44][21] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10675_));
 sky130_fd_sc_hd__mux4_2 _24842_ (.A0(_10672_),
    .A1(_10673_),
    .A2(_10674_),
    .A3(_10675_),
    .S0(net328),
    .S1(net321),
    .X(_10676_));
 sky130_fd_sc_hd__mux2i_1 _24843_ (.A0(_10670_),
    .A1(_10676_),
    .S(net295),
    .Y(_10677_));
 sky130_fd_sc_hd__nand2_4 _24844_ (.A(net356),
    .B(\w[0][21] ),
    .Y(_10678_));
 sky130_fd_sc_hd__o21ai_0 _24845_ (.A1(net291),
    .A2(_10677_),
    .B1(_10678_),
    .Y(_00013_));
 sky130_fd_sc_hd__mux4_2 _24846_ (.A0(\w[18][22] ),
    .A1(\w[16][22] ),
    .A2(\w[22][22] ),
    .A3(\w[20][22] ),
    .S0(net377),
    .S1(net312),
    .X(_10679_));
 sky130_fd_sc_hd__mux4_2 _24847_ (.A0(\w[26][22] ),
    .A1(\w[24][22] ),
    .A2(\w[30][22] ),
    .A3(\w[28][22] ),
    .S0(net377),
    .S1(net312),
    .X(_10680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_425 ();
 sky130_fd_sc_hd__mux4_2 _24849_ (.A0(\w[2][22] ),
    .A1(\w[0][22] ),
    .A2(\w[6][22] ),
    .A3(\w[4][22] ),
    .S0(net377),
    .S1(net312),
    .X(_10682_));
 sky130_fd_sc_hd__mux4_2 _24850_ (.A0(\w[10][22] ),
    .A1(\w[8][22] ),
    .A2(\w[14][22] ),
    .A3(\w[12][22] ),
    .S0(net377),
    .S1(net312),
    .X(_10683_));
 sky130_fd_sc_hd__mux4_2 _24851_ (.A0(_10679_),
    .A1(_10680_),
    .A2(_10682_),
    .A3(_10683_),
    .S0(net333),
    .S1(net322),
    .X(_10684_));
 sky130_fd_sc_hd__mux4_2 _24852_ (.A0(\w[50][22] ),
    .A1(\w[48][22] ),
    .A2(\w[54][22] ),
    .A3(\w[52][22] ),
    .S0(net541),
    .S1(net312),
    .X(_10685_));
 sky130_fd_sc_hd__mux4_2 _24853_ (.A0(\w[58][22] ),
    .A1(\w[56][22] ),
    .A2(\w[62][22] ),
    .A3(\w[60][22] ),
    .S0(net541),
    .S1(net312),
    .X(_10686_));
 sky130_fd_sc_hd__mux4_2 _24854_ (.A0(\w[34][22] ),
    .A1(\w[32][22] ),
    .A2(\w[38][22] ),
    .A3(\w[36][22] ),
    .S0(net541),
    .S1(net312),
    .X(_10687_));
 sky130_fd_sc_hd__mux4_2 _24855_ (.A0(\w[42][22] ),
    .A1(\w[40][22] ),
    .A2(\w[46][22] ),
    .A3(\w[44][22] ),
    .S0(net541),
    .S1(net312),
    .X(_10688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_424 ();
 sky130_fd_sc_hd__mux4_2 _24857_ (.A0(_10685_),
    .A1(_10686_),
    .A2(_10687_),
    .A3(_10688_),
    .S0(net331),
    .S1(net322),
    .X(_10690_));
 sky130_fd_sc_hd__mux2i_1 _24858_ (.A0(_10684_),
    .A1(_10690_),
    .S(net296),
    .Y(_10691_));
 sky130_fd_sc_hd__nand2_1 _24859_ (.A(net356),
    .B(\w[0][22] ),
    .Y(_10692_));
 sky130_fd_sc_hd__o21ai_0 _24860_ (.A1(_09875_),
    .A2(_10691_),
    .B1(_10692_),
    .Y(_00014_));
 sky130_fd_sc_hd__mux4_2 _24861_ (.A0(\w[18][23] ),
    .A1(\w[16][23] ),
    .A2(\w[22][23] ),
    .A3(\w[20][23] ),
    .S0(net379),
    .S1(net310),
    .X(_10693_));
 sky130_fd_sc_hd__mux4_2 _24862_ (.A0(\w[26][23] ),
    .A1(\w[24][23] ),
    .A2(\w[30][23] ),
    .A3(\w[28][23] ),
    .S0(net379),
    .S1(net310),
    .X(_10694_));
 sky130_fd_sc_hd__mux4_2 _24863_ (.A0(\w[2][23] ),
    .A1(\w[0][23] ),
    .A2(\w[6][23] ),
    .A3(\w[4][23] ),
    .S0(net379),
    .S1(net310),
    .X(_10695_));
 sky130_fd_sc_hd__mux4_2 _24864_ (.A0(\w[10][23] ),
    .A1(\w[8][23] ),
    .A2(\w[14][23] ),
    .A3(\w[12][23] ),
    .S0(net379),
    .S1(net310),
    .X(_10696_));
 sky130_fd_sc_hd__mux4_2 _24865_ (.A0(_10693_),
    .A1(_10694_),
    .A2(_10695_),
    .A3(_10696_),
    .S0(net330),
    .S1(net324),
    .X(_10697_));
 sky130_fd_sc_hd__mux4_2 _24866_ (.A0(\w[50][23] ),
    .A1(\w[48][23] ),
    .A2(\w[54][23] ),
    .A3(\w[52][23] ),
    .S0(net375),
    .S1(net308),
    .X(_10698_));
 sky130_fd_sc_hd__mux4_2 _24867_ (.A0(\w[58][23] ),
    .A1(\w[56][23] ),
    .A2(\w[62][23] ),
    .A3(\w[60][23] ),
    .S0(net375),
    .S1(net310),
    .X(_10699_));
 sky130_fd_sc_hd__mux4_2 _24868_ (.A0(\w[34][23] ),
    .A1(\w[32][23] ),
    .A2(\w[38][23] ),
    .A3(\w[36][23] ),
    .S0(net375),
    .S1(net308),
    .X(_10700_));
 sky130_fd_sc_hd__mux4_2 _24869_ (.A0(\w[42][23] ),
    .A1(\w[40][23] ),
    .A2(\w[46][23] ),
    .A3(\w[44][23] ),
    .S0(net375),
    .S1(net310),
    .X(_10701_));
 sky130_fd_sc_hd__mux4_2 _24870_ (.A0(_10698_),
    .A1(_10699_),
    .A2(_10700_),
    .A3(_10701_),
    .S0(net328),
    .S1(net324),
    .X(_10702_));
 sky130_fd_sc_hd__mux2i_1 _24871_ (.A0(_10697_),
    .A1(_10702_),
    .S(net293),
    .Y(_10703_));
 sky130_fd_sc_hd__nand2_4 _24872_ (.A(net356),
    .B(\w[0][23] ),
    .Y(_10704_));
 sky130_fd_sc_hd__o21ai_4 _24873_ (.A1(net290),
    .A2(_10703_),
    .B1(_10704_),
    .Y(_00015_));
 sky130_fd_sc_hd__mux4_2 _24874_ (.A0(\w[18][24] ),
    .A1(\w[16][24] ),
    .A2(\w[22][24] ),
    .A3(\w[20][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10705_));
 sky130_fd_sc_hd__mux4_2 _24875_ (.A0(\w[26][24] ),
    .A1(\w[24][24] ),
    .A2(\w[30][24] ),
    .A3(\w[28][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10706_));
 sky130_fd_sc_hd__mux4_2 _24876_ (.A0(\w[2][24] ),
    .A1(\w[0][24] ),
    .A2(\w[6][24] ),
    .A3(\w[4][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10707_));
 sky130_fd_sc_hd__mux4_2 _24877_ (.A0(\w[10][24] ),
    .A1(\w[8][24] ),
    .A2(\w[14][24] ),
    .A3(\w[12][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10708_));
 sky130_fd_sc_hd__mux4_2 _24878_ (.A0(_10705_),
    .A1(_10706_),
    .A2(_10707_),
    .A3(_10708_),
    .S0(net329),
    .S1(net323),
    .X(_10709_));
 sky130_fd_sc_hd__mux4_2 _24879_ (.A0(\w[50][24] ),
    .A1(\w[48][24] ),
    .A2(\w[54][24] ),
    .A3(\w[52][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10710_));
 sky130_fd_sc_hd__mux4_2 _24880_ (.A0(\w[58][24] ),
    .A1(\w[56][24] ),
    .A2(\w[62][24] ),
    .A3(\w[60][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10711_));
 sky130_fd_sc_hd__mux4_2 _24881_ (.A0(\w[34][24] ),
    .A1(\w[32][24] ),
    .A2(\w[38][24] ),
    .A3(\w[36][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10712_));
 sky130_fd_sc_hd__mux4_2 _24882_ (.A0(\w[42][24] ),
    .A1(\w[40][24] ),
    .A2(\w[46][24] ),
    .A3(\w[44][24] ),
    .S0(net376),
    .S1(net311),
    .X(_10713_));
 sky130_fd_sc_hd__mux4_2 _24883_ (.A0(_10710_),
    .A1(_10711_),
    .A2(_10712_),
    .A3(_10713_),
    .S0(net329),
    .S1(net323),
    .X(_10714_));
 sky130_fd_sc_hd__mux2i_1 _24884_ (.A0(_10709_),
    .A1(_10714_),
    .S(net296),
    .Y(_10715_));
 sky130_fd_sc_hd__nand2_1 _24885_ (.A(net356),
    .B(\w[0][24] ),
    .Y(_10716_));
 sky130_fd_sc_hd__o21ai_2 _24886_ (.A1(_09875_),
    .A2(_10715_),
    .B1(_10716_),
    .Y(_00016_));
 sky130_fd_sc_hd__mux4_2 _24887_ (.A0(\w[18][25] ),
    .A1(\w[16][25] ),
    .A2(\w[22][25] ),
    .A3(\w[20][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10717_));
 sky130_fd_sc_hd__mux4_2 _24888_ (.A0(\w[26][25] ),
    .A1(\w[24][25] ),
    .A2(\w[30][25] ),
    .A3(\w[28][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10718_));
 sky130_fd_sc_hd__mux4_2 _24889_ (.A0(\w[2][25] ),
    .A1(\w[0][25] ),
    .A2(\w[6][25] ),
    .A3(\w[4][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10719_));
 sky130_fd_sc_hd__mux4_2 _24890_ (.A0(\w[10][25] ),
    .A1(\w[8][25] ),
    .A2(\w[14][25] ),
    .A3(\w[12][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10720_));
 sky130_fd_sc_hd__mux4_2 _24891_ (.A0(_10717_),
    .A1(_10718_),
    .A2(_10719_),
    .A3(_10720_),
    .S0(net330),
    .S1(net321),
    .X(_10721_));
 sky130_fd_sc_hd__mux4_2 _24892_ (.A0(\w[50][25] ),
    .A1(\w[48][25] ),
    .A2(\w[54][25] ),
    .A3(\w[52][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10722_));
 sky130_fd_sc_hd__mux4_2 _24893_ (.A0(\w[58][25] ),
    .A1(\w[56][25] ),
    .A2(\w[62][25] ),
    .A3(\w[60][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10723_));
 sky130_fd_sc_hd__mux4_2 _24894_ (.A0(\w[34][25] ),
    .A1(\w[32][25] ),
    .A2(\w[38][25] ),
    .A3(\w[36][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10724_));
 sky130_fd_sc_hd__mux4_2 _24895_ (.A0(\w[42][25] ),
    .A1(\w[40][25] ),
    .A2(\w[46][25] ),
    .A3(\w[44][25] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_423 ();
 sky130_fd_sc_hd__mux4_2 _24897_ (.A0(_10722_),
    .A1(_10723_),
    .A2(_10724_),
    .A3(_10725_),
    .S0(net330),
    .S1(net321),
    .X(_10727_));
 sky130_fd_sc_hd__mux2i_1 _24898_ (.A0(_10721_),
    .A1(_10727_),
    .S(net295),
    .Y(_10728_));
 sky130_fd_sc_hd__nand2_1 _24899_ (.A(net356),
    .B(\w[0][25] ),
    .Y(_10729_));
 sky130_fd_sc_hd__o21ai_2 _24900_ (.A1(net291),
    .A2(_10728_),
    .B1(_10729_),
    .Y(_00017_));
 sky130_fd_sc_hd__mux4_2 _24901_ (.A0(\w[18][26] ),
    .A1(\w[16][26] ),
    .A2(\w[22][26] ),
    .A3(\w[20][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10730_));
 sky130_fd_sc_hd__mux4_2 _24902_ (.A0(\w[26][26] ),
    .A1(\w[24][26] ),
    .A2(\w[30][26] ),
    .A3(\w[28][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10731_));
 sky130_fd_sc_hd__mux4_2 _24903_ (.A0(\w[2][26] ),
    .A1(\w[0][26] ),
    .A2(\w[6][26] ),
    .A3(\w[4][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10732_));
 sky130_fd_sc_hd__mux4_2 _24904_ (.A0(\w[10][26] ),
    .A1(\w[8][26] ),
    .A2(\w[14][26] ),
    .A3(\w[12][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10733_));
 sky130_fd_sc_hd__mux4_2 _24905_ (.A0(_10730_),
    .A1(_10731_),
    .A2(_10732_),
    .A3(_10733_),
    .S0(net329),
    .S1(net323),
    .X(_10734_));
 sky130_fd_sc_hd__mux4_2 _24906_ (.A0(\w[50][26] ),
    .A1(\w[48][26] ),
    .A2(\w[54][26] ),
    .A3(\w[52][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10735_));
 sky130_fd_sc_hd__mux4_2 _24907_ (.A0(\w[58][26] ),
    .A1(\w[56][26] ),
    .A2(\w[62][26] ),
    .A3(\w[60][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10736_));
 sky130_fd_sc_hd__mux4_2 _24908_ (.A0(\w[34][26] ),
    .A1(\w[32][26] ),
    .A2(\w[38][26] ),
    .A3(\w[36][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10737_));
 sky130_fd_sc_hd__mux4_2 _24909_ (.A0(\w[42][26] ),
    .A1(\w[40][26] ),
    .A2(\w[46][26] ),
    .A3(\w[44][26] ),
    .S0(net376),
    .S1(net311),
    .X(_10738_));
 sky130_fd_sc_hd__mux4_2 _24910_ (.A0(_10735_),
    .A1(_10736_),
    .A2(_10737_),
    .A3(_10738_),
    .S0(net329),
    .S1(net323),
    .X(_10739_));
 sky130_fd_sc_hd__mux2i_1 _24911_ (.A0(_10734_),
    .A1(_10739_),
    .S(net295),
    .Y(_10740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_422 ();
 sky130_fd_sc_hd__nand2_1 _24913_ (.A(net356),
    .B(\w[0][26] ),
    .Y(_10742_));
 sky130_fd_sc_hd__o21ai_0 _24914_ (.A1(_09875_),
    .A2(_10740_),
    .B1(_10742_),
    .Y(_00018_));
 sky130_fd_sc_hd__mux4_2 _24915_ (.A0(\w[18][27] ),
    .A1(\w[16][27] ),
    .A2(\w[22][27] ),
    .A3(\w[20][27] ),
    .S0(net375),
    .S1(net310),
    .X(_10743_));
 sky130_fd_sc_hd__mux4_2 _24916_ (.A0(\w[26][27] ),
    .A1(\w[24][27] ),
    .A2(\w[30][27] ),
    .A3(\w[28][27] ),
    .S0(net375),
    .S1(net310),
    .X(_10744_));
 sky130_fd_sc_hd__mux4_2 _24917_ (.A0(\w[2][27] ),
    .A1(\w[0][27] ),
    .A2(\w[6][27] ),
    .A3(\w[4][27] ),
    .S0(net375),
    .S1(net310),
    .X(_10745_));
 sky130_fd_sc_hd__mux4_2 _24918_ (.A0(\w[10][27] ),
    .A1(\w[8][27] ),
    .A2(\w[14][27] ),
    .A3(\w[12][27] ),
    .S0(net375),
    .S1(net310),
    .X(_10746_));
 sky130_fd_sc_hd__mux4_2 _24919_ (.A0(_10743_),
    .A1(_10744_),
    .A2(_10745_),
    .A3(_10746_),
    .S0(net328),
    .S1(net324),
    .X(_10747_));
 sky130_fd_sc_hd__mux4_2 _24920_ (.A0(\w[50][27] ),
    .A1(\w[48][27] ),
    .A2(\w[54][27] ),
    .A3(\w[52][27] ),
    .S0(net375),
    .S1(net308),
    .X(_10748_));
 sky130_fd_sc_hd__mux4_2 _24921_ (.A0(\w[58][27] ),
    .A1(\w[56][27] ),
    .A2(\w[62][27] ),
    .A3(\w[60][27] ),
    .S0(net375),
    .S1(net308),
    .X(_10749_));
 sky130_fd_sc_hd__mux4_2 _24922_ (.A0(\w[34][27] ),
    .A1(\w[32][27] ),
    .A2(\w[38][27] ),
    .A3(\w[36][27] ),
    .S0(net375),
    .S1(net308),
    .X(_10750_));
 sky130_fd_sc_hd__mux4_2 _24923_ (.A0(\w[42][27] ),
    .A1(\w[40][27] ),
    .A2(\w[46][27] ),
    .A3(\w[44][27] ),
    .S0(net375),
    .S1(net308),
    .X(_10751_));
 sky130_fd_sc_hd__mux4_2 _24924_ (.A0(_10748_),
    .A1(_10749_),
    .A2(_10750_),
    .A3(_10751_),
    .S0(net328),
    .S1(net324),
    .X(_10752_));
 sky130_fd_sc_hd__mux2i_1 _24925_ (.A0(_10747_),
    .A1(_10752_),
    .S(net293),
    .Y(_10753_));
 sky130_fd_sc_hd__nand2_4 _24926_ (.A(net356),
    .B(\w[0][27] ),
    .Y(_10754_));
 sky130_fd_sc_hd__o21ai_4 _24927_ (.A1(net290),
    .A2(_10753_),
    .B1(_10754_),
    .Y(_00019_));
 sky130_fd_sc_hd__mux4_2 _24928_ (.A0(\w[18][28] ),
    .A1(\w[16][28] ),
    .A2(\w[22][28] ),
    .A3(\w[20][28] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10755_));
 sky130_fd_sc_hd__mux4_2 _24929_ (.A0(\w[26][28] ),
    .A1(\w[24][28] ),
    .A2(\w[30][28] ),
    .A3(\w[28][28] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10756_));
 sky130_fd_sc_hd__mux4_2 _24930_ (.A0(\w[2][28] ),
    .A1(\w[0][28] ),
    .A2(\w[6][28] ),
    .A3(\w[4][28] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10757_));
 sky130_fd_sc_hd__mux4_2 _24931_ (.A0(\w[10][28] ),
    .A1(\w[8][28] ),
    .A2(\w[14][28] ),
    .A3(\w[12][28] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10758_));
 sky130_fd_sc_hd__mux4_2 _24932_ (.A0(_10755_),
    .A1(_10756_),
    .A2(_10757_),
    .A3(_10758_),
    .S0(net330),
    .S1(net321),
    .X(_10759_));
 sky130_fd_sc_hd__mux4_2 _24933_ (.A0(\w[50][28] ),
    .A1(\w[48][28] ),
    .A2(\w[54][28] ),
    .A3(\w[52][28] ),
    .S0(net379),
    .S1(net310),
    .X(_10760_));
 sky130_fd_sc_hd__mux4_2 _24934_ (.A0(\w[58][28] ),
    .A1(\w[56][28] ),
    .A2(\w[62][28] ),
    .A3(\w[60][28] ),
    .S0(net379),
    .S1(net310),
    .X(_10761_));
 sky130_fd_sc_hd__mux4_2 _24935_ (.A0(\w[34][28] ),
    .A1(\w[32][28] ),
    .A2(\w[38][28] ),
    .A3(\w[36][28] ),
    .S0(net379),
    .S1(net310),
    .X(_10762_));
 sky130_fd_sc_hd__mux4_2 _24936_ (.A0(\w[42][28] ),
    .A1(\w[40][28] ),
    .A2(\w[46][28] ),
    .A3(\w[44][28] ),
    .S0(net379),
    .S1(net310),
    .X(_10763_));
 sky130_fd_sc_hd__mux4_2 _24937_ (.A0(_10760_),
    .A1(_10761_),
    .A2(_10762_),
    .A3(_10763_),
    .S0(net328),
    .S1(net321),
    .X(_10764_));
 sky130_fd_sc_hd__mux2i_1 _24938_ (.A0(_10759_),
    .A1(_10764_),
    .S(net293),
    .Y(_10765_));
 sky130_fd_sc_hd__nand2_4 _24939_ (.A(net356),
    .B(\w[0][28] ),
    .Y(_10766_));
 sky130_fd_sc_hd__o21ai_2 _24940_ (.A1(net290),
    .A2(_10765_),
    .B1(_10766_),
    .Y(_00020_));
 sky130_fd_sc_hd__mux4_2 _24941_ (.A0(\w[18][29] ),
    .A1(\w[16][29] ),
    .A2(\w[22][29] ),
    .A3(\w[20][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10767_));
 sky130_fd_sc_hd__mux4_2 _24942_ (.A0(\w[26][29] ),
    .A1(\w[24][29] ),
    .A2(\w[30][29] ),
    .A3(\w[28][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10768_));
 sky130_fd_sc_hd__mux4_2 _24943_ (.A0(\w[2][29] ),
    .A1(\w[0][29] ),
    .A2(\w[6][29] ),
    .A3(\w[4][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10769_));
 sky130_fd_sc_hd__mux4_2 _24944_ (.A0(\w[10][29] ),
    .A1(\w[8][29] ),
    .A2(\w[14][29] ),
    .A3(\w[12][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10770_));
 sky130_fd_sc_hd__mux4_2 _24945_ (.A0(_10767_),
    .A1(_10768_),
    .A2(_10769_),
    .A3(_10770_),
    .S0(net327),
    .S1(net320),
    .X(_10771_));
 sky130_fd_sc_hd__mux4_2 _24946_ (.A0(\w[50][29] ),
    .A1(\w[48][29] ),
    .A2(\w[54][29] ),
    .A3(\w[52][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10772_));
 sky130_fd_sc_hd__mux4_2 _24947_ (.A0(\w[58][29] ),
    .A1(\w[56][29] ),
    .A2(\w[62][29] ),
    .A3(\w[60][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10773_));
 sky130_fd_sc_hd__mux4_2 _24948_ (.A0(\w[34][29] ),
    .A1(\w[32][29] ),
    .A2(\w[38][29] ),
    .A3(\w[36][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10774_));
 sky130_fd_sc_hd__mux4_2 _24949_ (.A0(\w[42][29] ),
    .A1(\w[40][29] ),
    .A2(\w[46][29] ),
    .A3(\w[44][29] ),
    .S0(net374),
    .S1(net308),
    .X(_10775_));
 sky130_fd_sc_hd__mux4_2 _24950_ (.A0(_10772_),
    .A1(_10773_),
    .A2(_10774_),
    .A3(_10775_),
    .S0(net327),
    .S1(net320),
    .X(_10776_));
 sky130_fd_sc_hd__mux2i_1 _24951_ (.A0(_10771_),
    .A1(_10776_),
    .S(net293),
    .Y(_10777_));
 sky130_fd_sc_hd__nand2_2 _24952_ (.A(net356),
    .B(\w[0][29] ),
    .Y(_10778_));
 sky130_fd_sc_hd__o21ai_4 _24953_ (.A1(net290),
    .A2(_10777_),
    .B1(_10778_),
    .Y(_00021_));
 sky130_fd_sc_hd__mux4_2 _24954_ (.A0(\w[18][30] ),
    .A1(\w[16][30] ),
    .A2(\w[22][30] ),
    .A3(\w[20][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10779_));
 sky130_fd_sc_hd__mux4_2 _24955_ (.A0(\w[26][30] ),
    .A1(\w[24][30] ),
    .A2(\w[30][30] ),
    .A3(\w[28][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10780_));
 sky130_fd_sc_hd__mux4_2 _24956_ (.A0(\w[2][30] ),
    .A1(\w[0][30] ),
    .A2(\w[6][30] ),
    .A3(\w[4][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10781_));
 sky130_fd_sc_hd__mux4_2 _24957_ (.A0(\w[10][30] ),
    .A1(\w[8][30] ),
    .A2(\w[14][30] ),
    .A3(\w[12][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10782_));
 sky130_fd_sc_hd__mux4_2 _24958_ (.A0(_10779_),
    .A1(_10780_),
    .A2(_10781_),
    .A3(_10782_),
    .S0(net327),
    .S1(net320),
    .X(_10783_));
 sky130_fd_sc_hd__mux4_2 _24959_ (.A0(\w[50][30] ),
    .A1(\w[48][30] ),
    .A2(\w[54][30] ),
    .A3(\w[52][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10784_));
 sky130_fd_sc_hd__mux4_2 _24960_ (.A0(\w[58][30] ),
    .A1(\w[56][30] ),
    .A2(\w[62][30] ),
    .A3(\w[60][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10785_));
 sky130_fd_sc_hd__mux4_2 _24961_ (.A0(\w[34][30] ),
    .A1(\w[32][30] ),
    .A2(\w[38][30] ),
    .A3(\w[36][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10786_));
 sky130_fd_sc_hd__mux4_2 _24962_ (.A0(\w[42][30] ),
    .A1(\w[40][30] ),
    .A2(\w[46][30] ),
    .A3(\w[44][30] ),
    .S0(net374),
    .S1(net308),
    .X(_10787_));
 sky130_fd_sc_hd__mux4_2 _24963_ (.A0(_10784_),
    .A1(_10785_),
    .A2(_10786_),
    .A3(_10787_),
    .S0(net326),
    .S1(net319),
    .X(_10788_));
 sky130_fd_sc_hd__mux2i_1 _24964_ (.A0(_10783_),
    .A1(_10788_),
    .S(net293),
    .Y(_10789_));
 sky130_fd_sc_hd__nand2_2 _24965_ (.A(net356),
    .B(\w[0][30] ),
    .Y(_10790_));
 sky130_fd_sc_hd__o21ai_4 _24966_ (.A1(net290),
    .A2(_10789_),
    .B1(_10790_),
    .Y(_00023_));
 sky130_fd_sc_hd__mux4_2 _24967_ (.A0(\w[18][31] ),
    .A1(\w[16][31] ),
    .A2(\w[22][31] ),
    .A3(\w[20][31] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10791_));
 sky130_fd_sc_hd__mux4_2 _24968_ (.A0(\w[26][31] ),
    .A1(\w[24][31] ),
    .A2(\w[30][31] ),
    .A3(\w[28][31] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10792_));
 sky130_fd_sc_hd__mux4_2 _24969_ (.A0(\w[2][31] ),
    .A1(\w[0][31] ),
    .A2(\w[6][31] ),
    .A3(\w[4][31] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10793_));
 sky130_fd_sc_hd__mux4_2 _24970_ (.A0(\w[10][31] ),
    .A1(\w[8][31] ),
    .A2(\w[14][31] ),
    .A3(\w[12][31] ),
    .S0(net378),
    .S1(_00655_),
    .X(_10794_));
 sky130_fd_sc_hd__mux4_2 _24971_ (.A0(_10791_),
    .A1(_10792_),
    .A2(_10793_),
    .A3(_10794_),
    .S0(net328),
    .S1(net321),
    .X(_10795_));
 sky130_fd_sc_hd__mux4_2 _24972_ (.A0(\w[50][31] ),
    .A1(\w[48][31] ),
    .A2(\w[54][31] ),
    .A3(\w[52][31] ),
    .S0(net379),
    .S1(net310),
    .X(_10796_));
 sky130_fd_sc_hd__mux4_2 _24973_ (.A0(\w[58][31] ),
    .A1(\w[56][31] ),
    .A2(\w[62][31] ),
    .A3(\w[60][31] ),
    .S0(net379),
    .S1(net310),
    .X(_10797_));
 sky130_fd_sc_hd__mux4_2 _24974_ (.A0(\w[34][31] ),
    .A1(\w[32][31] ),
    .A2(\w[38][31] ),
    .A3(\w[36][31] ),
    .S0(net379),
    .S1(_00655_),
    .X(_10798_));
 sky130_fd_sc_hd__mux4_2 _24975_ (.A0(\w[42][31] ),
    .A1(\w[40][31] ),
    .A2(\w[46][31] ),
    .A3(\w[44][31] ),
    .S0(net379),
    .S1(_00655_),
    .X(_10799_));
 sky130_fd_sc_hd__mux4_2 _24976_ (.A0(_10796_),
    .A1(_10797_),
    .A2(_10798_),
    .A3(_10799_),
    .S0(net327),
    .S1(net324),
    .X(_10800_));
 sky130_fd_sc_hd__mux2i_1 _24977_ (.A0(_10795_),
    .A1(_10800_),
    .S(net293),
    .Y(_10801_));
 sky130_fd_sc_hd__nand2_1 _24978_ (.A(net356),
    .B(\w[0][31] ),
    .Y(_10802_));
 sky130_fd_sc_hd__o21ai_2 _24979_ (.A1(net290),
    .A2(_10801_),
    .B1(_10802_),
    .Y(_00024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_413 ();
 sky130_fd_sc_hd__mux4_2 _24989_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10812_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_409 ();
 sky130_fd_sc_hd__mux4_2 _24994_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10817_));
 sky130_fd_sc_hd__mux4_2 _24995_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10818_));
 sky130_fd_sc_hd__mux4_2 _24996_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_404 ();
 sky130_fd_sc_hd__mux4_2 _25002_ (.A0(_10812_),
    .A1(_10817_),
    .A2(_10818_),
    .A3(_10819_),
    .S0(net522),
    .S1(net521),
    .X(_10825_));
 sky130_fd_sc_hd__mux4_2 _25003_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10826_));
 sky130_fd_sc_hd__mux4_2 _25004_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10827_));
 sky130_fd_sc_hd__mux4_2 _25005_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10828_));
 sky130_fd_sc_hd__mux4_2 _25006_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net525),
    .S1(net536),
    .X(_10829_));
 sky130_fd_sc_hd__mux4_2 _25007_ (.A0(_10826_),
    .A1(_10827_),
    .A2(_10828_),
    .A3(_10829_),
    .S0(net524),
    .S1(net521),
    .X(_10830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_402 ();
 sky130_fd_sc_hd__mux2i_4 _25010_ (.A0(_10825_),
    .A1(_10830_),
    .S(net558),
    .Y(_10833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__mux4_2 _25014_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net531),
    .S1(net533),
    .X(_10837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_397 ();
 sky130_fd_sc_hd__mux4_2 _25017_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net531),
    .S1(net533),
    .X(_10840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_395 ();
 sky130_fd_sc_hd__mux4_2 _25020_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net531),
    .S1(net535),
    .X(_10843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_393 ();
 sky130_fd_sc_hd__mux4_2 _25023_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net531),
    .S1(net535),
    .X(_10846_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_391 ();
 sky130_fd_sc_hd__mux4_2 _25026_ (.A0(_10837_),
    .A1(_10840_),
    .A2(_10843_),
    .A3(_10846_),
    .S0(net523),
    .S1(net559),
    .X(_10849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__mux4_2 _25028_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net531),
    .S1(net533),
    .X(_10851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__mux4_2 _25031_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net531),
    .S1(net533),
    .X(_10854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__mux4_2 _25034_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net531),
    .S1(net533),
    .X(_10857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__mux4_2 _25037_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net531),
    .S1(net533),
    .X(_10860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__mux4_2 _25040_ (.A0(_10851_),
    .A1(_10854_),
    .A2(_10857_),
    .A3(_10860_),
    .S0(net523),
    .S1(net559),
    .X(_10863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__mux2i_4 _25042_ (.A0(_10849_),
    .A1(_10863_),
    .S(net519),
    .Y(_10865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_379 ();
 sky130_fd_sc_hd__mux4_2 _25045_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_10868_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_377 ();
 sky130_fd_sc_hd__mux4_2 _25048_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_10871_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_376 ();
 sky130_fd_sc_hd__mux4_2 _25050_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_10873_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__mux4_2 _25052_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_10875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__mux4_2 _25055_ (.A0(_10868_),
    .A1(_10871_),
    .A2(_10873_),
    .A3(_10875_),
    .S0(net524),
    .S1(net521),
    .X(_10878_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__mux4_2 _25058_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net529),
    .S1(net537),
    .X(_10881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__mux4_2 _25061_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net529),
    .S1(net537),
    .X(_10884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_368 ();
 sky130_fd_sc_hd__mux4_2 _25063_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net529),
    .S1(net537),
    .X(_10886_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_366 ();
 sky130_fd_sc_hd__mux4_2 _25066_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net529),
    .S1(net537),
    .X(_10889_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_364 ();
 sky130_fd_sc_hd__mux4_2 _25069_ (.A0(_10881_),
    .A1(_10884_),
    .A2(_10886_),
    .A3(_10889_),
    .S0(\count15_1[3] ),
    .S1(net520),
    .X(_10892_));
 sky130_fd_sc_hd__mux2i_4 _25070_ (.A0(_10878_),
    .A1(_10892_),
    .S(net518),
    .Y(_10893_));
 sky130_fd_sc_hd__xnor2_1 _25071_ (.A(_10865_),
    .B(_10893_),
    .Y(_10894_));
 sky130_fd_sc_hd__xnor2_1 _25072_ (.A(_10833_),
    .B(_10894_),
    .Y(_11579_));
 sky130_fd_sc_hd__mux4_2 _25073_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net526),
    .S1(net534),
    .X(_10895_));
 sky130_fd_sc_hd__mux4_2 _25074_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net526),
    .S1(net534),
    .X(_10896_));
 sky130_fd_sc_hd__mux4_2 _25075_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net526),
    .S1(net534),
    .X(_10897_));
 sky130_fd_sc_hd__mux4_2 _25076_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net526),
    .S1(net534),
    .X(_10898_));
 sky130_fd_sc_hd__mux4_2 _25077_ (.A0(_10895_),
    .A1(_10896_),
    .A2(_10897_),
    .A3(_10898_),
    .S0(net522),
    .S1(net520),
    .X(_10899_));
 sky130_fd_sc_hd__mux4_2 _25078_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net528),
    .S1(net534),
    .X(_10900_));
 sky130_fd_sc_hd__mux4_2 _25079_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net528),
    .S1(net534),
    .X(_10901_));
 sky130_fd_sc_hd__mux4_2 _25080_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net528),
    .S1(net534),
    .X(_10902_));
 sky130_fd_sc_hd__mux4_2 _25081_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net528),
    .S1(net534),
    .X(_10903_));
 sky130_fd_sc_hd__mux4_2 _25082_ (.A0(_10900_),
    .A1(_10901_),
    .A2(_10902_),
    .A3(_10903_),
    .S0(net522),
    .S1(net520),
    .X(_10904_));
 sky130_fd_sc_hd__mux2i_4 _25083_ (.A0(_10899_),
    .A1(_10904_),
    .S(net518),
    .Y(_10905_));
 sky130_fd_sc_hd__mux4_2 _25084_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net527),
    .S1(net533),
    .X(_10906_));
 sky130_fd_sc_hd__mux4_2 _25085_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net527),
    .S1(net533),
    .X(_10907_));
 sky130_fd_sc_hd__mux4_2 _25086_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net527),
    .S1(net533),
    .X(_10908_));
 sky130_fd_sc_hd__mux4_2 _25087_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net527),
    .S1(net533),
    .X(_10909_));
 sky130_fd_sc_hd__mux4_2 _25088_ (.A0(_10906_),
    .A1(_10907_),
    .A2(_10908_),
    .A3(_10909_),
    .S0(net522),
    .S1(net520),
    .X(_10910_));
 sky130_fd_sc_hd__mux4_2 _25089_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net529),
    .S1(net535),
    .X(_10911_));
 sky130_fd_sc_hd__mux4_2 _25090_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net529),
    .S1(net535),
    .X(_10912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_363 ();
 sky130_fd_sc_hd__mux4_2 _25092_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net529),
    .S1(net535),
    .X(_10914_));
 sky130_fd_sc_hd__mux4_2 _25093_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net529),
    .S1(net535),
    .X(_10915_));
 sky130_fd_sc_hd__mux4_2 _25094_ (.A0(_10911_),
    .A1(_10912_),
    .A2(_10914_),
    .A3(_10915_),
    .S0(\count15_1[3] ),
    .S1(net520),
    .X(_10916_));
 sky130_fd_sc_hd__mux2i_4 _25095_ (.A0(_10910_),
    .A1(_10916_),
    .S(net518),
    .Y(_10917_));
 sky130_fd_sc_hd__mux4_2 _25096_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net527),
    .S1(net533),
    .X(_10918_));
 sky130_fd_sc_hd__mux4_2 _25097_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net527),
    .S1(net533),
    .X(_10919_));
 sky130_fd_sc_hd__mux4_2 _25098_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net527),
    .S1(net533),
    .X(_10920_));
 sky130_fd_sc_hd__mux4_2 _25099_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net527),
    .S1(net533),
    .X(_10921_));
 sky130_fd_sc_hd__mux4_2 _25100_ (.A0(_10918_),
    .A1(_10919_),
    .A2(_10920_),
    .A3(_10921_),
    .S0(net523),
    .S1(net520),
    .X(_10922_));
 sky130_fd_sc_hd__mux4_2 _25101_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net531),
    .S1(net535),
    .X(_10923_));
 sky130_fd_sc_hd__mux4_2 _25102_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net531),
    .S1(net535),
    .X(_10924_));
 sky130_fd_sc_hd__mux4_2 _25103_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net531),
    .S1(net535),
    .X(_10925_));
 sky130_fd_sc_hd__mux4_2 _25104_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net531),
    .S1(net535),
    .X(_10926_));
 sky130_fd_sc_hd__mux4_2 _25105_ (.A0(_10923_),
    .A1(_10924_),
    .A2(_10925_),
    .A3(_10926_),
    .S0(net523),
    .S1(net559),
    .X(_10927_));
 sky130_fd_sc_hd__mux2i_4 _25106_ (.A0(_10922_),
    .A1(_10927_),
    .S(net519),
    .Y(_10928_));
 sky130_fd_sc_hd__xnor2_1 _25107_ (.A(_10917_),
    .B(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__xnor2_1 _25108_ (.A(_10905_),
    .B(_10929_),
    .Y(_11584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 ();
 sky130_fd_sc_hd__mux4_2 _25119_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net444),
    .S1(net451),
    .X(_10940_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_351 ();
 sky130_fd_sc_hd__mux4_2 _25122_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net444),
    .S1(net451),
    .X(_10943_));
 sky130_fd_sc_hd__mux4_2 _25123_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net444),
    .S1(net451),
    .X(_10944_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_349 ();
 sky130_fd_sc_hd__mux4_2 _25126_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net444),
    .S1(net451),
    .X(_10947_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 ();
 sky130_fd_sc_hd__mux4_2 _25132_ (.A0(_10940_),
    .A1(_10943_),
    .A2(_10944_),
    .A3(_10947_),
    .S0(net442),
    .S1(net440),
    .X(_10953_));
 sky130_fd_sc_hd__mux4_2 _25133_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net450),
    .S1(net455),
    .X(_10954_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_342 ();
 sky130_fd_sc_hd__mux4_2 _25136_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net450),
    .S1(net455),
    .X(_10957_));
 sky130_fd_sc_hd__mux4_2 _25137_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net450),
    .S1(net455),
    .X(_10958_));
 sky130_fd_sc_hd__mux4_2 _25138_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net450),
    .S1(net455),
    .X(_10959_));
 sky130_fd_sc_hd__mux4_2 _25139_ (.A0(_10954_),
    .A1(_10957_),
    .A2(_10958_),
    .A3(_10959_),
    .S0(net441),
    .S1(net439),
    .X(_10960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_340 ();
 sky130_fd_sc_hd__mux2i_4 _25142_ (.A0(_10953_),
    .A1(_10960_),
    .S(net438),
    .Y(_10963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_337 ();
 sky130_fd_sc_hd__mux4_2 _25146_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net447),
    .S1(net453),
    .X(_10967_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_335 ();
 sky130_fd_sc_hd__mux4_2 _25149_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net447),
    .S1(net453),
    .X(_10970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_333 ();
 sky130_fd_sc_hd__mux4_2 _25152_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net447),
    .S1(net453),
    .X(_10973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_331 ();
 sky130_fd_sc_hd__mux4_2 _25155_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net447),
    .S1(net453),
    .X(_10976_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_329 ();
 sky130_fd_sc_hd__mux4_2 _25158_ (.A0(_10967_),
    .A1(_10970_),
    .A2(_10973_),
    .A3(_10976_),
    .S0(net441),
    .S1(net439),
    .X(_10979_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_327 ();
 sky130_fd_sc_hd__mux4_2 _25161_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net450),
    .S1(net455),
    .X(_10982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_326 ();
 sky130_fd_sc_hd__mux4_2 _25163_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net450),
    .S1(net455),
    .X(_10984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_324 ();
 sky130_fd_sc_hd__mux4_2 _25166_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net450),
    .S1(net455),
    .X(_10987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_322 ();
 sky130_fd_sc_hd__mux4_2 _25169_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net450),
    .S1(net455),
    .X(_10990_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_320 ();
 sky130_fd_sc_hd__mux4_2 _25172_ (.A0(_10982_),
    .A1(_10984_),
    .A2(_10987_),
    .A3(_10990_),
    .S0(net441),
    .S1(net439),
    .X(_10993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_319 ();
 sky130_fd_sc_hd__mux2i_4 _25174_ (.A0(_10979_),
    .A1(_10993_),
    .S(net438),
    .Y(_10995_));
 sky130_fd_sc_hd__mux4_2 _25175_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net449),
    .S1(net455),
    .X(_10996_));
 sky130_fd_sc_hd__mux4_2 _25176_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net449),
    .S1(net455),
    .X(_10997_));
 sky130_fd_sc_hd__mux4_2 _25177_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net449),
    .S1(net455),
    .X(_10998_));
 sky130_fd_sc_hd__mux4_2 _25178_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net449),
    .S1(net455),
    .X(_10999_));
 sky130_fd_sc_hd__mux4_2 _25179_ (.A0(_10996_),
    .A1(_10997_),
    .A2(_10998_),
    .A3(_10999_),
    .S0(net441),
    .S1(net439),
    .X(_11000_));
 sky130_fd_sc_hd__mux4_2 _25180_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net450),
    .S1(net455),
    .X(_11001_));
 sky130_fd_sc_hd__mux4_2 _25181_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net450),
    .S1(net455),
    .X(_11002_));
 sky130_fd_sc_hd__mux4_2 _25182_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net450),
    .S1(net455),
    .X(_11003_));
 sky130_fd_sc_hd__mux4_2 _25183_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net450),
    .S1(net455),
    .X(_11004_));
 sky130_fd_sc_hd__mux4_2 _25184_ (.A0(_11001_),
    .A1(_11002_),
    .A2(_11003_),
    .A3(_11004_),
    .S0(net441),
    .S1(net439),
    .X(_11005_));
 sky130_fd_sc_hd__mux2i_4 _25185_ (.A0(_11000_),
    .A1(_11005_),
    .S(net438),
    .Y(_11006_));
 sky130_fd_sc_hd__xnor2_1 _25186_ (.A(_10995_),
    .B(_11006_),
    .Y(_11007_));
 sky130_fd_sc_hd__xnor2_1 _25187_ (.A(_10963_),
    .B(_11007_),
    .Y(_11589_));
 sky130_fd_sc_hd__mux4_2 _25188_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_318 ();
 sky130_fd_sc_hd__mux4_2 _25190_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11010_));
 sky130_fd_sc_hd__mux4_2 _25191_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11011_));
 sky130_fd_sc_hd__mux4_2 _25192_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11012_));
 sky130_fd_sc_hd__mux4_2 _25193_ (.A0(_11008_),
    .A1(_11010_),
    .A2(_11011_),
    .A3(_11012_),
    .S0(net523),
    .S1(net559),
    .X(_11013_));
 sky130_fd_sc_hd__mux4_2 _25194_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11014_));
 sky130_fd_sc_hd__mux4_2 _25195_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_317 ();
 sky130_fd_sc_hd__mux4_2 _25197_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_315 ();
 sky130_fd_sc_hd__mux4_2 _25200_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net532),
    .S1(net537),
    .X(_11020_));
 sky130_fd_sc_hd__mux4_2 _25201_ (.A0(_11014_),
    .A1(_11015_),
    .A2(_11017_),
    .A3(_11020_),
    .S0(net523),
    .S1(net559),
    .X(_11021_));
 sky130_fd_sc_hd__mux2i_4 _25202_ (.A0(_11013_),
    .A1(_11021_),
    .S(net519),
    .Y(_11022_));
 sky130_fd_sc_hd__mux4_2 _25203_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11023_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_314 ();
 sky130_fd_sc_hd__mux4_2 _25205_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11025_));
 sky130_fd_sc_hd__mux4_2 _25206_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11026_));
 sky130_fd_sc_hd__mux4_2 _25207_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11027_));
 sky130_fd_sc_hd__mux4_2 _25208_ (.A0(_11023_),
    .A1(_11025_),
    .A2(_11026_),
    .A3(_11027_),
    .S0(net524),
    .S1(net521),
    .X(_11028_));
 sky130_fd_sc_hd__mux4_2 _25209_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11029_));
 sky130_fd_sc_hd__mux4_2 _25210_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11030_));
 sky130_fd_sc_hd__mux4_2 _25211_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11031_));
 sky130_fd_sc_hd__mux4_2 _25212_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net525),
    .S1(net536),
    .X(_11032_));
 sky130_fd_sc_hd__mux4_2 _25213_ (.A0(_11029_),
    .A1(_11030_),
    .A2(_11031_),
    .A3(_11032_),
    .S0(net524),
    .S1(net521),
    .X(_11033_));
 sky130_fd_sc_hd__mux2i_4 _25214_ (.A0(_11028_),
    .A1(_11033_),
    .S(net558),
    .Y(_11034_));
 sky130_fd_sc_hd__mux4_2 _25215_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11035_));
 sky130_fd_sc_hd__mux4_2 _25216_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11036_));
 sky130_fd_sc_hd__mux4_2 _25217_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11037_));
 sky130_fd_sc_hd__mux4_2 _25218_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11038_));
 sky130_fd_sc_hd__mux4_2 _25219_ (.A0(_11035_),
    .A1(_11036_),
    .A2(_11037_),
    .A3(_11038_),
    .S0(net523),
    .S1(net559),
    .X(_11039_));
 sky130_fd_sc_hd__mux4_2 _25220_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11040_));
 sky130_fd_sc_hd__mux4_2 _25221_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11041_));
 sky130_fd_sc_hd__mux4_2 _25222_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11042_));
 sky130_fd_sc_hd__mux4_2 _25223_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net532),
    .S1(net537),
    .X(_11043_));
 sky130_fd_sc_hd__mux4_2 _25224_ (.A0(_11040_),
    .A1(_11041_),
    .A2(_11042_),
    .A3(_11043_),
    .S0(net523),
    .S1(net559),
    .X(_11044_));
 sky130_fd_sc_hd__mux2i_4 _25225_ (.A0(_11039_),
    .A1(_11044_),
    .S(net519),
    .Y(_11045_));
 sky130_fd_sc_hd__xnor2_1 _25226_ (.A(_11034_),
    .B(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__xnor2_1 _25227_ (.A(_11022_),
    .B(_11046_),
    .Y(_11592_));
 sky130_fd_sc_hd__mux4_2 _25228_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net444),
    .S1(net451),
    .X(_11047_));
 sky130_fd_sc_hd__mux4_2 _25229_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net444),
    .S1(net451),
    .X(_11048_));
 sky130_fd_sc_hd__mux4_2 _25230_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net444),
    .S1(net451),
    .X(_11049_));
 sky130_fd_sc_hd__mux4_2 _25231_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net444),
    .S1(net451),
    .X(_11050_));
 sky130_fd_sc_hd__mux4_2 _25232_ (.A0(_11047_),
    .A1(_11048_),
    .A2(_11049_),
    .A3(_11050_),
    .S0(net443),
    .S1(net550),
    .X(_11051_));
 sky130_fd_sc_hd__mux4_2 _25233_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net450),
    .S1(net456),
    .X(_11052_));
 sky130_fd_sc_hd__mux4_2 _25234_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net450),
    .S1(net456),
    .X(_11053_));
 sky130_fd_sc_hd__mux4_2 _25235_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net450),
    .S1(net456),
    .X(_11054_));
 sky130_fd_sc_hd__mux4_2 _25236_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net450),
    .S1(net456),
    .X(_11055_));
 sky130_fd_sc_hd__mux4_2 _25237_ (.A0(_11052_),
    .A1(_11053_),
    .A2(_11054_),
    .A3(_11055_),
    .S0(net442),
    .S1(net440),
    .X(_11056_));
 sky130_fd_sc_hd__mux2i_4 _25238_ (.A0(_11051_),
    .A1(_11056_),
    .S(net438),
    .Y(_11057_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_313 ();
 sky130_fd_sc_hd__mux4_2 _25240_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net444),
    .S1(net451),
    .X(_11059_));
 sky130_fd_sc_hd__mux4_2 _25241_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net444),
    .S1(net451),
    .X(_11060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_312 ();
 sky130_fd_sc_hd__mux4_2 _25243_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net444),
    .S1(net451),
    .X(_11062_));
 sky130_fd_sc_hd__mux4_2 _25244_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net444),
    .S1(net451),
    .X(_11063_));
 sky130_fd_sc_hd__mux4_2 _25245_ (.A0(_11059_),
    .A1(_11060_),
    .A2(_11062_),
    .A3(_11063_),
    .S0(net442),
    .S1(net440),
    .X(_11064_));
 sky130_fd_sc_hd__mux4_2 _25246_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net448),
    .S1(net454),
    .X(_11065_));
 sky130_fd_sc_hd__mux4_2 _25247_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net448),
    .S1(net454),
    .X(_11066_));
 sky130_fd_sc_hd__mux4_2 _25248_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net449),
    .S1(net455),
    .X(_11067_));
 sky130_fd_sc_hd__mux4_2 _25249_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net449),
    .S1(net455),
    .X(_11068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_311 ();
 sky130_fd_sc_hd__mux4_2 _25251_ (.A0(_11065_),
    .A1(_11066_),
    .A2(_11067_),
    .A3(_11068_),
    .S0(net441),
    .S1(net439),
    .X(_11070_));
 sky130_fd_sc_hd__mux2i_4 _25252_ (.A0(_11064_),
    .A1(_11070_),
    .S(net437),
    .Y(_11071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_310 ();
 sky130_fd_sc_hd__mux4_2 _25254_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net448),
    .S1(net454),
    .X(_11073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_309 ();
 sky130_fd_sc_hd__mux4_2 _25256_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net448),
    .S1(net454),
    .X(_11075_));
 sky130_fd_sc_hd__mux4_2 _25257_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net448),
    .S1(net454),
    .X(_11076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_307 ();
 sky130_fd_sc_hd__mux4_2 _25260_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net448),
    .S1(net454),
    .X(_11079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_305 ();
 sky130_fd_sc_hd__mux4_2 _25263_ (.A0(_11073_),
    .A1(_11075_),
    .A2(_11076_),
    .A3(_11079_),
    .S0(net442),
    .S1(net440),
    .X(_11082_));
 sky130_fd_sc_hd__mux4_2 _25264_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net447),
    .S1(net453),
    .X(_11083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_303 ();
 sky130_fd_sc_hd__mux4_2 _25267_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net448),
    .S1(net454),
    .X(_11086_));
 sky130_fd_sc_hd__mux4_2 _25268_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net448),
    .S1(net454),
    .X(_11087_));
 sky130_fd_sc_hd__mux4_2 _25269_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net448),
    .S1(net454),
    .X(_11088_));
 sky130_fd_sc_hd__mux4_2 _25270_ (.A0(_11083_),
    .A1(_11086_),
    .A2(_11087_),
    .A3(_11088_),
    .S0(net441),
    .S1(net439),
    .X(_11089_));
 sky130_fd_sc_hd__mux2i_4 _25271_ (.A0(_11082_),
    .A1(_11089_),
    .S(net437),
    .Y(_11090_));
 sky130_fd_sc_hd__xnor2_1 _25272_ (.A(_11071_),
    .B(_11090_),
    .Y(_11091_));
 sky130_fd_sc_hd__xnor2_1 _25273_ (.A(_11057_),
    .B(_11091_),
    .Y(_11597_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_301 ();
 sky130_fd_sc_hd__mux4_2 _25276_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_11094_));
 sky130_fd_sc_hd__mux4_2 _25277_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_11095_));
 sky130_fd_sc_hd__mux4_2 _25278_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_11096_));
 sky130_fd_sc_hd__mux4_2 _25279_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_11097_));
 sky130_fd_sc_hd__mux4_2 _25280_ (.A0(_11094_),
    .A1(_11095_),
    .A2(_11096_),
    .A3(_11097_),
    .S0(net524),
    .S1(net521),
    .X(_11098_));
 sky130_fd_sc_hd__mux4_2 _25281_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net530),
    .S1(net537),
    .X(_11099_));
 sky130_fd_sc_hd__mux4_2 _25282_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net530),
    .S1(net537),
    .X(_11100_));
 sky130_fd_sc_hd__mux4_2 _25283_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(\count15_1[2] ),
    .S1(net537),
    .X(_11101_));
 sky130_fd_sc_hd__mux4_2 _25284_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(\count15_1[2] ),
    .S1(net537),
    .X(_11102_));
 sky130_fd_sc_hd__mux4_2 _25285_ (.A0(_11099_),
    .A1(_11100_),
    .A2(_11101_),
    .A3(_11102_),
    .S0(net524),
    .S1(net521),
    .X(_11103_));
 sky130_fd_sc_hd__mux2i_4 _25286_ (.A0(_11098_),
    .A1(_11103_),
    .S(net558),
    .Y(_11104_));
 sky130_fd_sc_hd__mux4_2 _25287_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11105_));
 sky130_fd_sc_hd__mux4_2 _25288_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11106_));
 sky130_fd_sc_hd__mux4_2 _25289_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11107_));
 sky130_fd_sc_hd__mux4_2 _25290_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11108_));
 sky130_fd_sc_hd__mux4_2 _25291_ (.A0(_11105_),
    .A1(_11106_),
    .A2(_11107_),
    .A3(_11108_),
    .S0(net523),
    .S1(net559),
    .X(_11109_));
 sky130_fd_sc_hd__mux4_2 _25292_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11110_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_300 ();
 sky130_fd_sc_hd__mux4_2 _25294_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11112_));
 sky130_fd_sc_hd__mux4_2 _25295_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11113_));
 sky130_fd_sc_hd__mux4_2 _25296_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net531),
    .S1(net535),
    .X(_11114_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_299 ();
 sky130_fd_sc_hd__mux4_2 _25298_ (.A0(_11110_),
    .A1(_11112_),
    .A2(_11113_),
    .A3(_11114_),
    .S0(net523),
    .S1(net559),
    .X(_11116_));
 sky130_fd_sc_hd__mux2i_4 _25299_ (.A0(_11109_),
    .A1(_11116_),
    .S(net519),
    .Y(_11117_));
 sky130_fd_sc_hd__mux4_2 _25300_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net531),
    .S1(net535),
    .X(_11118_));
 sky130_fd_sc_hd__mux4_2 _25301_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net531),
    .S1(net535),
    .X(_11119_));
 sky130_fd_sc_hd__mux4_2 _25302_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net531),
    .S1(net535),
    .X(_11120_));
 sky130_fd_sc_hd__mux4_2 _25303_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net531),
    .S1(net535),
    .X(_11121_));
 sky130_fd_sc_hd__mux4_2 _25304_ (.A0(_11118_),
    .A1(_11119_),
    .A2(_11120_),
    .A3(_11121_),
    .S0(net523),
    .S1(net559),
    .X(_11122_));
 sky130_fd_sc_hd__mux4_2 _25305_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net531),
    .S1(net537),
    .X(_11123_));
 sky130_fd_sc_hd__mux4_2 _25306_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net531),
    .S1(net537),
    .X(_11124_));
 sky130_fd_sc_hd__mux4_2 _25307_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net531),
    .S1(net537),
    .X(_11125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_298 ();
 sky130_fd_sc_hd__mux4_2 _25309_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net531),
    .S1(net537),
    .X(_11127_));
 sky130_fd_sc_hd__mux4_2 _25310_ (.A0(_11123_),
    .A1(_11124_),
    .A2(_11125_),
    .A3(_11127_),
    .S0(net523),
    .S1(net559),
    .X(_11128_));
 sky130_fd_sc_hd__mux2i_4 _25311_ (.A0(_11122_),
    .A1(_11128_),
    .S(net519),
    .Y(_11129_));
 sky130_fd_sc_hd__xnor2_1 _25312_ (.A(_11117_),
    .B(_11129_),
    .Y(_11130_));
 sky130_fd_sc_hd__xnor2_1 _25313_ (.A(_11104_),
    .B(_11130_),
    .Y(_11603_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_297 ();
 sky130_fd_sc_hd__mux4_2 _25315_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net444),
    .S1(net451),
    .X(_11132_));
 sky130_fd_sc_hd__mux4_2 _25316_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net444),
    .S1(net451),
    .X(_11133_));
 sky130_fd_sc_hd__mux4_2 _25317_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net444),
    .S1(net451),
    .X(_11134_));
 sky130_fd_sc_hd__mux4_2 _25318_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net444),
    .S1(net451),
    .X(_11135_));
 sky130_fd_sc_hd__mux4_2 _25319_ (.A0(_11132_),
    .A1(_11133_),
    .A2(_11134_),
    .A3(_11135_),
    .S0(net443),
    .S1(net550),
    .X(_11136_));
 sky130_fd_sc_hd__mux4_2 _25320_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net450),
    .S1(net456),
    .X(_11137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_295 ();
 sky130_fd_sc_hd__mux4_2 _25323_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net450),
    .S1(net456),
    .X(_11140_));
 sky130_fd_sc_hd__mux4_2 _25324_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net450),
    .S1(net456),
    .X(_11141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_294 ();
 sky130_fd_sc_hd__mux4_2 _25326_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net450),
    .S1(net456),
    .X(_11143_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_293 ();
 sky130_fd_sc_hd__mux4_2 _25328_ (.A0(_11137_),
    .A1(_11140_),
    .A2(_11141_),
    .A3(_11143_),
    .S0(net442),
    .S1(net440),
    .X(_11145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_292 ();
 sky130_fd_sc_hd__mux2i_4 _25330_ (.A0(_11136_),
    .A1(_11145_),
    .S(net438),
    .Y(_11147_));
 sky130_fd_sc_hd__mux4_2 _25331_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net447),
    .S1(net453),
    .X(_11148_));
 sky130_fd_sc_hd__mux4_2 _25332_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net447),
    .S1(net453),
    .X(_11149_));
 sky130_fd_sc_hd__mux4_2 _25333_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net447),
    .S1(net453),
    .X(_11150_));
 sky130_fd_sc_hd__mux4_2 _25334_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net447),
    .S1(net453),
    .X(_11151_));
 sky130_fd_sc_hd__mux4_2 _25335_ (.A0(_11148_),
    .A1(_11149_),
    .A2(_11150_),
    .A3(_11151_),
    .S0(net441),
    .S1(net439),
    .X(_11152_));
 sky130_fd_sc_hd__mux4_2 _25336_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net449),
    .S1(net455),
    .X(_11153_));
 sky130_fd_sc_hd__mux4_2 _25337_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net449),
    .S1(net455),
    .X(_11154_));
 sky130_fd_sc_hd__mux4_2 _25338_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net449),
    .S1(net455),
    .X(_11155_));
 sky130_fd_sc_hd__mux4_2 _25339_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net449),
    .S1(net455),
    .X(_11156_));
 sky130_fd_sc_hd__mux4_2 _25340_ (.A0(_11153_),
    .A1(_11154_),
    .A2(_11155_),
    .A3(_11156_),
    .S0(net441),
    .S1(net439),
    .X(_11157_));
 sky130_fd_sc_hd__mux2i_4 _25341_ (.A0(_11152_),
    .A1(_11157_),
    .S(net437),
    .Y(_11158_));
 sky130_fd_sc_hd__xnor2_1 _25342_ (.A(_11147_),
    .B(_11158_),
    .Y(_11159_));
 sky130_fd_sc_hd__xnor2_1 _25343_ (.A(_10995_),
    .B(_11159_),
    .Y(_11608_));
 sky130_fd_sc_hd__mux4_2 _25344_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net531),
    .S1(net533),
    .X(_11160_));
 sky130_fd_sc_hd__mux4_2 _25345_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net531),
    .S1(net533),
    .X(_11161_));
 sky130_fd_sc_hd__mux4_2 _25346_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net531),
    .S1(net533),
    .X(_11162_));
 sky130_fd_sc_hd__mux4_2 _25347_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net531),
    .S1(net533),
    .X(_11163_));
 sky130_fd_sc_hd__mux4_2 _25348_ (.A0(_11160_),
    .A1(_11161_),
    .A2(_11162_),
    .A3(_11163_),
    .S0(net523),
    .S1(net559),
    .X(_11164_));
 sky130_fd_sc_hd__mux4_2 _25349_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net527),
    .S1(net533),
    .X(_11165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_291 ();
 sky130_fd_sc_hd__mux4_2 _25351_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net527),
    .S1(net533),
    .X(_11167_));
 sky130_fd_sc_hd__mux4_2 _25352_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net527),
    .S1(net533),
    .X(_11168_));
 sky130_fd_sc_hd__mux4_2 _25353_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net527),
    .S1(net533),
    .X(_11169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_290 ();
 sky130_fd_sc_hd__mux4_2 _25355_ (.A0(_11165_),
    .A1(_11167_),
    .A2(_11168_),
    .A3(_11169_),
    .S0(net522),
    .S1(net520),
    .X(_11171_));
 sky130_fd_sc_hd__mux2i_4 _25356_ (.A0(_11164_),
    .A1(_11171_),
    .S(net518),
    .Y(_11172_));
 sky130_fd_sc_hd__mux4_2 _25357_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net527),
    .S1(net533),
    .X(_11173_));
 sky130_fd_sc_hd__mux4_2 _25358_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net527),
    .S1(net533),
    .X(_11174_));
 sky130_fd_sc_hd__mux4_2 _25359_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net527),
    .S1(net533),
    .X(_11175_));
 sky130_fd_sc_hd__mux4_2 _25360_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net527),
    .S1(net533),
    .X(_11176_));
 sky130_fd_sc_hd__mux4_2 _25361_ (.A0(_11173_),
    .A1(_11174_),
    .A2(_11175_),
    .A3(_11176_),
    .S0(net523),
    .S1(net559),
    .X(_11177_));
 sky130_fd_sc_hd__mux4_2 _25362_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net532),
    .S1(net537),
    .X(_11178_));
 sky130_fd_sc_hd__mux4_2 _25363_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net532),
    .S1(net537),
    .X(_11179_));
 sky130_fd_sc_hd__mux4_2 _25364_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net532),
    .S1(net537),
    .X(_11180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_289 ();
 sky130_fd_sc_hd__mux4_2 _25366_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net532),
    .S1(net537),
    .X(_11182_));
 sky130_fd_sc_hd__mux4_2 _25367_ (.A0(_11178_),
    .A1(_11179_),
    .A2(_11180_),
    .A3(_11182_),
    .S0(net523),
    .S1(net559),
    .X(_11183_));
 sky130_fd_sc_hd__mux2i_4 _25368_ (.A0(_11177_),
    .A1(_11183_),
    .S(net519),
    .Y(_11184_));
 sky130_fd_sc_hd__xnor2_1 _25369_ (.A(_11172_),
    .B(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__xnor2_1 _25370_ (.A(_10893_),
    .B(_11185_),
    .Y(_11611_));
 sky130_fd_sc_hd__mux4_2 _25371_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net444),
    .S1(net451),
    .X(_11186_));
 sky130_fd_sc_hd__mux4_2 _25372_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net444),
    .S1(net451),
    .X(_11187_));
 sky130_fd_sc_hd__mux4_2 _25373_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net444),
    .S1(net451),
    .X(_11188_));
 sky130_fd_sc_hd__mux4_2 _25374_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net444),
    .S1(net451),
    .X(_11189_));
 sky130_fd_sc_hd__mux4_2 _25375_ (.A0(_11186_),
    .A1(_11187_),
    .A2(_11188_),
    .A3(_11189_),
    .S0(net443),
    .S1(net550),
    .X(_11190_));
 sky130_fd_sc_hd__mux4_2 _25376_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net450),
    .S1(net455),
    .X(_11191_));
 sky130_fd_sc_hd__mux4_2 _25377_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net450),
    .S1(net456),
    .X(_11192_));
 sky130_fd_sc_hd__mux4_2 _25378_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net450),
    .S1(net456),
    .X(_11193_));
 sky130_fd_sc_hd__mux4_2 _25379_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net450),
    .S1(net456),
    .X(_11194_));
 sky130_fd_sc_hd__mux4_2 _25380_ (.A0(_11191_),
    .A1(_11192_),
    .A2(_11193_),
    .A3(_11194_),
    .S0(net442),
    .S1(net440),
    .X(_11195_));
 sky130_fd_sc_hd__mux2i_4 _25381_ (.A0(_11190_),
    .A1(_11195_),
    .S(net437),
    .Y(_11196_));
 sky130_fd_sc_hd__mux4_2 _25382_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net444),
    .S1(net451),
    .X(_11197_));
 sky130_fd_sc_hd__mux4_2 _25383_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net444),
    .S1(net451),
    .X(_11198_));
 sky130_fd_sc_hd__mux4_2 _25384_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net444),
    .S1(net451),
    .X(_11199_));
 sky130_fd_sc_hd__mux4_2 _25385_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net444),
    .S1(net451),
    .X(_11200_));
 sky130_fd_sc_hd__mux4_2 _25386_ (.A0(_11197_),
    .A1(_11198_),
    .A2(_11199_),
    .A3(_11200_),
    .S0(net443),
    .S1(net550),
    .X(_11201_));
 sky130_fd_sc_hd__mux4_2 _25387_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net445),
    .S1(net451),
    .X(_11202_));
 sky130_fd_sc_hd__mux4_2 _25388_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net445),
    .S1(net451),
    .X(_11203_));
 sky130_fd_sc_hd__mux4_2 _25389_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net445),
    .S1(net451),
    .X(_11204_));
 sky130_fd_sc_hd__mux4_2 _25390_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net445),
    .S1(net451),
    .X(_11205_));
 sky130_fd_sc_hd__mux4_2 _25391_ (.A0(_11202_),
    .A1(_11203_),
    .A2(_11204_),
    .A3(_11205_),
    .S0(net443),
    .S1(net550),
    .X(_11206_));
 sky130_fd_sc_hd__mux2i_4 _25392_ (.A0(_11201_),
    .A1(_11206_),
    .S(net438),
    .Y(_11207_));
 sky130_fd_sc_hd__xnor2_1 _25393_ (.A(_11196_),
    .B(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__xnor2_1 _25394_ (.A(_11071_),
    .B(_11208_),
    .Y(_11616_));
 sky130_fd_sc_hd__mux4_2 _25395_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net530),
    .S1(net560),
    .X(_11209_));
 sky130_fd_sc_hd__mux4_2 _25396_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net530),
    .S1(net560),
    .X(_11210_));
 sky130_fd_sc_hd__mux4_2 _25397_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net530),
    .S1(net560),
    .X(_11211_));
 sky130_fd_sc_hd__mux4_2 _25398_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net530),
    .S1(net560),
    .X(_11212_));
 sky130_fd_sc_hd__mux4_2 _25399_ (.A0(_11209_),
    .A1(_11210_),
    .A2(_11211_),
    .A3(_11212_),
    .S0(net524),
    .S1(net521),
    .X(_11213_));
 sky130_fd_sc_hd__mux4_2 _25400_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net529),
    .S1(net535),
    .X(_11214_));
 sky130_fd_sc_hd__mux4_2 _25401_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net529),
    .S1(net535),
    .X(_11215_));
 sky130_fd_sc_hd__mux4_2 _25402_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net529),
    .S1(net535),
    .X(_11216_));
 sky130_fd_sc_hd__mux4_2 _25403_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net529),
    .S1(net535),
    .X(_11217_));
 sky130_fd_sc_hd__mux4_2 _25404_ (.A0(_11214_),
    .A1(_11215_),
    .A2(_11216_),
    .A3(_11217_),
    .S0(\count15_1[3] ),
    .S1(net520),
    .X(_11218_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_288 ();
 sky130_fd_sc_hd__mux2i_4 _25406_ (.A0(_11213_),
    .A1(_11218_),
    .S(net518),
    .Y(_11220_));
 sky130_fd_sc_hd__mux4_2 _25407_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net527),
    .S1(net533),
    .X(_11221_));
 sky130_fd_sc_hd__mux4_2 _25408_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net527),
    .S1(net533),
    .X(_11222_));
 sky130_fd_sc_hd__mux4_2 _25409_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net527),
    .S1(net533),
    .X(_11223_));
 sky130_fd_sc_hd__mux4_2 _25410_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net527),
    .S1(net533),
    .X(_11224_));
 sky130_fd_sc_hd__mux4_2 _25411_ (.A0(_11221_),
    .A1(_11222_),
    .A2(_11223_),
    .A3(_11224_),
    .S0(net522),
    .S1(net520),
    .X(_11225_));
 sky130_fd_sc_hd__mux4_2 _25412_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net529),
    .S1(net535),
    .X(_11226_));
 sky130_fd_sc_hd__mux4_2 _25413_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net529),
    .S1(net535),
    .X(_11227_));
 sky130_fd_sc_hd__mux4_2 _25414_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net529),
    .S1(net535),
    .X(_11228_));
 sky130_fd_sc_hd__mux4_2 _25415_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net529),
    .S1(net535),
    .X(_11229_));
 sky130_fd_sc_hd__mux4_2 _25416_ (.A0(_11226_),
    .A1(_11227_),
    .A2(_11228_),
    .A3(_11229_),
    .S0(\count15_1[3] ),
    .S1(net520),
    .X(_11230_));
 sky130_fd_sc_hd__mux2i_4 _25417_ (.A0(_11225_),
    .A1(_11230_),
    .S(net518),
    .Y(_11231_));
 sky130_fd_sc_hd__xnor2_1 _25418_ (.A(_11220_),
    .B(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__xnor2_1 _25419_ (.A(_10917_),
    .B(_11232_),
    .Y(_11619_));
 sky130_fd_sc_hd__mux4_2 _25420_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net446),
    .S1(net452),
    .X(_11233_));
 sky130_fd_sc_hd__mux4_2 _25421_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net446),
    .S1(net452),
    .X(_11234_));
 sky130_fd_sc_hd__mux4_2 _25422_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net446),
    .S1(net552),
    .X(_11235_));
 sky130_fd_sc_hd__mux4_2 _25423_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net446),
    .S1(net552),
    .X(_11236_));
 sky130_fd_sc_hd__mux4_2 _25424_ (.A0(_11233_),
    .A1(_11234_),
    .A2(_11235_),
    .A3(_11236_),
    .S0(net443),
    .S1(net550),
    .X(_11237_));
 sky130_fd_sc_hd__mux4_2 _25425_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net446),
    .S1(net552),
    .X(_11238_));
 sky130_fd_sc_hd__mux4_2 _25426_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net446),
    .S1(net552),
    .X(_11239_));
 sky130_fd_sc_hd__mux4_2 _25427_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net446),
    .S1(net552),
    .X(_11240_));
 sky130_fd_sc_hd__mux4_2 _25428_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net446),
    .S1(net552),
    .X(_11241_));
 sky130_fd_sc_hd__mux4_2 _25429_ (.A0(_11238_),
    .A1(_11239_),
    .A2(_11240_),
    .A3(_11241_),
    .S0(net443),
    .S1(net550),
    .X(_11242_));
 sky130_fd_sc_hd__mux2i_4 _25430_ (.A0(_11237_),
    .A1(_11242_),
    .S(net438),
    .Y(_11243_));
 sky130_fd_sc_hd__mux4_2 _25431_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11244_));
 sky130_fd_sc_hd__mux4_2 _25432_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11245_));
 sky130_fd_sc_hd__mux4_2 _25433_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11246_));
 sky130_fd_sc_hd__mux4_2 _25434_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11247_));
 sky130_fd_sc_hd__mux4_2 _25435_ (.A0(_11244_),
    .A1(_11245_),
    .A2(_11246_),
    .A3(_11247_),
    .S0(net442),
    .S1(net440),
    .X(_11248_));
 sky130_fd_sc_hd__mux4_2 _25436_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11249_));
 sky130_fd_sc_hd__mux4_2 _25437_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11250_));
 sky130_fd_sc_hd__mux4_2 _25438_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11251_));
 sky130_fd_sc_hd__mux4_2 _25439_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net448),
    .S1(net454),
    .X(_11252_));
 sky130_fd_sc_hd__mux4_2 _25440_ (.A0(_11249_),
    .A1(_11250_),
    .A2(_11251_),
    .A3(_11252_),
    .S0(net442),
    .S1(net440),
    .X(_11253_));
 sky130_fd_sc_hd__mux2i_4 _25441_ (.A0(_11248_),
    .A1(_11253_),
    .S(net437),
    .Y(_11254_));
 sky130_fd_sc_hd__xnor2_1 _25442_ (.A(_11243_),
    .B(_11254_),
    .Y(_11255_));
 sky130_fd_sc_hd__xnor2_2 _25443_ (.A(_11158_),
    .B(_11255_),
    .Y(_11624_));
 sky130_fd_sc_hd__mux4_2 _25444_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net530),
    .S1(net560),
    .X(_11256_));
 sky130_fd_sc_hd__mux4_2 _25445_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net530),
    .S1(net560),
    .X(_11257_));
 sky130_fd_sc_hd__mux4_2 _25446_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net530),
    .S1(net560),
    .X(_11258_));
 sky130_fd_sc_hd__mux4_2 _25447_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net530),
    .S1(net560),
    .X(_11259_));
 sky130_fd_sc_hd__mux4_2 _25448_ (.A0(_11256_),
    .A1(_11257_),
    .A2(_11258_),
    .A3(_11259_),
    .S0(net524),
    .S1(net521),
    .X(_11260_));
 sky130_fd_sc_hd__mux4_2 _25449_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net525),
    .S1(net534),
    .X(_11261_));
 sky130_fd_sc_hd__mux4_2 _25450_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net525),
    .S1(net534),
    .X(_11262_));
 sky130_fd_sc_hd__mux4_2 _25451_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net525),
    .S1(net536),
    .X(_11263_));
 sky130_fd_sc_hd__mux4_2 _25452_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net525),
    .S1(net536),
    .X(_11264_));
 sky130_fd_sc_hd__mux4_2 _25453_ (.A0(_11261_),
    .A1(_11262_),
    .A2(_11263_),
    .A3(_11264_),
    .S0(net524),
    .S1(net521),
    .X(_11265_));
 sky130_fd_sc_hd__mux2i_4 _25454_ (.A0(_11260_),
    .A1(_11265_),
    .S(net558),
    .Y(_11266_));
 sky130_fd_sc_hd__mux4_2 _25455_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net531),
    .S1(net535),
    .X(_11267_));
 sky130_fd_sc_hd__mux4_2 _25456_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net531),
    .S1(net535),
    .X(_11268_));
 sky130_fd_sc_hd__mux4_2 _25457_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net531),
    .S1(net535),
    .X(_11269_));
 sky130_fd_sc_hd__mux4_2 _25458_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net531),
    .S1(net535),
    .X(_11270_));
 sky130_fd_sc_hd__mux4_2 _25459_ (.A0(_11267_),
    .A1(_11268_),
    .A2(_11269_),
    .A3(_11270_),
    .S0(net523),
    .S1(net559),
    .X(_11271_));
 sky130_fd_sc_hd__mux4_2 _25460_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net531),
    .S1(net537),
    .X(_11272_));
 sky130_fd_sc_hd__mux4_2 _25461_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net531),
    .S1(net537),
    .X(_11273_));
 sky130_fd_sc_hd__mux4_2 _25462_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net531),
    .S1(net537),
    .X(_11274_));
 sky130_fd_sc_hd__mux4_2 _25463_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net532),
    .S1(net537),
    .X(_11275_));
 sky130_fd_sc_hd__mux4_2 _25464_ (.A0(_11272_),
    .A1(_11273_),
    .A2(_11274_),
    .A3(_11275_),
    .S0(net523),
    .S1(net559),
    .X(_11276_));
 sky130_fd_sc_hd__mux2i_4 _25465_ (.A0(_11271_),
    .A1(_11276_),
    .S(net519),
    .Y(_11277_));
 sky130_fd_sc_hd__xnor2_1 _25466_ (.A(_11266_),
    .B(_11277_),
    .Y(_11278_));
 sky130_fd_sc_hd__xnor2_1 _25467_ (.A(_11045_),
    .B(_11278_),
    .Y(_11627_));
 sky130_fd_sc_hd__mux4_2 _25468_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11279_));
 sky130_fd_sc_hd__mux4_2 _25469_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11280_));
 sky130_fd_sc_hd__mux4_2 _25470_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11281_));
 sky130_fd_sc_hd__mux4_2 _25471_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11282_));
 sky130_fd_sc_hd__mux4_2 _25472_ (.A0(_11279_),
    .A1(_11280_),
    .A2(_11281_),
    .A3(_11282_),
    .S0(net442),
    .S1(net440),
    .X(_11283_));
 sky130_fd_sc_hd__mux4_2 _25473_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11284_));
 sky130_fd_sc_hd__mux4_2 _25474_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11285_));
 sky130_fd_sc_hd__mux4_2 _25475_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11286_));
 sky130_fd_sc_hd__mux4_2 _25476_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net445),
    .S1(net454),
    .X(_11287_));
 sky130_fd_sc_hd__mux4_2 _25477_ (.A0(_11284_),
    .A1(_11285_),
    .A2(_11286_),
    .A3(_11287_),
    .S0(net442),
    .S1(net440),
    .X(_11288_));
 sky130_fd_sc_hd__mux2i_4 _25478_ (.A0(_11283_),
    .A1(_11288_),
    .S(net437),
    .Y(_11289_));
 sky130_fd_sc_hd__mux4_2 _25479_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net446),
    .S1(net552),
    .X(_11290_));
 sky130_fd_sc_hd__mux4_2 _25480_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net446),
    .S1(net552),
    .X(_11291_));
 sky130_fd_sc_hd__mux4_2 _25481_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net446),
    .S1(net552),
    .X(_11292_));
 sky130_fd_sc_hd__mux4_2 _25482_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net446),
    .S1(net552),
    .X(_11293_));
 sky130_fd_sc_hd__mux4_2 _25483_ (.A0(_11290_),
    .A1(_11291_),
    .A2(_11292_),
    .A3(_11293_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11294_));
 sky130_fd_sc_hd__mux4_2 _25484_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net450),
    .S1(net456),
    .X(_11295_));
 sky130_fd_sc_hd__mux4_2 _25485_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_11296_));
 sky130_fd_sc_hd__mux4_2 _25486_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_11297_));
 sky130_fd_sc_hd__mux4_2 _25487_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_11298_));
 sky130_fd_sc_hd__mux4_2 _25488_ (.A0(_11295_),
    .A1(_11296_),
    .A2(_11297_),
    .A3(_11298_),
    .S0(net442),
    .S1(net440),
    .X(_11299_));
 sky130_fd_sc_hd__mux2i_4 _25489_ (.A0(_11294_),
    .A1(_11299_),
    .S(net438),
    .Y(_11300_));
 sky130_fd_sc_hd__xnor2_1 _25490_ (.A(_11289_),
    .B(_11300_),
    .Y(_11301_));
 sky130_fd_sc_hd__xnor2_1 _25491_ (.A(_11207_),
    .B(_11301_),
    .Y(_11632_));
 sky130_fd_sc_hd__mux4_2 _25492_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11302_));
 sky130_fd_sc_hd__mux4_2 _25493_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11303_));
 sky130_fd_sc_hd__mux4_2 _25494_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11304_));
 sky130_fd_sc_hd__mux4_2 _25495_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11305_));
 sky130_fd_sc_hd__mux4_2 _25496_ (.A0(_11302_),
    .A1(_11303_),
    .A2(_11304_),
    .A3(_11305_),
    .S0(net522),
    .S1(net520),
    .X(_11306_));
 sky130_fd_sc_hd__mux4_2 _25497_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11307_));
 sky130_fd_sc_hd__mux4_2 _25498_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11308_));
 sky130_fd_sc_hd__mux4_2 _25499_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11309_));
 sky130_fd_sc_hd__mux4_2 _25500_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net527),
    .S1(net533),
    .X(_11310_));
 sky130_fd_sc_hd__mux4_2 _25501_ (.A0(_11307_),
    .A1(_11308_),
    .A2(_11309_),
    .A3(_11310_),
    .S0(net522),
    .S1(net520),
    .X(_11311_));
 sky130_fd_sc_hd__mux2i_4 _25502_ (.A0(_11306_),
    .A1(_11311_),
    .S(net518),
    .Y(_11312_));
 sky130_fd_sc_hd__mux4_2 _25503_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net527),
    .S1(net533),
    .X(_11313_));
 sky130_fd_sc_hd__mux4_2 _25504_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net527),
    .S1(net533),
    .X(_11314_));
 sky130_fd_sc_hd__mux4_2 _25505_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net527),
    .S1(net533),
    .X(_11315_));
 sky130_fd_sc_hd__mux4_2 _25506_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net527),
    .S1(net533),
    .X(_11316_));
 sky130_fd_sc_hd__mux4_2 _25507_ (.A0(_11313_),
    .A1(_11314_),
    .A2(_11315_),
    .A3(_11316_),
    .S0(net522),
    .S1(net520),
    .X(_11317_));
 sky130_fd_sc_hd__mux4_2 _25508_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net528),
    .S1(net533),
    .X(_11318_));
 sky130_fd_sc_hd__mux4_2 _25509_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net528),
    .S1(net533),
    .X(_11319_));
 sky130_fd_sc_hd__mux4_2 _25510_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net528),
    .S1(net533),
    .X(_11320_));
 sky130_fd_sc_hd__mux4_2 _25511_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net528),
    .S1(net533),
    .X(_11321_));
 sky130_fd_sc_hd__mux4_2 _25512_ (.A0(_11318_),
    .A1(_11319_),
    .A2(_11320_),
    .A3(_11321_),
    .S0(net522),
    .S1(net520),
    .X(_11322_));
 sky130_fd_sc_hd__mux2i_4 _25513_ (.A0(_11317_),
    .A1(_11322_),
    .S(net518),
    .Y(_11323_));
 sky130_fd_sc_hd__xnor2_1 _25514_ (.A(_11312_),
    .B(_11323_),
    .Y(_11324_));
 sky130_fd_sc_hd__xnor2_1 _25515_ (.A(_11129_),
    .B(_11324_),
    .Y(_11635_));
 sky130_fd_sc_hd__mux4_2 _25516_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net445),
    .S1(net451),
    .X(_11325_));
 sky130_fd_sc_hd__mux4_2 _25517_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net445),
    .S1(net451),
    .X(_11326_));
 sky130_fd_sc_hd__mux4_2 _25518_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net445),
    .S1(net451),
    .X(_11327_));
 sky130_fd_sc_hd__mux4_2 _25519_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net445),
    .S1(net451),
    .X(_11328_));
 sky130_fd_sc_hd__mux4_2 _25520_ (.A0(_11325_),
    .A1(_11326_),
    .A2(_11327_),
    .A3(_11328_),
    .S0(net442),
    .S1(net440),
    .X(_11329_));
 sky130_fd_sc_hd__mux4_2 _25521_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net445),
    .S1(net456),
    .X(_11330_));
 sky130_fd_sc_hd__mux4_2 _25522_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net445),
    .S1(net456),
    .X(_11331_));
 sky130_fd_sc_hd__mux4_2 _25523_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net445),
    .S1(net456),
    .X(_11332_));
 sky130_fd_sc_hd__mux4_2 _25524_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net445),
    .S1(net456),
    .X(_11333_));
 sky130_fd_sc_hd__mux4_2 _25525_ (.A0(_11330_),
    .A1(_11331_),
    .A2(_11332_),
    .A3(_11333_),
    .S0(net442),
    .S1(net440),
    .X(_11334_));
 sky130_fd_sc_hd__mux2i_4 _25526_ (.A0(_11329_),
    .A1(_11334_),
    .S(net437),
    .Y(_11335_));
 sky130_fd_sc_hd__mux4_2 _25527_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11336_));
 sky130_fd_sc_hd__mux4_2 _25528_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11337_));
 sky130_fd_sc_hd__mux4_2 _25529_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11338_));
 sky130_fd_sc_hd__mux4_2 _25530_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11339_));
 sky130_fd_sc_hd__mux4_2 _25531_ (.A0(_11336_),
    .A1(_11337_),
    .A2(_11338_),
    .A3(_11339_),
    .S0(net442),
    .S1(net440),
    .X(_11340_));
 sky130_fd_sc_hd__mux4_2 _25532_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11341_));
 sky130_fd_sc_hd__mux4_2 _25533_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11342_));
 sky130_fd_sc_hd__mux4_2 _25534_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11343_));
 sky130_fd_sc_hd__mux4_2 _25535_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net448),
    .S1(net454),
    .X(_11344_));
 sky130_fd_sc_hd__mux4_2 _25536_ (.A0(_11341_),
    .A1(_11342_),
    .A2(_11343_),
    .A3(_11344_),
    .S0(net442),
    .S1(net440),
    .X(_11345_));
 sky130_fd_sc_hd__mux2i_4 _25537_ (.A0(_11340_),
    .A1(_11345_),
    .S(net437),
    .Y(_11346_));
 sky130_fd_sc_hd__xnor2_1 _25538_ (.A(_11335_),
    .B(_11346_),
    .Y(_11347_));
 sky130_fd_sc_hd__xnor2_1 _25539_ (.A(_11254_),
    .B(_11347_),
    .Y(_11640_));
 sky130_fd_sc_hd__mux4_2 _25540_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net530),
    .S1(net560),
    .X(_11348_));
 sky130_fd_sc_hd__mux4_2 _25541_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net530),
    .S1(net560),
    .X(_11349_));
 sky130_fd_sc_hd__mux4_2 _25542_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net530),
    .S1(net560),
    .X(_11350_));
 sky130_fd_sc_hd__mux4_2 _25543_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net530),
    .S1(net560),
    .X(_11351_));
 sky130_fd_sc_hd__mux4_2 _25544_ (.A0(_11348_),
    .A1(_11349_),
    .A2(_11350_),
    .A3(_11351_),
    .S0(net524),
    .S1(net521),
    .X(_11352_));
 sky130_fd_sc_hd__mux4_2 _25545_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net529),
    .S1(net535),
    .X(_11353_));
 sky130_fd_sc_hd__mux4_2 _25546_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net529),
    .S1(net535),
    .X(_11354_));
 sky130_fd_sc_hd__mux4_2 _25547_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net529),
    .S1(net535),
    .X(_11355_));
 sky130_fd_sc_hd__mux4_2 _25548_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net529),
    .S1(net535),
    .X(_11356_));
 sky130_fd_sc_hd__mux4_2 _25549_ (.A0(_11353_),
    .A1(_11354_),
    .A2(_11355_),
    .A3(_11356_),
    .S0(\count15_1[3] ),
    .S1(net520),
    .X(_11357_));
 sky130_fd_sc_hd__mux2i_4 _25550_ (.A0(_11352_),
    .A1(_11357_),
    .S(net518),
    .Y(_11358_));
 sky130_fd_sc_hd__mux4_2 _25551_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net530),
    .S1(net560),
    .X(_11359_));
 sky130_fd_sc_hd__mux4_2 _25552_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(\count15_1[2] ),
    .S1(net560),
    .X(_11360_));
 sky130_fd_sc_hd__mux4_2 _25553_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net530),
    .S1(net560),
    .X(_11361_));
 sky130_fd_sc_hd__mux4_2 _25554_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net530),
    .S1(net560),
    .X(_11362_));
 sky130_fd_sc_hd__mux4_2 _25555_ (.A0(_11359_),
    .A1(_11360_),
    .A2(_11361_),
    .A3(_11362_),
    .S0(net524),
    .S1(net521),
    .X(_11363_));
 sky130_fd_sc_hd__mux4_2 _25556_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net525),
    .S1(net535),
    .X(_11364_));
 sky130_fd_sc_hd__mux4_2 _25557_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net525),
    .S1(net536),
    .X(_11365_));
 sky130_fd_sc_hd__mux4_2 _25558_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net530),
    .S1(net536),
    .X(_11366_));
 sky130_fd_sc_hd__mux4_2 _25559_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net530),
    .S1(net536),
    .X(_11367_));
 sky130_fd_sc_hd__mux4_2 _25560_ (.A0(_11364_),
    .A1(_11365_),
    .A2(_11366_),
    .A3(_11367_),
    .S0(net524),
    .S1(net521),
    .X(_11368_));
 sky130_fd_sc_hd__mux2i_4 _25561_ (.A0(_11363_),
    .A1(_11368_),
    .S(net558),
    .Y(_11369_));
 sky130_fd_sc_hd__xnor2_1 _25562_ (.A(_11358_),
    .B(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__xnor2_1 _25563_ (.A(_11184_),
    .B(_11370_),
    .Y(_11643_));
 sky130_fd_sc_hd__mux4_2 _25564_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net444),
    .S1(net451),
    .X(_11371_));
 sky130_fd_sc_hd__mux4_2 _25565_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net444),
    .S1(net451),
    .X(_11372_));
 sky130_fd_sc_hd__mux4_2 _25566_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net444),
    .S1(net451),
    .X(_11373_));
 sky130_fd_sc_hd__mux4_2 _25567_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net444),
    .S1(net451),
    .X(_11374_));
 sky130_fd_sc_hd__mux4_2 _25568_ (.A0(_11371_),
    .A1(_11372_),
    .A2(_11373_),
    .A3(_11374_),
    .S0(net443),
    .S1(net550),
    .X(_11375_));
 sky130_fd_sc_hd__mux4_2 _25569_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net444),
    .S1(net451),
    .X(_11376_));
 sky130_fd_sc_hd__mux4_2 _25570_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net444),
    .S1(net451),
    .X(_11377_));
 sky130_fd_sc_hd__mux4_2 _25571_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net444),
    .S1(net451),
    .X(_11378_));
 sky130_fd_sc_hd__mux4_2 _25572_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net445),
    .S1(net451),
    .X(_11379_));
 sky130_fd_sc_hd__mux4_2 _25573_ (.A0(_11376_),
    .A1(_11377_),
    .A2(_11378_),
    .A3(_11379_),
    .S0(net443),
    .S1(net550),
    .X(_11380_));
 sky130_fd_sc_hd__mux2i_4 _25574_ (.A0(_11375_),
    .A1(_11380_),
    .S(net438),
    .Y(_11381_));
 sky130_fd_sc_hd__xnor2_1 _25575_ (.A(_11289_),
    .B(_11381_),
    .Y(_11382_));
 sky130_fd_sc_hd__xnor2_1 _25576_ (.A(_11006_),
    .B(_11382_),
    .Y(_11648_));
 sky130_fd_sc_hd__mux4_2 _25577_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net526),
    .S1(net534),
    .X(_11383_));
 sky130_fd_sc_hd__mux4_2 _25578_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net526),
    .S1(net534),
    .X(_11384_));
 sky130_fd_sc_hd__mux4_2 _25579_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net526),
    .S1(net534),
    .X(_11385_));
 sky130_fd_sc_hd__mux4_2 _25580_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net526),
    .S1(net534),
    .X(_11386_));
 sky130_fd_sc_hd__mux4_2 _25581_ (.A0(_11383_),
    .A1(_11384_),
    .A2(_11385_),
    .A3(_11386_),
    .S0(net522),
    .S1(net520),
    .X(_11387_));
 sky130_fd_sc_hd__mux4_2 _25582_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net528),
    .S1(net535),
    .X(_11388_));
 sky130_fd_sc_hd__mux4_2 _25583_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net528),
    .S1(net535),
    .X(_11389_));
 sky130_fd_sc_hd__mux4_2 _25584_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net528),
    .S1(net535),
    .X(_11390_));
 sky130_fd_sc_hd__mux4_2 _25585_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net529),
    .S1(net535),
    .X(_11391_));
 sky130_fd_sc_hd__mux4_2 _25586_ (.A0(_11388_),
    .A1(_11389_),
    .A2(_11390_),
    .A3(_11391_),
    .S0(net522),
    .S1(net520),
    .X(_11392_));
 sky130_fd_sc_hd__mux2i_4 _25587_ (.A0(_11387_),
    .A1(_11392_),
    .S(net518),
    .Y(_11393_));
 sky130_fd_sc_hd__mux4_2 _25588_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net526),
    .S1(net534),
    .X(_11394_));
 sky130_fd_sc_hd__mux4_2 _25589_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net526),
    .S1(net534),
    .X(_11395_));
 sky130_fd_sc_hd__mux4_2 _25590_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net526),
    .S1(net534),
    .X(_11396_));
 sky130_fd_sc_hd__mux4_2 _25591_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net526),
    .S1(net534),
    .X(_11397_));
 sky130_fd_sc_hd__mux4_2 _25592_ (.A0(_11394_),
    .A1(_11395_),
    .A2(_11396_),
    .A3(_11397_),
    .S0(net522),
    .S1(net520),
    .X(_11398_));
 sky130_fd_sc_hd__mux4_2 _25593_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net529),
    .S1(net535),
    .X(_11399_));
 sky130_fd_sc_hd__mux4_2 _25594_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net529),
    .S1(net535),
    .X(_11400_));
 sky130_fd_sc_hd__mux4_2 _25595_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net529),
    .S1(net535),
    .X(_11401_));
 sky130_fd_sc_hd__mux4_2 _25596_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net529),
    .S1(net535),
    .X(_11402_));
 sky130_fd_sc_hd__mux4_2 _25597_ (.A0(_11399_),
    .A1(_11400_),
    .A2(_11401_),
    .A3(_11402_),
    .S0(net522),
    .S1(net520),
    .X(_11403_));
 sky130_fd_sc_hd__mux2i_4 _25598_ (.A0(_11398_),
    .A1(_11403_),
    .S(net518),
    .Y(_11404_));
 sky130_fd_sc_hd__xnor2_1 _25599_ (.A(_11393_),
    .B(_11404_),
    .Y(_11405_));
 sky130_fd_sc_hd__xnor2_1 _25600_ (.A(_11231_),
    .B(_11405_),
    .Y(_11651_));
 sky130_fd_sc_hd__mux4_2 _25601_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net444),
    .S1(net451),
    .X(_11406_));
 sky130_fd_sc_hd__mux4_2 _25602_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net444),
    .S1(net451),
    .X(_11407_));
 sky130_fd_sc_hd__mux4_2 _25603_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net444),
    .S1(net451),
    .X(_11408_));
 sky130_fd_sc_hd__mux4_2 _25604_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net444),
    .S1(net451),
    .X(_11409_));
 sky130_fd_sc_hd__mux4_2 _25605_ (.A0(_11406_),
    .A1(_11407_),
    .A2(_11408_),
    .A3(_11409_),
    .S0(net442),
    .S1(net440),
    .X(_11410_));
 sky130_fd_sc_hd__mux4_2 _25606_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net450),
    .S1(net455),
    .X(_11411_));
 sky130_fd_sc_hd__mux4_2 _25607_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net449),
    .S1(net455),
    .X(_11412_));
 sky130_fd_sc_hd__mux4_2 _25608_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net449),
    .S1(net455),
    .X(_11413_));
 sky130_fd_sc_hd__mux4_2 _25609_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net450),
    .S1(net455),
    .X(_11414_));
 sky130_fd_sc_hd__mux4_2 _25610_ (.A0(_11411_),
    .A1(_11412_),
    .A2(_11413_),
    .A3(_11414_),
    .S0(net441),
    .S1(net439),
    .X(_11415_));
 sky130_fd_sc_hd__mux2i_4 _25611_ (.A0(_11410_),
    .A1(_11415_),
    .S(net437),
    .Y(_11416_));
 sky130_fd_sc_hd__xnor2_1 _25612_ (.A(_11346_),
    .B(_11416_),
    .Y(_11417_));
 sky130_fd_sc_hd__xnor2_1 _25613_ (.A(_11090_),
    .B(_11417_),
    .Y(_11656_));
 sky130_fd_sc_hd__mux4_2 _25614_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net528),
    .S1(net536),
    .X(_11418_));
 sky130_fd_sc_hd__mux4_2 _25615_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net528),
    .S1(net536),
    .X(_11419_));
 sky130_fd_sc_hd__mux4_2 _25616_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net528),
    .S1(net536),
    .X(_11420_));
 sky130_fd_sc_hd__mux4_2 _25617_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net528),
    .S1(net536),
    .X(_11421_));
 sky130_fd_sc_hd__mux4_2 _25618_ (.A0(_11418_),
    .A1(_11419_),
    .A2(_11420_),
    .A3(_11421_),
    .S0(net522),
    .S1(net521),
    .X(_11422_));
 sky130_fd_sc_hd__mux4_2 _25619_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net528),
    .S1(net534),
    .X(_11423_));
 sky130_fd_sc_hd__mux4_2 _25620_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net528),
    .S1(net534),
    .X(_11424_));
 sky130_fd_sc_hd__mux4_2 _25621_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net528),
    .S1(net534),
    .X(_11425_));
 sky130_fd_sc_hd__mux4_2 _25622_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net528),
    .S1(net534),
    .X(_11426_));
 sky130_fd_sc_hd__mux4_2 _25623_ (.A0(_11423_),
    .A1(_11424_),
    .A2(_11425_),
    .A3(_11426_),
    .S0(net522),
    .S1(net520),
    .X(_11427_));
 sky130_fd_sc_hd__mux2i_4 _25624_ (.A0(_11422_),
    .A1(_11427_),
    .S(net518),
    .Y(_11428_));
 sky130_fd_sc_hd__mux4_2 _25625_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net530),
    .S1(net560),
    .X(_11429_));
 sky130_fd_sc_hd__mux4_2 _25626_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net530),
    .S1(net560),
    .X(_11430_));
 sky130_fd_sc_hd__mux4_2 _25627_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net530),
    .S1(net560),
    .X(_11431_));
 sky130_fd_sc_hd__mux4_2 _25628_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net530),
    .S1(net560),
    .X(_11432_));
 sky130_fd_sc_hd__mux4_2 _25629_ (.A0(_11429_),
    .A1(_11430_),
    .A2(_11431_),
    .A3(_11432_),
    .S0(net524),
    .S1(net521),
    .X(_11433_));
 sky130_fd_sc_hd__mux4_2 _25630_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net525),
    .S1(net536),
    .X(_11434_));
 sky130_fd_sc_hd__mux4_2 _25631_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net525),
    .S1(net536),
    .X(_11435_));
 sky130_fd_sc_hd__mux4_2 _25632_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net525),
    .S1(net536),
    .X(_11436_));
 sky130_fd_sc_hd__mux4_2 _25633_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net525),
    .S1(net536),
    .X(_11437_));
 sky130_fd_sc_hd__mux4_2 _25634_ (.A0(_11434_),
    .A1(_11435_),
    .A2(_11436_),
    .A3(_11437_),
    .S0(net524),
    .S1(net521),
    .X(_11438_));
 sky130_fd_sc_hd__mux2i_4 _25635_ (.A0(_11433_),
    .A1(_11438_),
    .S(net558),
    .Y(_11439_));
 sky130_fd_sc_hd__xnor2_1 _25636_ (.A(_11428_),
    .B(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__xnor2_1 _25637_ (.A(_11277_),
    .B(_11440_),
    .Y(_11659_));
 sky130_fd_sc_hd__mux4_2 _25638_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net551),
    .S1(net452),
    .X(_11441_));
 sky130_fd_sc_hd__mux4_2 _25639_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net551),
    .S1(net452),
    .X(_11442_));
 sky130_fd_sc_hd__mux4_2 _25640_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net551),
    .S1(net452),
    .X(_11443_));
 sky130_fd_sc_hd__mux4_2 _25641_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net551),
    .S1(net452),
    .X(_11444_));
 sky130_fd_sc_hd__mux4_2 _25642_ (.A0(_11441_),
    .A1(_11442_),
    .A2(_11443_),
    .A3(_11444_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11445_));
 sky130_fd_sc_hd__mux4_2 _25643_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net446),
    .S1(net452),
    .X(_11446_));
 sky130_fd_sc_hd__mux4_2 _25644_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net446),
    .S1(net452),
    .X(_11447_));
 sky130_fd_sc_hd__mux4_2 _25645_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net446),
    .S1(net452),
    .X(_11448_));
 sky130_fd_sc_hd__mux4_2 _25646_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net446),
    .S1(net452),
    .X(_11449_));
 sky130_fd_sc_hd__mux4_2 _25647_ (.A0(_11446_),
    .A1(_11447_),
    .A2(_11448_),
    .A3(_11449_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11450_));
 sky130_fd_sc_hd__mux2i_4 _25648_ (.A0(_11445_),
    .A1(_11450_),
    .S(\count2_1[5] ),
    .Y(_11451_));
 sky130_fd_sc_hd__xnor2_1 _25649_ (.A(_11381_),
    .B(_11451_),
    .Y(_11452_));
 sky130_fd_sc_hd__xnor2_1 _25650_ (.A(_10995_),
    .B(_11452_),
    .Y(_11664_));
 sky130_fd_sc_hd__mux4_2 _25651_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net530),
    .S1(net560),
    .X(_11453_));
 sky130_fd_sc_hd__mux4_2 _25652_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net530),
    .S1(net560),
    .X(_11454_));
 sky130_fd_sc_hd__mux4_2 _25653_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net530),
    .S1(net560),
    .X(_11455_));
 sky130_fd_sc_hd__mux4_2 _25654_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net530),
    .S1(net560),
    .X(_11456_));
 sky130_fd_sc_hd__mux4_2 _25655_ (.A0(_11453_),
    .A1(_11454_),
    .A2(_11455_),
    .A3(_11456_),
    .S0(net524),
    .S1(net521),
    .X(_11457_));
 sky130_fd_sc_hd__mux4_2 _25656_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net525),
    .S1(net536),
    .X(_11458_));
 sky130_fd_sc_hd__mux4_2 _25657_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net525),
    .S1(net536),
    .X(_11459_));
 sky130_fd_sc_hd__mux4_2 _25658_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net525),
    .S1(net536),
    .X(_11460_));
 sky130_fd_sc_hd__mux4_2 _25659_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net525),
    .S1(net536),
    .X(_11461_));
 sky130_fd_sc_hd__mux4_2 _25660_ (.A0(_11458_),
    .A1(_11459_),
    .A2(_11460_),
    .A3(_11461_),
    .S0(net524),
    .S1(net521),
    .X(_11462_));
 sky130_fd_sc_hd__mux2i_4 _25661_ (.A0(_11457_),
    .A1(_11462_),
    .S(net558),
    .Y(_11463_));
 sky130_fd_sc_hd__xnor2_1 _25662_ (.A(_11312_),
    .B(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__xnor2_1 _25663_ (.A(_10865_),
    .B(_11464_),
    .Y(_11667_));
 sky130_fd_sc_hd__mux4_2 _25664_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net551),
    .S1(net452),
    .X(_11465_));
 sky130_fd_sc_hd__mux4_2 _25665_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net551),
    .S1(net452),
    .X(_11466_));
 sky130_fd_sc_hd__mux4_2 _25666_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net551),
    .S1(net452),
    .X(_11467_));
 sky130_fd_sc_hd__mux4_2 _25667_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net551),
    .S1(net452),
    .X(_11468_));
 sky130_fd_sc_hd__mux4_2 _25668_ (.A0(_11465_),
    .A1(_11466_),
    .A2(_11467_),
    .A3(_11468_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11469_));
 sky130_fd_sc_hd__mux4_2 _25669_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net446),
    .S1(net452),
    .X(_11470_));
 sky130_fd_sc_hd__mux4_2 _25670_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net446),
    .S1(net452),
    .X(_11471_));
 sky130_fd_sc_hd__mux4_2 _25671_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net446),
    .S1(net452),
    .X(_11472_));
 sky130_fd_sc_hd__mux4_2 _25672_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net446),
    .S1(net452),
    .X(_11473_));
 sky130_fd_sc_hd__mux4_2 _25673_ (.A0(_11470_),
    .A1(_11471_),
    .A2(_11472_),
    .A3(_11473_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11474_));
 sky130_fd_sc_hd__mux2i_4 _25674_ (.A0(_11469_),
    .A1(_11474_),
    .S(\count2_1[5] ),
    .Y(_11475_));
 sky130_fd_sc_hd__xnor2_1 _25675_ (.A(_11416_),
    .B(_11475_),
    .Y(_11476_));
 sky130_fd_sc_hd__xnor2_1 _25676_ (.A(_11071_),
    .B(_11476_),
    .Y(_11672_));
 sky130_fd_sc_hd__mux4_2 _25677_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(\count15_1[2] ),
    .S1(net536),
    .X(_11477_));
 sky130_fd_sc_hd__mux4_2 _25678_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(\count15_1[2] ),
    .S1(net536),
    .X(_11478_));
 sky130_fd_sc_hd__mux4_2 _25679_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(\count15_1[2] ),
    .S1(net537),
    .X(_11479_));
 sky130_fd_sc_hd__mux4_2 _25680_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(\count15_1[2] ),
    .S1(net537),
    .X(_11480_));
 sky130_fd_sc_hd__mux4_2 _25681_ (.A0(_11477_),
    .A1(_11478_),
    .A2(_11479_),
    .A3(_11480_),
    .S0(net524),
    .S1(net521),
    .X(_11481_));
 sky130_fd_sc_hd__mux4_2 _25682_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net532),
    .S1(net537),
    .X(_11482_));
 sky130_fd_sc_hd__mux4_2 _25683_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net532),
    .S1(net537),
    .X(_11483_));
 sky130_fd_sc_hd__mux4_2 _25684_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net532),
    .S1(net537),
    .X(_11484_));
 sky130_fd_sc_hd__mux4_2 _25685_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net532),
    .S1(net537),
    .X(_11485_));
 sky130_fd_sc_hd__mux4_2 _25686_ (.A0(_11482_),
    .A1(_11483_),
    .A2(_11484_),
    .A3(_11485_),
    .S0(net523),
    .S1(net559),
    .X(_11486_));
 sky130_fd_sc_hd__mux2i_4 _25687_ (.A0(_11481_),
    .A1(_11486_),
    .S(net519),
    .Y(_11487_));
 sky130_fd_sc_hd__xnor2_1 _25688_ (.A(_11369_),
    .B(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__xnor2_1 _25689_ (.A(_10928_),
    .B(_11488_),
    .Y(_11675_));
 sky130_fd_sc_hd__mux4_2 _25690_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net445),
    .S1(net456),
    .X(_11489_));
 sky130_fd_sc_hd__mux4_2 _25691_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net445),
    .S1(net456),
    .X(_11490_));
 sky130_fd_sc_hd__mux4_2 _25692_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net445),
    .S1(net456),
    .X(_11491_));
 sky130_fd_sc_hd__mux4_2 _25693_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net445),
    .S1(net456),
    .X(_11492_));
 sky130_fd_sc_hd__mux4_2 _25694_ (.A0(_11489_),
    .A1(_11490_),
    .A2(_11491_),
    .A3(_11492_),
    .S0(net442),
    .S1(net440),
    .X(_11493_));
 sky130_fd_sc_hd__mux4_2 _25695_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net450),
    .S1(net455),
    .X(_11494_));
 sky130_fd_sc_hd__mux4_2 _25696_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net450),
    .S1(net455),
    .X(_11495_));
 sky130_fd_sc_hd__mux4_2 _25697_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net450),
    .S1(net455),
    .X(_11496_));
 sky130_fd_sc_hd__mux4_2 _25698_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net450),
    .S1(net455),
    .X(_11497_));
 sky130_fd_sc_hd__mux4_2 _25699_ (.A0(_11494_),
    .A1(_11495_),
    .A2(_11496_),
    .A3(_11497_),
    .S0(net441),
    .S1(net439),
    .X(_11498_));
 sky130_fd_sc_hd__mux2i_4 _25700_ (.A0(_11493_),
    .A1(_11498_),
    .S(net438),
    .Y(_11499_));
 sky130_fd_sc_hd__xnor2_1 _25701_ (.A(_11451_),
    .B(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__xnor2_1 _25702_ (.A(_11158_),
    .B(_11500_),
    .Y(_11680_));
 sky130_fd_sc_hd__mux4_2 _25703_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11501_));
 sky130_fd_sc_hd__mux4_2 _25704_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11502_));
 sky130_fd_sc_hd__mux4_2 _25705_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11503_));
 sky130_fd_sc_hd__mux4_2 _25706_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11504_));
 sky130_fd_sc_hd__mux4_2 _25707_ (.A0(_11501_),
    .A1(_11502_),
    .A2(_11503_),
    .A3(_11504_),
    .S0(net522),
    .S1(net521),
    .X(_11505_));
 sky130_fd_sc_hd__mux4_2 _25708_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11506_));
 sky130_fd_sc_hd__mux4_2 _25709_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11507_));
 sky130_fd_sc_hd__mux4_2 _25710_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11508_));
 sky130_fd_sc_hd__mux4_2 _25711_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net528),
    .S1(net536),
    .X(_11509_));
 sky130_fd_sc_hd__mux4_2 _25712_ (.A0(_11506_),
    .A1(_11507_),
    .A2(_11508_),
    .A3(_11509_),
    .S0(net522),
    .S1(net521),
    .X(_11510_));
 sky130_fd_sc_hd__mux2i_4 _25713_ (.A0(_11505_),
    .A1(_11510_),
    .S(net558),
    .Y(_11511_));
 sky130_fd_sc_hd__xnor2_1 _25714_ (.A(_11404_),
    .B(_11511_),
    .Y(_11512_));
 sky130_fd_sc_hd__xnor2_1 _25715_ (.A(_11022_),
    .B(_11512_),
    .Y(_11683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_286 ();
 sky130_fd_sc_hd__mux4_2 _25718_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_284 ();
 sky130_fd_sc_hd__mux4_2 _25721_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11518_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_282 ();
 sky130_fd_sc_hd__mux4_2 _25724_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_280 ();
 sky130_fd_sc_hd__mux4_2 _25727_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11524_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_278 ();
 sky130_fd_sc_hd__mux4_2 _25730_ (.A0(_11515_),
    .A1(_11518_),
    .A2(_11521_),
    .A3(_11524_),
    .S0(net441),
    .S1(net439),
    .X(_11527_));
 sky130_fd_sc_hd__mux4_2 _25731_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11528_));
 sky130_fd_sc_hd__mux4_2 _25732_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11529_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_276 ();
 sky130_fd_sc_hd__mux4_2 _25735_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_274 ();
 sky130_fd_sc_hd__mux4_2 _25738_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net447),
    .S1(net453),
    .X(_11535_));
 sky130_fd_sc_hd__mux4_2 _25739_ (.A0(_11528_),
    .A1(_11529_),
    .A2(_11532_),
    .A3(_11535_),
    .S0(net441),
    .S1(net439),
    .X(_11536_));
 sky130_fd_sc_hd__mux2i_4 _25740_ (.A0(_11527_),
    .A1(_11536_),
    .S(net437),
    .Y(_11537_));
 sky130_fd_sc_hd__xnor2_1 _25741_ (.A(_11475_),
    .B(_11537_),
    .Y(_11538_));
 sky130_fd_sc_hd__xnor2_1 _25742_ (.A(_11207_),
    .B(_11538_),
    .Y(_11688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_272 ();
 sky130_fd_sc_hd__mux4_2 _25745_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11541_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_270 ();
 sky130_fd_sc_hd__mux4_2 _25748_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11544_));
 sky130_fd_sc_hd__mux4_2 _25749_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11545_));
 sky130_fd_sc_hd__mux4_2 _25750_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11546_));
 sky130_fd_sc_hd__mux4_2 _25751_ (.A0(_11541_),
    .A1(_11544_),
    .A2(_11545_),
    .A3(_11546_),
    .S0(net522),
    .S1(net520),
    .X(_11547_));
 sky130_fd_sc_hd__mux4_2 _25752_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11548_));
 sky130_fd_sc_hd__mux4_2 _25753_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11549_));
 sky130_fd_sc_hd__mux4_2 _25754_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11550_));
 sky130_fd_sc_hd__mux4_2 _25755_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net526),
    .S1(net534),
    .X(_11551_));
 sky130_fd_sc_hd__mux4_2 _25756_ (.A0(_11548_),
    .A1(_11549_),
    .A2(_11550_),
    .A3(_11551_),
    .S0(net522),
    .S1(net520),
    .X(_11552_));
 sky130_fd_sc_hd__mux2i_4 _25757_ (.A0(_11547_),
    .A1(_11552_),
    .S(net518),
    .Y(_11553_));
 sky130_fd_sc_hd__xnor2_1 _25758_ (.A(_11428_),
    .B(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__xnor2_1 _25759_ (.A(_11117_),
    .B(_11554_),
    .Y(_11691_));
 sky130_fd_sc_hd__mux4_2 _25760_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net448),
    .S1(net454),
    .X(_11555_));
 sky130_fd_sc_hd__mux4_2 _25761_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net444),
    .S1(net454),
    .X(_11556_));
 sky130_fd_sc_hd__mux4_2 _25762_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net448),
    .S1(net454),
    .X(_11557_));
 sky130_fd_sc_hd__mux4_2 _25763_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net448),
    .S1(net454),
    .X(_11558_));
 sky130_fd_sc_hd__mux4_2 _25764_ (.A0(_11555_),
    .A1(_11556_),
    .A2(_11557_),
    .A3(_11558_),
    .S0(net442),
    .S1(net440),
    .X(_11559_));
 sky130_fd_sc_hd__mux4_2 _25765_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net449),
    .S1(net455),
    .X(_11560_));
 sky130_fd_sc_hd__mux4_2 _25766_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net449),
    .S1(net455),
    .X(_11561_));
 sky130_fd_sc_hd__mux4_2 _25767_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net449),
    .S1(net455),
    .X(_11562_));
 sky130_fd_sc_hd__mux4_2 _25768_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net449),
    .S1(net455),
    .X(_11563_));
 sky130_fd_sc_hd__mux4_2 _25769_ (.A0(_11560_),
    .A1(_11561_),
    .A2(_11562_),
    .A3(_11563_),
    .S0(net441),
    .S1(net439),
    .X(_11564_));
 sky130_fd_sc_hd__mux2i_4 _25770_ (.A0(_11559_),
    .A1(_11564_),
    .S(net437),
    .Y(_11565_));
 sky130_fd_sc_hd__xnor2_1 _25771_ (.A(_11499_),
    .B(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__xnor2_1 _25772_ (.A(_11254_),
    .B(_11566_),
    .Y(_11696_));
 sky130_fd_sc_hd__mux4_2 _25773_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net526),
    .S1(net534),
    .X(_11567_));
 sky130_fd_sc_hd__mux4_2 _25774_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net526),
    .S1(net534),
    .X(_11568_));
 sky130_fd_sc_hd__mux4_2 _25775_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net526),
    .S1(net534),
    .X(_11569_));
 sky130_fd_sc_hd__mux4_2 _25776_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net526),
    .S1(net534),
    .X(_11570_));
 sky130_fd_sc_hd__mux4_2 _25777_ (.A0(_11567_),
    .A1(_11568_),
    .A2(_11569_),
    .A3(_11570_),
    .S0(net522),
    .S1(net520),
    .X(_11571_));
 sky130_fd_sc_hd__mux4_2 _25778_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net526),
    .S1(net534),
    .X(_11572_));
 sky130_fd_sc_hd__mux4_2 _25779_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net526),
    .S1(net534),
    .X(_11573_));
 sky130_fd_sc_hd__mux4_2 _25780_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net526),
    .S1(net534),
    .X(_11574_));
 sky130_fd_sc_hd__mux4_2 _25781_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net526),
    .S1(net534),
    .X(_02570_));
 sky130_fd_sc_hd__mux4_2 _25782_ (.A0(_11572_),
    .A1(_11573_),
    .A2(_11574_),
    .A3(_02570_),
    .S0(net522),
    .S1(net520),
    .X(_02571_));
 sky130_fd_sc_hd__mux2i_4 _25783_ (.A0(_11571_),
    .A1(_02571_),
    .S(net558),
    .Y(_02572_));
 sky130_fd_sc_hd__xnor2_1 _25784_ (.A(_11172_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_1 _25785_ (.A(_10865_),
    .B(_02573_),
    .Y(_11699_));
 sky130_fd_sc_hd__mux4_2 _25786_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net446),
    .S1(net452),
    .X(_02574_));
 sky130_fd_sc_hd__mux4_2 _25787_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net446),
    .S1(net452),
    .X(_02575_));
 sky130_fd_sc_hd__mux4_2 _25788_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net446),
    .S1(net452),
    .X(_02576_));
 sky130_fd_sc_hd__mux4_2 _25789_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net446),
    .S1(net452),
    .X(_02577_));
 sky130_fd_sc_hd__mux4_2 _25790_ (.A0(_02574_),
    .A1(_02575_),
    .A2(_02576_),
    .A3(_02577_),
    .S0(net443),
    .S1(net550),
    .X(_02578_));
 sky130_fd_sc_hd__mux4_2 _25791_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net446),
    .S1(net552),
    .X(_02579_));
 sky130_fd_sc_hd__mux4_2 _25792_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net446),
    .S1(net552),
    .X(_02580_));
 sky130_fd_sc_hd__mux4_2 _25793_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net446),
    .S1(net552),
    .X(_02581_));
 sky130_fd_sc_hd__mux4_2 _25794_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net446),
    .S1(net552),
    .X(_02582_));
 sky130_fd_sc_hd__mux4_2 _25795_ (.A0(_02579_),
    .A1(_02580_),
    .A2(_02581_),
    .A3(_02582_),
    .S0(net443),
    .S1(net550),
    .X(_02583_));
 sky130_fd_sc_hd__mux2i_4 _25796_ (.A0(_02578_),
    .A1(_02583_),
    .S(net438),
    .Y(_02584_));
 sky130_fd_sc_hd__xnor2_1 _25797_ (.A(_11537_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__xnor2_1 _25798_ (.A(_11289_),
    .B(_02585_),
    .Y(_11704_));
 sky130_fd_sc_hd__mux4_2 _25799_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net526),
    .S1(net534),
    .X(_02586_));
 sky130_fd_sc_hd__mux4_2 _25800_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net526),
    .S1(net534),
    .X(_02587_));
 sky130_fd_sc_hd__mux4_2 _25801_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net526),
    .S1(net534),
    .X(_02588_));
 sky130_fd_sc_hd__mux4_2 _25802_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net526),
    .S1(net534),
    .X(_02589_));
 sky130_fd_sc_hd__mux4_2 _25803_ (.A0(_02586_),
    .A1(_02587_),
    .A2(_02588_),
    .A3(_02589_),
    .S0(net522),
    .S1(net520),
    .X(_02590_));
 sky130_fd_sc_hd__mux4_2 _25804_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net528),
    .S1(net533),
    .X(_02591_));
 sky130_fd_sc_hd__mux4_2 _25805_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net527),
    .S1(net533),
    .X(_02592_));
 sky130_fd_sc_hd__mux4_2 _25806_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net527),
    .S1(net533),
    .X(_02593_));
 sky130_fd_sc_hd__mux4_2 _25807_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net528),
    .S1(net533),
    .X(_02594_));
 sky130_fd_sc_hd__mux4_2 _25808_ (.A0(_02591_),
    .A1(_02592_),
    .A2(_02593_),
    .A3(_02594_),
    .S0(net522),
    .S1(net520),
    .X(_02595_));
 sky130_fd_sc_hd__mux2i_4 _25809_ (.A0(_02590_),
    .A1(_02595_),
    .S(net518),
    .Y(_02596_));
 sky130_fd_sc_hd__xnor2_1 _25810_ (.A(_11220_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__xnor2_1 _25811_ (.A(_10928_),
    .B(_02597_),
    .Y(_11707_));
 sky130_fd_sc_hd__mux4_2 _25812_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net551),
    .S1(net552),
    .X(_02598_));
 sky130_fd_sc_hd__mux4_2 _25813_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net551),
    .S1(\count2_1[1] ),
    .X(_02599_));
 sky130_fd_sc_hd__mux4_2 _25814_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net551),
    .S1(\count2_1[1] ),
    .X(_02600_));
 sky130_fd_sc_hd__mux4_2 _25815_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net551),
    .S1(\count2_1[1] ),
    .X(_02601_));
 sky130_fd_sc_hd__mux4_2 _25816_ (.A0(_02598_),
    .A1(_02599_),
    .A2(_02600_),
    .A3(_02601_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02602_));
 sky130_fd_sc_hd__mux4_2 _25817_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_02603_));
 sky130_fd_sc_hd__mux4_2 _25818_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_02604_));
 sky130_fd_sc_hd__mux4_2 _25819_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_02605_));
 sky130_fd_sc_hd__mux4_2 _25820_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_02606_));
 sky130_fd_sc_hd__mux4_2 _25821_ (.A0(_02603_),
    .A1(_02604_),
    .A2(_02605_),
    .A3(_02606_),
    .S0(net442),
    .S1(net440),
    .X(_02607_));
 sky130_fd_sc_hd__mux2i_4 _25822_ (.A0(_02602_),
    .A1(_02607_),
    .S(net438),
    .Y(_02608_));
 sky130_fd_sc_hd__xnor2_1 _25823_ (.A(_11565_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__xnor2_1 _25824_ (.A(_11346_),
    .B(_02609_),
    .Y(_11712_));
 sky130_fd_sc_hd__xnor2_1 _25825_ (.A(_11022_),
    .B(_11266_),
    .Y(_02610_));
 sky130_fd_sc_hd__xnor2_1 _25826_ (.A(_10833_),
    .B(_02610_),
    .Y(_11715_));
 sky130_fd_sc_hd__mux4_2 _25827_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net551),
    .S1(net452),
    .X(_02611_));
 sky130_fd_sc_hd__mux4_2 _25828_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net551),
    .S1(net452),
    .X(_02612_));
 sky130_fd_sc_hd__mux4_2 _25829_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net551),
    .S1(net452),
    .X(_02613_));
 sky130_fd_sc_hd__mux4_2 _25830_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net551),
    .S1(net452),
    .X(_02614_));
 sky130_fd_sc_hd__mux4_2 _25831_ (.A0(_02611_),
    .A1(_02612_),
    .A2(_02613_),
    .A3(_02614_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02615_));
 sky130_fd_sc_hd__mux4_2 _25832_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net446),
    .S1(net552),
    .X(_02616_));
 sky130_fd_sc_hd__mux4_2 _25833_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net446),
    .S1(net552),
    .X(_02617_));
 sky130_fd_sc_hd__mux4_2 _25834_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net446),
    .S1(net552),
    .X(_02618_));
 sky130_fd_sc_hd__mux4_2 _25835_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net446),
    .S1(net552),
    .X(_02619_));
 sky130_fd_sc_hd__mux4_2 _25836_ (.A0(_02616_),
    .A1(_02617_),
    .A2(_02618_),
    .A3(_02619_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02620_));
 sky130_fd_sc_hd__mux2i_4 _25837_ (.A0(_02615_),
    .A1(_02620_),
    .S(\count2_1[5] ),
    .Y(_02621_));
 sky130_fd_sc_hd__xnor2_1 _25838_ (.A(_02584_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__xnor2_1 _25839_ (.A(_11381_),
    .B(_02622_),
    .Y(_11720_));
 sky130_fd_sc_hd__xnor2_1 _25840_ (.A(_11117_),
    .B(_11323_),
    .Y(_02623_));
 sky130_fd_sc_hd__xnor2_1 _25841_ (.A(_10905_),
    .B(_02623_),
    .Y(_11723_));
 sky130_fd_sc_hd__mux4_2 _25842_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net551),
    .S1(net452),
    .X(_02624_));
 sky130_fd_sc_hd__mux4_2 _25843_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net551),
    .S1(net452),
    .X(_02625_));
 sky130_fd_sc_hd__mux4_2 _25844_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net551),
    .S1(net452),
    .X(_02626_));
 sky130_fd_sc_hd__mux4_2 _25845_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net551),
    .S1(net452),
    .X(_02627_));
 sky130_fd_sc_hd__mux4_2 _25846_ (.A0(_02624_),
    .A1(_02625_),
    .A2(_02626_),
    .A3(_02627_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02628_));
 sky130_fd_sc_hd__mux4_2 _25847_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net446),
    .S1(net552),
    .X(_02629_));
 sky130_fd_sc_hd__mux4_2 _25848_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net446),
    .S1(net552),
    .X(_02630_));
 sky130_fd_sc_hd__mux4_2 _25849_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net446),
    .S1(net552),
    .X(_02631_));
 sky130_fd_sc_hd__mux4_2 _25850_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net446),
    .S1(net552),
    .X(_02632_));
 sky130_fd_sc_hd__mux4_2 _25851_ (.A0(_02629_),
    .A1(_02630_),
    .A2(_02631_),
    .A3(_02632_),
    .S0(net443),
    .S1(net550),
    .X(_02633_));
 sky130_fd_sc_hd__mux2i_4 _25852_ (.A0(_02628_),
    .A1(_02633_),
    .S(net438),
    .Y(_02634_));
 sky130_fd_sc_hd__xnor2_1 _25853_ (.A(_02608_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__xnor2_1 _25854_ (.A(_11416_),
    .B(_02635_),
    .Y(_11728_));
 sky130_fd_sc_hd__xnor2_1 _25855_ (.A(_11172_),
    .B(_11358_),
    .Y(_02636_));
 sky130_fd_sc_hd__xnor2_2 _25856_ (.A(_11034_),
    .B(_02636_),
    .Y(_11731_));
 sky130_fd_sc_hd__mux4_2 _25857_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net551),
    .S1(\count2_1[1] ),
    .X(_02637_));
 sky130_fd_sc_hd__mux4_2 _25858_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net551),
    .S1(\count2_1[1] ),
    .X(_02638_));
 sky130_fd_sc_hd__mux4_2 _25859_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net551),
    .S1(\count2_1[1] ),
    .X(_02639_));
 sky130_fd_sc_hd__mux4_2 _25860_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net551),
    .S1(net452),
    .X(_02640_));
 sky130_fd_sc_hd__mux4_2 _25861_ (.A0(_02637_),
    .A1(_02638_),
    .A2(_02639_),
    .A3(_02640_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02641_));
 sky130_fd_sc_hd__mux4_2 _25862_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net446),
    .S1(net456),
    .X(_02642_));
 sky130_fd_sc_hd__mux4_2 _25863_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net446),
    .S1(net456),
    .X(_02643_));
 sky130_fd_sc_hd__mux4_2 _25864_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net551),
    .S1(net456),
    .X(_02644_));
 sky130_fd_sc_hd__mux4_2 _25865_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count2_1[2] ),
    .S1(net456),
    .X(_02645_));
 sky130_fd_sc_hd__mux4_2 _25866_ (.A0(_02642_),
    .A1(_02643_),
    .A2(_02644_),
    .A3(_02645_),
    .S0(net443),
    .S1(\count2_1[4] ),
    .X(_02646_));
 sky130_fd_sc_hd__mux2i_4 _25867_ (.A0(_02641_),
    .A1(_02646_),
    .S(net438),
    .Y(_02647_));
 sky130_fd_sc_hd__xnor2_1 _25868_ (.A(_02621_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__xnor2_1 _25869_ (.A(_11451_),
    .B(_02648_),
    .Y(_11736_));
 sky130_fd_sc_hd__xnor2_1 _25870_ (.A(_11220_),
    .B(_11393_),
    .Y(_02649_));
 sky130_fd_sc_hd__xnor2_2 _25871_ (.A(_11104_),
    .B(_02649_),
    .Y(_11739_));
 sky130_fd_sc_hd__mux4_2 _25872_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net445),
    .S1(net451),
    .X(_02650_));
 sky130_fd_sc_hd__mux4_2 _25873_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net445),
    .S1(net451),
    .X(_02651_));
 sky130_fd_sc_hd__mux4_2 _25874_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net445),
    .S1(net451),
    .X(_02652_));
 sky130_fd_sc_hd__mux4_2 _25875_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net445),
    .S1(net451),
    .X(_02653_));
 sky130_fd_sc_hd__mux4_2 _25876_ (.A0(_02650_),
    .A1(_02651_),
    .A2(_02652_),
    .A3(_02653_),
    .S0(net443),
    .S1(net550),
    .X(_02654_));
 sky130_fd_sc_hd__mux4_2 _25877_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net450),
    .S1(net456),
    .X(_02655_));
 sky130_fd_sc_hd__mux4_2 _25878_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net450),
    .S1(net456),
    .X(_02656_));
 sky130_fd_sc_hd__mux4_2 _25879_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net450),
    .S1(net456),
    .X(_02657_));
 sky130_fd_sc_hd__mux4_2 _25880_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net450),
    .S1(net456),
    .X(_02658_));
 sky130_fd_sc_hd__mux4_2 _25881_ (.A0(_02655_),
    .A1(_02656_),
    .A2(_02657_),
    .A3(_02658_),
    .S0(net442),
    .S1(net440),
    .X(_02659_));
 sky130_fd_sc_hd__mux2i_2 _25882_ (.A0(_02654_),
    .A1(_02659_),
    .S(net438),
    .Y(_02660_));
 sky130_fd_sc_hd__xnor2_1 _25883_ (.A(_02634_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__xnor2_1 _25884_ (.A(_11475_),
    .B(_02661_),
    .Y(_11744_));
 sky130_fd_sc_hd__xnor2_1 _25885_ (.A(_11266_),
    .B(_11439_),
    .Y(_02662_));
 sky130_fd_sc_hd__xnor2_2 _25886_ (.A(_10893_),
    .B(_02662_),
    .Y(_11747_));
 sky130_fd_sc_hd__mux4_2 _25887_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02663_));
 sky130_fd_sc_hd__mux4_2 _25888_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02664_));
 sky130_fd_sc_hd__mux4_2 _25889_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02665_));
 sky130_fd_sc_hd__mux4_2 _25890_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02666_));
 sky130_fd_sc_hd__mux4_2 _25891_ (.A0(_02663_),
    .A1(_02664_),
    .A2(_02665_),
    .A3(_02666_),
    .S0(net441),
    .S1(net439),
    .X(_02667_));
 sky130_fd_sc_hd__mux4_2 _25892_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02668_));
 sky130_fd_sc_hd__mux4_2 _25893_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02669_));
 sky130_fd_sc_hd__mux4_2 _25894_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02670_));
 sky130_fd_sc_hd__mux4_2 _25895_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net447),
    .S1(net453),
    .X(_02671_));
 sky130_fd_sc_hd__mux4_2 _25896_ (.A0(_02668_),
    .A1(_02669_),
    .A2(_02670_),
    .A3(_02671_),
    .S0(net442),
    .S1(net440),
    .X(_02672_));
 sky130_fd_sc_hd__mux2i_4 _25897_ (.A0(_02667_),
    .A1(_02672_),
    .S(net437),
    .Y(_02673_));
 sky130_fd_sc_hd__xnor2_1 _25898_ (.A(_02647_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__xnor2_1 _25899_ (.A(_11499_),
    .B(_02674_),
    .Y(_11752_));
 sky130_fd_sc_hd__xnor2_1 _25900_ (.A(_11323_),
    .B(_11463_),
    .Y(_02675_));
 sky130_fd_sc_hd__xnor2_1 _25901_ (.A(_10917_),
    .B(_02675_),
    .Y(_11755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_269 ();
 sky130_fd_sc_hd__mux4_2 _25903_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02677_));
 sky130_fd_sc_hd__mux4_2 _25904_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02678_));
 sky130_fd_sc_hd__mux4_2 _25905_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02679_));
 sky130_fd_sc_hd__mux4_2 _25906_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02680_));
 sky130_fd_sc_hd__mux4_2 _25907_ (.A0(_02677_),
    .A1(_02678_),
    .A2(_02679_),
    .A3(_02680_),
    .S0(net441),
    .S1(net439),
    .X(_02681_));
 sky130_fd_sc_hd__mux4_2 _25908_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02682_));
 sky130_fd_sc_hd__mux4_2 _25909_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02683_));
 sky130_fd_sc_hd__mux4_2 _25910_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02684_));
 sky130_fd_sc_hd__mux4_2 _25911_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net447),
    .S1(net453),
    .X(_02685_));
 sky130_fd_sc_hd__mux4_2 _25912_ (.A0(_02682_),
    .A1(_02683_),
    .A2(_02684_),
    .A3(_02685_),
    .S0(net441),
    .S1(net439),
    .X(_02686_));
 sky130_fd_sc_hd__mux2i_4 _25913_ (.A0(_02681_),
    .A1(_02686_),
    .S(net437),
    .Y(_02687_));
 sky130_fd_sc_hd__xnor2_1 _25914_ (.A(_02660_),
    .B(_02687_),
    .Y(_11760_));
 sky130_fd_sc_hd__xnor2_1 _25915_ (.A(_11358_),
    .B(_11487_),
    .Y(_02688_));
 sky130_fd_sc_hd__xnor2_1 _25916_ (.A(_11045_),
    .B(_02688_),
    .Y(_11763_));
 sky130_fd_sc_hd__mux4_2 _25917_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net447),
    .S1(net453),
    .X(_02689_));
 sky130_fd_sc_hd__mux4_2 _25918_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net447),
    .S1(net453),
    .X(_02690_));
 sky130_fd_sc_hd__mux4_2 _25919_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net447),
    .S1(net453),
    .X(_02691_));
 sky130_fd_sc_hd__mux4_2 _25920_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net447),
    .S1(net453),
    .X(_02692_));
 sky130_fd_sc_hd__mux4_2 _25921_ (.A0(_02689_),
    .A1(_02690_),
    .A2(_02691_),
    .A3(_02692_),
    .S0(net441),
    .S1(net439),
    .X(_02693_));
 sky130_fd_sc_hd__mux4_2 _25922_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net449),
    .S1(net455),
    .X(_02694_));
 sky130_fd_sc_hd__mux4_2 _25923_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net449),
    .S1(net455),
    .X(_02695_));
 sky130_fd_sc_hd__mux4_2 _25924_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net449),
    .S1(net455),
    .X(_02696_));
 sky130_fd_sc_hd__mux4_2 _25925_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net449),
    .S1(net455),
    .X(_02697_));
 sky130_fd_sc_hd__mux4_2 _25926_ (.A0(_02694_),
    .A1(_02695_),
    .A2(_02696_),
    .A3(_02697_),
    .S0(net441),
    .S1(net439),
    .X(_02698_));
 sky130_fd_sc_hd__mux2i_4 _25927_ (.A0(_02693_),
    .A1(_02698_),
    .S(net437),
    .Y(_02699_));
 sky130_fd_sc_hd__xnor2_1 _25928_ (.A(_02673_),
    .B(_02699_),
    .Y(_11768_));
 sky130_fd_sc_hd__xnor2_1 _25929_ (.A(_11393_),
    .B(_11511_),
    .Y(_02700_));
 sky130_fd_sc_hd__xnor2_1 _25930_ (.A(_11129_),
    .B(_02700_),
    .Y(_11771_));
 sky130_fd_sc_hd__xnor2_1 _25931_ (.A(_10963_),
    .B(_02687_),
    .Y(_11776_));
 sky130_fd_sc_hd__xnor2_1 _25932_ (.A(_11439_),
    .B(_11553_),
    .Y(_02701_));
 sky130_fd_sc_hd__xnor2_1 _25933_ (.A(_11184_),
    .B(_02701_),
    .Y(_11779_));
 sky130_fd_sc_hd__xnor2_1 _25934_ (.A(_11057_),
    .B(_02699_),
    .Y(_11784_));
 sky130_fd_sc_hd__xnor2_1 _25935_ (.A(_11463_),
    .B(_02572_),
    .Y(_02702_));
 sky130_fd_sc_hd__xnor2_1 _25936_ (.A(_11231_),
    .B(_02702_),
    .Y(_11787_));
 sky130_fd_sc_hd__xnor2_1 _25937_ (.A(_10963_),
    .B(_11147_),
    .Y(_11792_));
 sky130_fd_sc_hd__xnor2_1 _25938_ (.A(_11487_),
    .B(_02596_),
    .Y(_02703_));
 sky130_fd_sc_hd__xnor2_1 _25939_ (.A(_11277_),
    .B(_02703_),
    .Y(_11795_));
 sky130_fd_sc_hd__xnor2_1 _25940_ (.A(_11057_),
    .B(_11196_),
    .Y(_11800_));
 sky130_fd_sc_hd__xnor2_1 _25941_ (.A(_11312_),
    .B(_11511_),
    .Y(_02704_));
 sky130_fd_sc_hd__xnor2_1 _25942_ (.A(_10833_),
    .B(_02704_),
    .Y(_11803_));
 sky130_fd_sc_hd__xnor2_1 _25943_ (.A(_11147_),
    .B(_11243_),
    .Y(_11808_));
 sky130_fd_sc_hd__xnor2_1 _25944_ (.A(_10905_),
    .B(_11369_),
    .Y(_11811_));
 sky130_fd_sc_hd__xnor2_1 _25945_ (.A(_11196_),
    .B(_11300_),
    .Y(_11816_));
 sky130_fd_sc_hd__xnor2_1 _25946_ (.A(_11034_),
    .B(_11404_),
    .Y(_11819_));
 sky130_fd_sc_hd__xnor2_1 _25947_ (.A(_11243_),
    .B(_11335_),
    .Y(_11824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_260 ();
 sky130_fd_sc_hd__mux4_2 _25957_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_258 ();
 sky130_fd_sc_hd__mux4_2 _25960_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02717_));
 sky130_fd_sc_hd__mux4_2 _25961_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02718_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_255 ();
 sky130_fd_sc_hd__mux4_2 _25965_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_250 ();
 sky130_fd_sc_hd__mux4_2 _25971_ (.A0(_02714_),
    .A1(_02717_),
    .A2(_02718_),
    .A3(_02722_),
    .S0(net422),
    .S1(net420),
    .X(_02728_));
 sky130_fd_sc_hd__mux4_2 _25972_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02729_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_248 ();
 sky130_fd_sc_hd__mux4_2 _25975_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02732_));
 sky130_fd_sc_hd__mux4_2 _25976_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02733_));
 sky130_fd_sc_hd__mux4_2 _25977_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net428),
    .S1(net434),
    .X(_02734_));
 sky130_fd_sc_hd__mux4_2 _25978_ (.A0(_02729_),
    .A1(_02732_),
    .A2(_02733_),
    .A3(_02734_),
    .S0(net422),
    .S1(net420),
    .X(_02735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_246 ();
 sky130_fd_sc_hd__mux2i_4 _25981_ (.A0(_02728_),
    .A1(_02735_),
    .S(net418),
    .Y(_02738_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_243 ();
 sky130_fd_sc_hd__mux4_2 _25985_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net427),
    .S1(net432),
    .X(_02742_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_241 ();
 sky130_fd_sc_hd__mux4_2 _25988_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net427),
    .S1(net432),
    .X(_02745_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_239 ();
 sky130_fd_sc_hd__mux4_2 _25991_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net427),
    .S1(net432),
    .X(_02748_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_237 ();
 sky130_fd_sc_hd__mux4_2 _25994_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net427),
    .S1(net432),
    .X(_02751_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_235 ();
 sky130_fd_sc_hd__mux4_2 _25997_ (.A0(_02742_),
    .A1(_02745_),
    .A2(_02748_),
    .A3(_02751_),
    .S0(net423),
    .S1(net421),
    .X(_02754_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_234 ();
 sky130_fd_sc_hd__mux4_2 _25999_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net428),
    .S1(net433),
    .X(_02756_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_232 ();
 sky130_fd_sc_hd__mux4_2 _26002_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net428),
    .S1(net433),
    .X(_02759_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_230 ();
 sky130_fd_sc_hd__mux4_2 _26005_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net428),
    .S1(net433),
    .X(_02762_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_228 ();
 sky130_fd_sc_hd__mux4_2 _26008_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net428),
    .S1(net433),
    .X(_02765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_226 ();
 sky130_fd_sc_hd__mux4_2 _26011_ (.A0(_02756_),
    .A1(_02759_),
    .A2(_02762_),
    .A3(_02765_),
    .S0(net422),
    .S1(net420),
    .X(_02768_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_225 ();
 sky130_fd_sc_hd__mux2i_4 _26013_ (.A0(_02754_),
    .A1(_02768_),
    .S(net418),
    .Y(_02770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_224 ();
 sky130_fd_sc_hd__mux4_2 _26015_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net426),
    .S1(net431),
    .X(_02772_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_222 ();
 sky130_fd_sc_hd__mux4_2 _26018_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net424),
    .S1(net435),
    .X(_02775_));
 sky130_fd_sc_hd__mux4_2 _26019_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net426),
    .S1(net431),
    .X(_02776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_220 ();
 sky130_fd_sc_hd__mux4_2 _26022_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net426),
    .S1(net431),
    .X(_02779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_218 ();
 sky130_fd_sc_hd__mux4_2 _26025_ (.A0(_02772_),
    .A1(_02775_),
    .A2(_02776_),
    .A3(_02779_),
    .S0(net549),
    .S1(net421),
    .X(_02782_));
 sky130_fd_sc_hd__mux4_2 _26026_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net429),
    .S1(net431),
    .X(_02783_));
 sky130_fd_sc_hd__mux4_2 _26027_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net429),
    .S1(net431),
    .X(_02784_));
 sky130_fd_sc_hd__mux4_2 _26028_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net429),
    .S1(net431),
    .X(_02785_));
 sky130_fd_sc_hd__mux4_2 _26029_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net429),
    .S1(net432),
    .X(_02786_));
 sky130_fd_sc_hd__mux4_2 _26030_ (.A0(_02783_),
    .A1(_02784_),
    .A2(_02785_),
    .A3(_02786_),
    .S0(net423),
    .S1(net421),
    .X(_02787_));
 sky130_fd_sc_hd__mux2i_4 _26031_ (.A0(_02782_),
    .A1(_02787_),
    .S(\count2_2[5] ),
    .Y(_02788_));
 sky130_fd_sc_hd__xnor2_1 _26032_ (.A(_02770_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__xnor2_1 _26033_ (.A(_02738_),
    .B(_02789_),
    .Y(_11829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__mux4_2 _26043_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net557),
    .S1(net517),
    .X(_02799_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_205 ();
 sky130_fd_sc_hd__mux4_2 _26048_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net557),
    .S1(net517),
    .X(_02804_));
 sky130_fd_sc_hd__mux4_2 _26049_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net557),
    .S1(net517),
    .X(_02805_));
 sky130_fd_sc_hd__mux4_2 _26050_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net557),
    .S1(net517),
    .X(_02806_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_200 ();
 sky130_fd_sc_hd__mux4_2 _26056_ (.A0(_02799_),
    .A1(_02804_),
    .A2(_02805_),
    .A3(_02806_),
    .S0(net504),
    .S1(net501),
    .X(_02812_));
 sky130_fd_sc_hd__mux4_2 _26057_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net511),
    .S1(net516),
    .X(_02813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_196 ();
 sky130_fd_sc_hd__mux4_2 _26062_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net511),
    .S1(net516),
    .X(_02818_));
 sky130_fd_sc_hd__mux4_2 _26063_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net511),
    .S1(net516),
    .X(_02819_));
 sky130_fd_sc_hd__mux4_2 _26064_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net511),
    .S1(net516),
    .X(_02820_));
 sky130_fd_sc_hd__mux4_2 _26065_ (.A0(_02813_),
    .A1(_02818_),
    .A2(_02819_),
    .A3(_02820_),
    .S0(\count15_2[3] ),
    .S1(net501),
    .X(_02821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_194 ();
 sky130_fd_sc_hd__mux2i_4 _26068_ (.A0(_02812_),
    .A1(_02821_),
    .S(net498),
    .Y(_02824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_192 ();
 sky130_fd_sc_hd__mux4_2 _26071_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net509),
    .S1(net514),
    .X(_02827_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_190 ();
 sky130_fd_sc_hd__mux4_2 _26074_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net509),
    .S1(net514),
    .X(_02830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_188 ();
 sky130_fd_sc_hd__mux4_2 _26077_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net509),
    .S1(net514),
    .X(_02833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_186 ();
 sky130_fd_sc_hd__mux4_2 _26080_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net509),
    .S1(net514),
    .X(_02836_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_184 ();
 sky130_fd_sc_hd__mux4_2 _26083_ (.A0(_02827_),
    .A1(_02830_),
    .A2(_02833_),
    .A3(_02836_),
    .S0(net503),
    .S1(net500),
    .X(_02839_));
 sky130_fd_sc_hd__mux4_2 _26084_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net510),
    .S1(net514),
    .X(_02840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_183 ();
 sky130_fd_sc_hd__mux4_2 _26086_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net510),
    .S1(net514),
    .X(_02842_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_181 ();
 sky130_fd_sc_hd__mux4_2 _26089_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net510),
    .S1(net514),
    .X(_02845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_179 ();
 sky130_fd_sc_hd__mux4_2 _26092_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net510),
    .S1(net514),
    .X(_02848_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_177 ();
 sky130_fd_sc_hd__mux4_2 _26095_ (.A0(_02840_),
    .A1(_02842_),
    .A2(_02845_),
    .A3(_02848_),
    .S0(net503),
    .S1(net500),
    .X(_02851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_176 ();
 sky130_fd_sc_hd__mux2i_4 _26097_ (.A0(_02839_),
    .A1(_02851_),
    .S(net498),
    .Y(_02853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_174 ();
 sky130_fd_sc_hd__mux4_2 _26100_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net511),
    .S1(net515),
    .X(_02856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_172 ();
 sky130_fd_sc_hd__mux4_2 _26103_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net511),
    .S1(net515),
    .X(_02859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_171 ();
 sky130_fd_sc_hd__mux4_2 _26105_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net511),
    .S1(net515),
    .X(_02861_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_170 ();
 sky130_fd_sc_hd__mux4_2 _26107_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net511),
    .S1(net515),
    .X(_02863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_168 ();
 sky130_fd_sc_hd__mux4_2 _26110_ (.A0(_02856_),
    .A1(_02859_),
    .A2(_02861_),
    .A3(_02863_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_02866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_166 ();
 sky130_fd_sc_hd__mux4_2 _26113_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net510),
    .S1(net516),
    .X(_02869_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_164 ();
 sky130_fd_sc_hd__mux4_2 _26116_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net510),
    .S1(net516),
    .X(_02872_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_162 ();
 sky130_fd_sc_hd__mux4_2 _26119_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net511),
    .S1(net516),
    .X(_02875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_160 ();
 sky130_fd_sc_hd__mux4_2 _26122_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net510),
    .S1(net516),
    .X(_02878_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_158 ();
 sky130_fd_sc_hd__mux4_2 _26125_ (.A0(_02869_),
    .A1(_02872_),
    .A2(_02875_),
    .A3(_02878_),
    .S0(net503),
    .S1(net500),
    .X(_02881_));
 sky130_fd_sc_hd__mux2i_4 _26126_ (.A0(_02866_),
    .A1(_02881_),
    .S(net498),
    .Y(_02882_));
 sky130_fd_sc_hd__xnor2_1 _26127_ (.A(_02853_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__xnor2_2 _26128_ (.A(_02824_),
    .B(_02883_),
    .Y(_11828_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_150 ();
 sky130_fd_sc_hd__mux4_2 _26137_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_146 ();
 sky130_fd_sc_hd__mux4_2 _26142_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02897_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_144 ();
 sky130_fd_sc_hd__mux4_2 _26145_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_141 ();
 sky130_fd_sc_hd__mux4_2 _26149_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_136 ();
 sky130_fd_sc_hd__mux4_2 _26155_ (.A0(_02892_),
    .A1(_02897_),
    .A2(_02900_),
    .A3(_02904_),
    .S0(net384),
    .S1(net542),
    .X(_02910_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_134 ();
 sky130_fd_sc_hd__mux4_2 _26158_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__mux4_2 _26161_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02916_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__mux4_2 _26164_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02919_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_128 ();
 sky130_fd_sc_hd__mux4_2 _26167_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net390),
    .S1(net395),
    .X(_02922_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_126 ();
 sky130_fd_sc_hd__mux4_2 _26170_ (.A0(_02913_),
    .A1(_02916_),
    .A2(_02919_),
    .A3(_02922_),
    .S0(net384),
    .S1(net542),
    .X(_02925_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_124 ();
 sky130_fd_sc_hd__mux2i_4 _26173_ (.A0(_02910_),
    .A1(_02925_),
    .S(net380),
    .Y(_11827_));
 sky130_fd_sc_hd__mux4_2 _26174_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net427),
    .S1(net432),
    .X(_02928_));
 sky130_fd_sc_hd__mux4_2 _26175_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net427),
    .S1(net432),
    .X(_02929_));
 sky130_fd_sc_hd__mux4_2 _26176_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net427),
    .S1(net432),
    .X(_02930_));
 sky130_fd_sc_hd__mux4_2 _26177_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net427),
    .S1(net432),
    .X(_02931_));
 sky130_fd_sc_hd__mux4_2 _26178_ (.A0(_02928_),
    .A1(_02929_),
    .A2(_02930_),
    .A3(_02931_),
    .S0(net422),
    .S1(net420),
    .X(_02932_));
 sky130_fd_sc_hd__mux4_2 _26179_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net430),
    .S1(net434),
    .X(_02933_));
 sky130_fd_sc_hd__mux4_2 _26180_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net430),
    .S1(net434),
    .X(_02934_));
 sky130_fd_sc_hd__mux4_2 _26181_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net430),
    .S1(net434),
    .X(_02935_));
 sky130_fd_sc_hd__mux4_2 _26182_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net430),
    .S1(net434),
    .X(_02936_));
 sky130_fd_sc_hd__mux4_2 _26183_ (.A0(_02933_),
    .A1(_02934_),
    .A2(_02935_),
    .A3(_02936_),
    .S0(net422),
    .S1(net420),
    .X(_02937_));
 sky130_fd_sc_hd__mux2i_4 _26184_ (.A0(_02932_),
    .A1(_02937_),
    .S(net418),
    .Y(_02938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_123 ();
 sky130_fd_sc_hd__mux4_2 _26186_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02940_));
 sky130_fd_sc_hd__mux4_2 _26187_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02941_));
 sky130_fd_sc_hd__mux4_2 _26188_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02942_));
 sky130_fd_sc_hd__mux4_2 _26189_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02943_));
 sky130_fd_sc_hd__mux4_2 _26190_ (.A0(_02940_),
    .A1(_02941_),
    .A2(_02942_),
    .A3(_02943_),
    .S0(net423),
    .S1(net420),
    .X(_02944_));
 sky130_fd_sc_hd__mux4_2 _26191_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_122 ();
 sky130_fd_sc_hd__mux4_2 _26193_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02947_));
 sky130_fd_sc_hd__mux4_2 _26194_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02948_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_121 ();
 sky130_fd_sc_hd__mux4_2 _26196_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_02950_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_120 ();
 sky130_fd_sc_hd__mux4_2 _26198_ (.A0(_02945_),
    .A1(_02947_),
    .A2(_02948_),
    .A3(_02950_),
    .S0(net423),
    .S1(net420),
    .X(_02952_));
 sky130_fd_sc_hd__mux2i_4 _26199_ (.A0(_02944_),
    .A1(_02952_),
    .S(net418),
    .Y(_02953_));
 sky130_fd_sc_hd__mux4_2 _26200_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02954_));
 sky130_fd_sc_hd__mux4_2 _26201_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02955_));
 sky130_fd_sc_hd__mux4_2 _26202_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02956_));
 sky130_fd_sc_hd__mux4_2 _26203_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02957_));
 sky130_fd_sc_hd__mux4_2 _26204_ (.A0(_02954_),
    .A1(_02955_),
    .A2(_02956_),
    .A3(_02957_),
    .S0(net422),
    .S1(net420),
    .X(_02958_));
 sky130_fd_sc_hd__mux4_2 _26205_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02959_));
 sky130_fd_sc_hd__mux4_2 _26206_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02960_));
 sky130_fd_sc_hd__mux4_2 _26207_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02961_));
 sky130_fd_sc_hd__mux4_2 _26208_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net428),
    .S1(net434),
    .X(_02962_));
 sky130_fd_sc_hd__mux4_2 _26209_ (.A0(_02959_),
    .A1(_02960_),
    .A2(_02961_),
    .A3(_02962_),
    .S0(net422),
    .S1(net420),
    .X(_02963_));
 sky130_fd_sc_hd__mux2i_4 _26210_ (.A0(_02958_),
    .A1(_02963_),
    .S(net419),
    .Y(_02964_));
 sky130_fd_sc_hd__xnor2_1 _26211_ (.A(_02953_),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__xnor2_1 _26212_ (.A(_02938_),
    .B(_02965_),
    .Y(_11834_));
 sky130_fd_sc_hd__mux4_2 _26213_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net505),
    .S1(net517),
    .X(_02966_));
 sky130_fd_sc_hd__mux4_2 _26214_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net505),
    .S1(net517),
    .X(_02967_));
 sky130_fd_sc_hd__mux4_2 _26215_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net505),
    .S1(net517),
    .X(_02968_));
 sky130_fd_sc_hd__mux4_2 _26216_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net505),
    .S1(net517),
    .X(_02969_));
 sky130_fd_sc_hd__mux4_2 _26217_ (.A0(_02966_),
    .A1(_02967_),
    .A2(_02968_),
    .A3(_02969_),
    .S0(net504),
    .S1(net501),
    .X(_02970_));
 sky130_fd_sc_hd__mux4_2 _26218_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_02971_));
 sky130_fd_sc_hd__mux4_2 _26219_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_02972_));
 sky130_fd_sc_hd__mux4_2 _26220_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_02973_));
 sky130_fd_sc_hd__mux4_2 _26221_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_02974_));
 sky130_fd_sc_hd__mux4_2 _26222_ (.A0(_02971_),
    .A1(_02972_),
    .A2(_02973_),
    .A3(_02974_),
    .S0(net504),
    .S1(net501),
    .X(_02975_));
 sky130_fd_sc_hd__mux2i_4 _26223_ (.A0(_02970_),
    .A1(_02975_),
    .S(\count15_2[5] ),
    .Y(_02976_));
 sky130_fd_sc_hd__mux4_2 _26224_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_118 ();
 sky130_fd_sc_hd__mux4_2 _26227_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02980_));
 sky130_fd_sc_hd__mux4_2 _26228_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_117 ();
 sky130_fd_sc_hd__mux4_2 _26230_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02983_));
 sky130_fd_sc_hd__mux4_2 _26231_ (.A0(_02977_),
    .A1(_02980_),
    .A2(_02981_),
    .A3(_02983_),
    .S0(net502),
    .S1(net499),
    .X(_02984_));
 sky130_fd_sc_hd__mux4_2 _26232_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02985_));
 sky130_fd_sc_hd__mux4_2 _26233_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02986_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_115 ();
 sky130_fd_sc_hd__mux4_2 _26236_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_113 ();
 sky130_fd_sc_hd__mux4_2 _26239_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net507),
    .S1(net512),
    .X(_02992_));
 sky130_fd_sc_hd__mux4_2 _26240_ (.A0(_02985_),
    .A1(_02986_),
    .A2(_02989_),
    .A3(_02992_),
    .S0(net502),
    .S1(net499),
    .X(_02993_));
 sky130_fd_sc_hd__mux2i_4 _26241_ (.A0(_02984_),
    .A1(_02993_),
    .S(net497),
    .Y(_02994_));
 sky130_fd_sc_hd__mux4_2 _26242_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net508),
    .S1(net513),
    .X(_02995_));
 sky130_fd_sc_hd__mux4_2 _26243_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net508),
    .S1(net513),
    .X(_02996_));
 sky130_fd_sc_hd__mux4_2 _26244_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net508),
    .S1(net513),
    .X(_02997_));
 sky130_fd_sc_hd__mux4_2 _26245_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net508),
    .S1(net513),
    .X(_02998_));
 sky130_fd_sc_hd__mux4_2 _26246_ (.A0(_02995_),
    .A1(_02996_),
    .A2(_02997_),
    .A3(_02998_),
    .S0(net502),
    .S1(net499),
    .X(_02999_));
 sky130_fd_sc_hd__mux4_2 _26247_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net507),
    .S1(net512),
    .X(_03000_));
 sky130_fd_sc_hd__mux4_2 _26248_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net508),
    .S1(net513),
    .X(_03001_));
 sky130_fd_sc_hd__mux4_2 _26249_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net508),
    .S1(net513),
    .X(_03002_));
 sky130_fd_sc_hd__mux4_2 _26250_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net508),
    .S1(net513),
    .X(_03003_));
 sky130_fd_sc_hd__mux4_2 _26251_ (.A0(_03000_),
    .A1(_03001_),
    .A2(_03002_),
    .A3(_03003_),
    .S0(net503),
    .S1(net500),
    .X(_03004_));
 sky130_fd_sc_hd__mux2i_4 _26252_ (.A0(_02999_),
    .A1(_03004_),
    .S(net497),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor2_1 _26253_ (.A(net1131),
    .B(net1140),
    .Y(_03006_));
 sky130_fd_sc_hd__xnor2_2 _26254_ (.A(_02976_),
    .B(_03006_),
    .Y(_11833_));
 sky130_fd_sc_hd__mux4_2 _26255_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net387),
    .S1(net396),
    .X(_03007_));
 sky130_fd_sc_hd__mux4_2 _26256_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net387),
    .S1(net396),
    .X(_03008_));
 sky130_fd_sc_hd__mux4_2 _26257_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net387),
    .S1(net396),
    .X(_03009_));
 sky130_fd_sc_hd__mux4_2 _26258_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net387),
    .S1(net396),
    .X(_03010_));
 sky130_fd_sc_hd__mux4_2 _26259_ (.A0(_03007_),
    .A1(_03008_),
    .A2(_03009_),
    .A3(_03010_),
    .S0(net385),
    .S1(net382),
    .X(_03011_));
 sky130_fd_sc_hd__mux4_2 _26260_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net391),
    .S1(net397),
    .X(_03012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_112 ();
 sky130_fd_sc_hd__mux4_2 _26262_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net391),
    .S1(net397),
    .X(_03014_));
 sky130_fd_sc_hd__mux4_2 _26263_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net391),
    .S1(net397),
    .X(_03015_));
 sky130_fd_sc_hd__mux4_2 _26264_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net391),
    .S1(net397),
    .X(_03016_));
 sky130_fd_sc_hd__mux4_2 _26265_ (.A0(_03012_),
    .A1(_03014_),
    .A2(_03015_),
    .A3(_03016_),
    .S0(net384),
    .S1(net542),
    .X(_03017_));
 sky130_fd_sc_hd__mux2i_4 _26266_ (.A0(_03011_),
    .A1(_03017_),
    .S(net380),
    .Y(_11832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__mux4_2 _26275_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net465),
    .S1(net475),
    .X(_03026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__mux4_2 _26280_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net465),
    .S1(net475),
    .X(_03031_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_98 ();
 sky130_fd_sc_hd__mux4_2 _26283_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net465),
    .S1(net475),
    .X(_03034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_95 ();
 sky130_fd_sc_hd__mux4_2 _26287_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net465),
    .S1(net475),
    .X(_03038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_90 ();
 sky130_fd_sc_hd__mux4_2 _26293_ (.A0(_03026_),
    .A1(_03031_),
    .A2(_03034_),
    .A3(_03038_),
    .S0(net462),
    .S1(net460),
    .X(_03044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_88 ();
 sky130_fd_sc_hd__mux4_2 _26296_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net465),
    .S1(net476),
    .X(_03047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_86 ();
 sky130_fd_sc_hd__mux4_2 _26299_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net465),
    .S1(net476),
    .X(_03050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_84 ();
 sky130_fd_sc_hd__mux4_2 _26302_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net465),
    .S1(net476),
    .X(_03053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_82 ();
 sky130_fd_sc_hd__mux4_2 _26305_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net465),
    .S1(net476),
    .X(_03056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_80 ();
 sky130_fd_sc_hd__mux4_2 _26308_ (.A0(_03047_),
    .A1(_03050_),
    .A2(_03053_),
    .A3(_03056_),
    .S0(net462),
    .S1(net460),
    .X(_03059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_78 ();
 sky130_fd_sc_hd__mux2i_4 _26311_ (.A0(_03044_),
    .A1(_03059_),
    .S(net458),
    .Y(_11837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_77 ();
 sky130_fd_sc_hd__mux4_2 _26313_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net427),
    .S1(net432),
    .X(_03063_));
 sky130_fd_sc_hd__mux4_2 _26314_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net427),
    .S1(net432),
    .X(_03064_));
 sky130_fd_sc_hd__mux4_2 _26315_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net427),
    .S1(net432),
    .X(_03065_));
 sky130_fd_sc_hd__mux4_2 _26316_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net427),
    .S1(net432),
    .X(_03066_));
 sky130_fd_sc_hd__mux4_2 _26317_ (.A0(_03063_),
    .A1(_03064_),
    .A2(_03065_),
    .A3(_03066_),
    .S0(net422),
    .S1(net420),
    .X(_03067_));
 sky130_fd_sc_hd__mux4_2 _26318_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net428),
    .S1(net433),
    .X(_03068_));
 sky130_fd_sc_hd__mux4_2 _26319_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net428),
    .S1(net433),
    .X(_03069_));
 sky130_fd_sc_hd__mux4_2 _26320_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net429),
    .S1(net433),
    .X(_03070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_76 ();
 sky130_fd_sc_hd__mux4_2 _26322_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net428),
    .S1(net433),
    .X(_03072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__mux4_2 _26324_ (.A0(_03068_),
    .A1(_03069_),
    .A2(_03070_),
    .A3(_03072_),
    .S0(net422),
    .S1(net420),
    .X(_03074_));
 sky130_fd_sc_hd__mux2i_4 _26325_ (.A0(_03067_),
    .A1(_03074_),
    .S(net418),
    .Y(_03075_));
 sky130_fd_sc_hd__mux4_2 _26326_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03076_));
 sky130_fd_sc_hd__mux4_2 _26327_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03077_));
 sky130_fd_sc_hd__mux4_2 _26328_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03078_));
 sky130_fd_sc_hd__mux4_2 _26329_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03079_));
 sky130_fd_sc_hd__mux4_2 _26330_ (.A0(_03076_),
    .A1(_03077_),
    .A2(_03078_),
    .A3(_03079_),
    .S0(net422),
    .S1(net420),
    .X(_03080_));
 sky130_fd_sc_hd__mux4_2 _26331_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03081_));
 sky130_fd_sc_hd__mux4_2 _26332_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03082_));
 sky130_fd_sc_hd__mux4_2 _26333_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03083_));
 sky130_fd_sc_hd__mux4_2 _26334_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net428),
    .S1(net434),
    .X(_03084_));
 sky130_fd_sc_hd__mux4_2 _26335_ (.A0(_03081_),
    .A1(_03082_),
    .A2(_03083_),
    .A3(_03084_),
    .S0(net422),
    .S1(net420),
    .X(_03085_));
 sky130_fd_sc_hd__mux2i_4 _26336_ (.A0(_03080_),
    .A1(_03085_),
    .S(net418),
    .Y(_03086_));
 sky130_fd_sc_hd__xnor2_1 _26337_ (.A(_03075_),
    .B(_03086_),
    .Y(_03087_));
 sky130_fd_sc_hd__xnor2_1 _26338_ (.A(_02770_),
    .B(_03087_),
    .Y(_11842_));
 sky130_fd_sc_hd__mux4_2 _26339_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net505),
    .S1(net517),
    .X(_03088_));
 sky130_fd_sc_hd__mux4_2 _26340_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net505),
    .S1(net517),
    .X(_03089_));
 sky130_fd_sc_hd__mux4_2 _26341_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net505),
    .S1(net517),
    .X(_03090_));
 sky130_fd_sc_hd__mux4_2 _26342_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net505),
    .S1(net517),
    .X(_03091_));
 sky130_fd_sc_hd__mux4_2 _26343_ (.A0(_03088_),
    .A1(_03089_),
    .A2(_03090_),
    .A3(_03091_),
    .S0(net504),
    .S1(net501),
    .X(_03092_));
 sky130_fd_sc_hd__mux4_2 _26344_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03093_));
 sky130_fd_sc_hd__mux4_2 _26345_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03094_));
 sky130_fd_sc_hd__mux4_2 _26346_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03095_));
 sky130_fd_sc_hd__mux4_2 _26347_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03096_));
 sky130_fd_sc_hd__mux4_2 _26348_ (.A0(_03093_),
    .A1(_03094_),
    .A2(_03095_),
    .A3(_03096_),
    .S0(net504),
    .S1(net501),
    .X(_03097_));
 sky130_fd_sc_hd__mux2i_4 _26349_ (.A0(_03092_),
    .A1(_03097_),
    .S(\count15_2[5] ),
    .Y(_03098_));
 sky130_fd_sc_hd__mux4_2 _26350_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net507),
    .S1(net512),
    .X(_03099_));
 sky130_fd_sc_hd__mux4_2 _26351_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net507),
    .S1(net512),
    .X(_03100_));
 sky130_fd_sc_hd__mux4_2 _26352_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net507),
    .S1(net512),
    .X(_03101_));
 sky130_fd_sc_hd__mux4_2 _26353_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net507),
    .S1(net512),
    .X(_03102_));
 sky130_fd_sc_hd__mux4_2 _26354_ (.A0(_03099_),
    .A1(_03100_),
    .A2(_03101_),
    .A3(_03102_),
    .S0(net503),
    .S1(net500),
    .X(_03103_));
 sky130_fd_sc_hd__mux4_2 _26355_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net510),
    .S1(net514),
    .X(_03104_));
 sky130_fd_sc_hd__mux4_2 _26356_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net510),
    .S1(net514),
    .X(_03105_));
 sky130_fd_sc_hd__mux4_2 _26357_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net510),
    .S1(net514),
    .X(_03106_));
 sky130_fd_sc_hd__mux4_2 _26358_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net510),
    .S1(net514),
    .X(_03107_));
 sky130_fd_sc_hd__mux4_2 _26359_ (.A0(_03104_),
    .A1(_03105_),
    .A2(_03106_),
    .A3(_03107_),
    .S0(net503),
    .S1(net500),
    .X(_03108_));
 sky130_fd_sc_hd__mux2i_4 _26360_ (.A0(_03103_),
    .A1(_03108_),
    .S(net498),
    .Y(_03109_));
 sky130_fd_sc_hd__mux4_2 _26361_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03110_));
 sky130_fd_sc_hd__mux4_2 _26362_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03111_));
 sky130_fd_sc_hd__mux4_2 _26363_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03112_));
 sky130_fd_sc_hd__mux4_2 _26364_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03113_));
 sky130_fd_sc_hd__mux4_2 _26365_ (.A0(_03110_),
    .A1(_03111_),
    .A2(_03112_),
    .A3(_03113_),
    .S0(net503),
    .S1(net500),
    .X(_03114_));
 sky130_fd_sc_hd__mux4_2 _26366_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03115_));
 sky130_fd_sc_hd__mux4_2 _26367_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03116_));
 sky130_fd_sc_hd__mux4_2 _26368_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03117_));
 sky130_fd_sc_hd__mux4_2 _26369_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net507),
    .S1(net512),
    .X(_03118_));
 sky130_fd_sc_hd__mux4_2 _26370_ (.A0(_03115_),
    .A1(_03116_),
    .A2(_03117_),
    .A3(_03118_),
    .S0(net503),
    .S1(net500),
    .X(_03119_));
 sky130_fd_sc_hd__mux2i_4 _26371_ (.A0(_03114_),
    .A1(_03119_),
    .S(net497),
    .Y(_03120_));
 sky130_fd_sc_hd__xnor2_1 _26372_ (.A(_03109_),
    .B(net1130),
    .Y(_03121_));
 sky130_fd_sc_hd__xnor2_2 _26373_ (.A(_03098_),
    .B(_03121_),
    .Y(_11841_));
 sky130_fd_sc_hd__mux4_2 _26374_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_74 ();
 sky130_fd_sc_hd__mux4_2 _26376_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03124_));
 sky130_fd_sc_hd__mux4_2 _26377_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03125_));
 sky130_fd_sc_hd__mux4_2 _26378_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03126_));
 sky130_fd_sc_hd__mux4_2 _26379_ (.A0(_03122_),
    .A1(_03124_),
    .A2(_03125_),
    .A3(_03126_),
    .S0(net386),
    .S1(net383),
    .X(_03127_));
 sky130_fd_sc_hd__mux4_2 _26380_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__mux4_2 _26382_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03130_));
 sky130_fd_sc_hd__mux4_2 _26383_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03131_));
 sky130_fd_sc_hd__mux4_2 _26384_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net389),
    .S1(net394),
    .X(_03132_));
 sky130_fd_sc_hd__mux4_2 _26385_ (.A0(_03128_),
    .A1(_03130_),
    .A2(_03131_),
    .A3(_03132_),
    .S0(net386),
    .S1(net383),
    .X(_03133_));
 sky130_fd_sc_hd__mux2i_4 _26386_ (.A0(_03127_),
    .A1(_03133_),
    .S(\count7_2[5] ),
    .Y(_11840_));
 sky130_fd_sc_hd__mux4_2 _26387_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net465),
    .S1(net476),
    .X(_03134_));
 sky130_fd_sc_hd__mux4_2 _26388_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net465),
    .S1(net476),
    .X(_03135_));
 sky130_fd_sc_hd__mux4_2 _26389_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net465),
    .S1(net476),
    .X(_03136_));
 sky130_fd_sc_hd__mux4_2 _26390_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net465),
    .S1(net476),
    .X(_03137_));
 sky130_fd_sc_hd__mux4_2 _26391_ (.A0(_03134_),
    .A1(_03135_),
    .A2(_03136_),
    .A3(_03137_),
    .S0(net462),
    .S1(net460),
    .X(_03138_));
 sky130_fd_sc_hd__mux4_2 _26392_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net467),
    .S1(net474),
    .X(_03139_));
 sky130_fd_sc_hd__mux4_2 _26393_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net466),
    .S1(net474),
    .X(_03140_));
 sky130_fd_sc_hd__mux4_2 _26394_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net466),
    .S1(net474),
    .X(_03141_));
 sky130_fd_sc_hd__mux4_2 _26395_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net467),
    .S1(net476),
    .X(_03142_));
 sky130_fd_sc_hd__mux4_2 _26396_ (.A0(_03139_),
    .A1(_03140_),
    .A2(_03141_),
    .A3(_03142_),
    .S0(net463),
    .S1(net459),
    .X(_03143_));
 sky130_fd_sc_hd__mux2i_4 _26397_ (.A0(_03138_),
    .A1(_03143_),
    .S(net458),
    .Y(_11845_));
 sky130_fd_sc_hd__mux4_2 _26398_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__mux4_2 _26401_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03147_));
 sky130_fd_sc_hd__mux4_2 _26402_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03148_));
 sky130_fd_sc_hd__mux4_2 _26403_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03149_));
 sky130_fd_sc_hd__mux4_2 _26404_ (.A0(_03144_),
    .A1(_03147_),
    .A2(_03148_),
    .A3(_03149_),
    .S0(net422),
    .S1(net420),
    .X(_03150_));
 sky130_fd_sc_hd__mux4_2 _26405_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03151_));
 sky130_fd_sc_hd__mux4_2 _26406_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03152_));
 sky130_fd_sc_hd__mux4_2 _26407_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03153_));
 sky130_fd_sc_hd__mux4_2 _26408_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net428),
    .S1(net434),
    .X(_03154_));
 sky130_fd_sc_hd__mux4_2 _26409_ (.A0(_03151_),
    .A1(_03152_),
    .A2(_03153_),
    .A3(_03154_),
    .S0(net422),
    .S1(net420),
    .X(_03155_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_70 ();
 sky130_fd_sc_hd__mux2i_4 _26411_ (.A0(_03150_),
    .A1(_03155_),
    .S(net418),
    .Y(_03157_));
 sky130_fd_sc_hd__mux4_2 _26412_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net427),
    .S1(net434),
    .X(_03158_));
 sky130_fd_sc_hd__mux4_2 _26413_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net427),
    .S1(net434),
    .X(_03159_));
 sky130_fd_sc_hd__mux4_2 _26414_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net427),
    .S1(net434),
    .X(_03160_));
 sky130_fd_sc_hd__mux4_2 _26415_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net427),
    .S1(net434),
    .X(_03161_));
 sky130_fd_sc_hd__mux4_2 _26416_ (.A0(_03158_),
    .A1(_03159_),
    .A2(_03160_),
    .A3(_03161_),
    .S0(net422),
    .S1(net420),
    .X(_03162_));
 sky130_fd_sc_hd__mux4_2 _26417_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net427),
    .S1(net432),
    .X(_03163_));
 sky130_fd_sc_hd__mux4_2 _26418_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net427),
    .S1(net432),
    .X(_03164_));
 sky130_fd_sc_hd__mux4_2 _26419_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net427),
    .S1(net432),
    .X(_03165_));
 sky130_fd_sc_hd__mux4_2 _26420_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net427),
    .S1(net432),
    .X(_03166_));
 sky130_fd_sc_hd__mux4_2 _26421_ (.A0(_03163_),
    .A1(_03164_),
    .A2(_03165_),
    .A3(_03166_),
    .S0(net422),
    .S1(net420),
    .X(_03167_));
 sky130_fd_sc_hd__mux2i_4 _26422_ (.A0(_03162_),
    .A1(_03167_),
    .S(net419),
    .Y(_03168_));
 sky130_fd_sc_hd__xnor2_1 _26423_ (.A(_03157_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__xnor2_1 _26424_ (.A(_02953_),
    .B(_03169_),
    .Y(_11853_));
 sky130_fd_sc_hd__mux4_2 _26425_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net506),
    .S1(net515),
    .X(_03170_));
 sky130_fd_sc_hd__mux4_2 _26426_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net506),
    .S1(net515),
    .X(_03171_));
 sky130_fd_sc_hd__mux4_2 _26427_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net506),
    .S1(net515),
    .X(_03172_));
 sky130_fd_sc_hd__mux4_2 _26428_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net506),
    .S1(net515),
    .X(_03173_));
 sky130_fd_sc_hd__mux4_2 _26429_ (.A0(_03170_),
    .A1(_03171_),
    .A2(_03172_),
    .A3(_03173_),
    .S0(net502),
    .S1(net499),
    .X(_03174_));
 sky130_fd_sc_hd__mux4_2 _26430_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net508),
    .S1(net513),
    .X(_03175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_69 ();
 sky130_fd_sc_hd__mux4_2 _26432_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net509),
    .S1(net514),
    .X(_03177_));
 sky130_fd_sc_hd__mux4_2 _26433_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net509),
    .S1(net514),
    .X(_03178_));
 sky130_fd_sc_hd__mux4_2 _26434_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net509),
    .S1(net514),
    .X(_03179_));
 sky130_fd_sc_hd__mux4_2 _26435_ (.A0(_03175_),
    .A1(_03177_),
    .A2(_03178_),
    .A3(_03179_),
    .S0(net503),
    .S1(net500),
    .X(_03180_));
 sky130_fd_sc_hd__mux2i_4 _26436_ (.A0(_03174_),
    .A1(_03180_),
    .S(net497),
    .Y(_03181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_67 ();
 sky130_fd_sc_hd__mux4_2 _26439_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net557),
    .S1(net517),
    .X(_03184_));
 sky130_fd_sc_hd__mux4_2 _26440_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net557),
    .S1(net517),
    .X(_03185_));
 sky130_fd_sc_hd__mux4_2 _26441_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net557),
    .S1(net517),
    .X(_03186_));
 sky130_fd_sc_hd__mux4_2 _26442_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net505),
    .S1(net517),
    .X(_03187_));
 sky130_fd_sc_hd__mux4_2 _26443_ (.A0(_03184_),
    .A1(_03185_),
    .A2(_03186_),
    .A3(_03187_),
    .S0(net504),
    .S1(net501),
    .X(_03188_));
 sky130_fd_sc_hd__mux4_2 _26444_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net511),
    .S1(\count15_2[1] ),
    .X(_03189_));
 sky130_fd_sc_hd__mux4_2 _26445_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net511),
    .S1(\count15_2[1] ),
    .X(_03190_));
 sky130_fd_sc_hd__mux4_2 _26446_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net511),
    .S1(\count15_2[1] ),
    .X(_03191_));
 sky130_fd_sc_hd__mux4_2 _26447_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net511),
    .S1(\count15_2[1] ),
    .X(_03192_));
 sky130_fd_sc_hd__mux4_2 _26448_ (.A0(_03189_),
    .A1(_03190_),
    .A2(_03191_),
    .A3(_03192_),
    .S0(\count15_2[3] ),
    .S1(net501),
    .X(_03193_));
 sky130_fd_sc_hd__mux2i_4 _26449_ (.A0(_03188_),
    .A1(_03193_),
    .S(\count15_2[5] ),
    .Y(_03194_));
 sky130_fd_sc_hd__mux4_2 _26450_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net507),
    .S1(net512),
    .X(_03195_));
 sky130_fd_sc_hd__mux4_2 _26451_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net507),
    .S1(net512),
    .X(_03196_));
 sky130_fd_sc_hd__mux4_2 _26452_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net507),
    .S1(net512),
    .X(_03197_));
 sky130_fd_sc_hd__mux4_2 _26453_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net507),
    .S1(net512),
    .X(_03198_));
 sky130_fd_sc_hd__mux4_2 _26454_ (.A0(_03195_),
    .A1(_03196_),
    .A2(_03197_),
    .A3(_03198_),
    .S0(net503),
    .S1(net500),
    .X(_03199_));
 sky130_fd_sc_hd__mux4_2 _26455_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net509),
    .S1(net514),
    .X(_03200_));
 sky130_fd_sc_hd__mux4_2 _26456_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net509),
    .S1(net514),
    .X(_03201_));
 sky130_fd_sc_hd__mux4_2 _26457_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net509),
    .S1(net514),
    .X(_03202_));
 sky130_fd_sc_hd__mux4_2 _26458_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net509),
    .S1(net514),
    .X(_03203_));
 sky130_fd_sc_hd__mux4_2 _26459_ (.A0(_03200_),
    .A1(_03201_),
    .A2(_03202_),
    .A3(_03203_),
    .S0(net503),
    .S1(net500),
    .X(_03204_));
 sky130_fd_sc_hd__mux2i_4 _26460_ (.A0(_03199_),
    .A1(_03204_),
    .S(net497),
    .Y(_03205_));
 sky130_fd_sc_hd__xnor2_1 _26461_ (.A(_03194_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__xnor2_2 _26462_ (.A(_03181_),
    .B(_03206_),
    .Y(_11852_));
 sky130_fd_sc_hd__mux4_2 _26463_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net543),
    .S1(\count7_2[1] ),
    .X(_03207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_66 ();
 sky130_fd_sc_hd__mux4_2 _26465_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net543),
    .S1(\count7_2[1] ),
    .X(_03209_));
 sky130_fd_sc_hd__mux4_2 _26466_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net543),
    .S1(\count7_2[1] ),
    .X(_03210_));
 sky130_fd_sc_hd__mux4_2 _26467_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net543),
    .S1(\count7_2[1] ),
    .X(_03211_));
 sky130_fd_sc_hd__mux4_2 _26468_ (.A0(_03207_),
    .A1(_03209_),
    .A2(_03210_),
    .A3(_03211_),
    .S0(\count7_2[3] ),
    .S1(net383),
    .X(_03212_));
 sky130_fd_sc_hd__mux4_2 _26469_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net393),
    .S1(net544),
    .X(_03213_));
 sky130_fd_sc_hd__mux4_2 _26470_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net393),
    .S1(net544),
    .X(_03214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_65 ();
 sky130_fd_sc_hd__mux4_2 _26472_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net393),
    .S1(net544),
    .X(_03216_));
 sky130_fd_sc_hd__mux4_2 _26473_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net393),
    .S1(net544),
    .X(_03217_));
 sky130_fd_sc_hd__mux4_2 _26474_ (.A0(_03213_),
    .A1(_03214_),
    .A2(_03216_),
    .A3(_03217_),
    .S0(net385),
    .S1(net383),
    .X(_03218_));
 sky130_fd_sc_hd__mux2i_4 _26475_ (.A0(_03212_),
    .A1(_03218_),
    .S(net381),
    .Y(_11851_));
 sky130_fd_sc_hd__mux4_2 _26476_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03219_));
 sky130_fd_sc_hd__mux4_2 _26477_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03220_));
 sky130_fd_sc_hd__mux4_2 _26478_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03221_));
 sky130_fd_sc_hd__mux4_2 _26479_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03222_));
 sky130_fd_sc_hd__mux4_2 _26480_ (.A0(_03219_),
    .A1(_03220_),
    .A2(_03221_),
    .A3(_03222_),
    .S0(net462),
    .S1(net460),
    .X(_03223_));
 sky130_fd_sc_hd__mux4_2 _26481_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03224_));
 sky130_fd_sc_hd__mux4_2 _26482_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03225_));
 sky130_fd_sc_hd__mux4_2 _26483_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03226_));
 sky130_fd_sc_hd__mux4_2 _26484_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net468),
    .S1(net475),
    .X(_03227_));
 sky130_fd_sc_hd__mux4_2 _26485_ (.A0(_03224_),
    .A1(_03225_),
    .A2(_03226_),
    .A3(_03227_),
    .S0(net464),
    .S1(net461),
    .X(_03228_));
 sky130_fd_sc_hd__mux2i_4 _26486_ (.A0(_03223_),
    .A1(_03228_),
    .S(\count16_2[5] ),
    .Y(_11856_));
 sky130_fd_sc_hd__mux4_2 _26487_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03229_));
 sky130_fd_sc_hd__mux4_2 _26488_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03230_));
 sky130_fd_sc_hd__mux4_2 _26489_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03231_));
 sky130_fd_sc_hd__mux4_2 _26490_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03232_));
 sky130_fd_sc_hd__mux4_2 _26491_ (.A0(_03229_),
    .A1(_03230_),
    .A2(_03231_),
    .A3(_03232_),
    .S0(net423),
    .S1(net421),
    .X(_03233_));
 sky130_fd_sc_hd__mux4_2 _26492_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03234_));
 sky130_fd_sc_hd__mux4_2 _26493_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03235_));
 sky130_fd_sc_hd__mux4_2 _26494_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03236_));
 sky130_fd_sc_hd__mux4_2 _26495_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net427),
    .S1(net432),
    .X(_03237_));
 sky130_fd_sc_hd__mux4_2 _26496_ (.A0(_03234_),
    .A1(_03235_),
    .A2(_03236_),
    .A3(_03237_),
    .S0(net422),
    .S1(net420),
    .X(_03238_));
 sky130_fd_sc_hd__mux2i_4 _26497_ (.A0(_03233_),
    .A1(_03238_),
    .S(net419),
    .Y(_03239_));
 sky130_fd_sc_hd__mux4_2 _26498_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net425),
    .S1(net436),
    .X(_03240_));
 sky130_fd_sc_hd__mux4_2 _26499_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net425),
    .S1(net436),
    .X(_03241_));
 sky130_fd_sc_hd__mux4_2 _26500_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net425),
    .S1(net436),
    .X(_03242_));
 sky130_fd_sc_hd__mux4_2 _26501_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net425),
    .S1(net436),
    .X(_03243_));
 sky130_fd_sc_hd__mux4_2 _26502_ (.A0(_03240_),
    .A1(_03241_),
    .A2(_03242_),
    .A3(_03243_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_03244_));
 sky130_fd_sc_hd__mux4_2 _26503_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net429),
    .S1(net433),
    .X(_03245_));
 sky130_fd_sc_hd__mux4_2 _26504_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net429),
    .S1(net433),
    .X(_03246_));
 sky130_fd_sc_hd__mux4_2 _26505_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net429),
    .S1(net433),
    .X(_03247_));
 sky130_fd_sc_hd__mux4_2 _26506_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net429),
    .S1(net433),
    .X(_03248_));
 sky130_fd_sc_hd__mux4_2 _26507_ (.A0(_03245_),
    .A1(_03246_),
    .A2(_03247_),
    .A3(_03248_),
    .S0(net422),
    .S1(net421),
    .X(_03249_));
 sky130_fd_sc_hd__mux2i_4 _26508_ (.A0(_03244_),
    .A1(_03249_),
    .S(net419),
    .Y(_03250_));
 sky130_fd_sc_hd__xnor2_1 _26509_ (.A(_03239_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__xnor2_1 _26510_ (.A(_03086_),
    .B(_03251_),
    .Y(_11861_));
 sky130_fd_sc_hd__mux4_2 _26511_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net507),
    .S1(net512),
    .X(_03252_));
 sky130_fd_sc_hd__mux4_2 _26512_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net507),
    .S1(net512),
    .X(_03253_));
 sky130_fd_sc_hd__mux4_2 _26513_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net507),
    .S1(net512),
    .X(_03254_));
 sky130_fd_sc_hd__mux4_2 _26514_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net507),
    .S1(net512),
    .X(_03255_));
 sky130_fd_sc_hd__mux4_2 _26515_ (.A0(_03252_),
    .A1(_03253_),
    .A2(_03254_),
    .A3(_03255_),
    .S0(net503),
    .S1(net500),
    .X(_03256_));
 sky130_fd_sc_hd__mux4_2 _26516_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net509),
    .S1(net514),
    .X(_03257_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__mux4_2 _26518_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net509),
    .S1(net514),
    .X(_03259_));
 sky130_fd_sc_hd__mux4_2 _26519_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net509),
    .S1(net514),
    .X(_03260_));
 sky130_fd_sc_hd__mux4_2 _26520_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net509),
    .S1(net514),
    .X(_03261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_63 ();
 sky130_fd_sc_hd__mux4_2 _26522_ (.A0(_03257_),
    .A1(_03259_),
    .A2(_03260_),
    .A3(_03261_),
    .S0(net503),
    .S1(net500),
    .X(_03263_));
 sky130_fd_sc_hd__mux2i_4 _26523_ (.A0(_03256_),
    .A1(_03263_),
    .S(net497),
    .Y(_03264_));
 sky130_fd_sc_hd__mux4_2 _26524_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net506),
    .S1(net515),
    .X(_03265_));
 sky130_fd_sc_hd__mux4_2 _26525_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net506),
    .S1(net515),
    .X(_03266_));
 sky130_fd_sc_hd__mux4_2 _26526_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net506),
    .S1(net515),
    .X(_03267_));
 sky130_fd_sc_hd__mux4_2 _26527_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net506),
    .S1(net515),
    .X(_03268_));
 sky130_fd_sc_hd__mux4_2 _26528_ (.A0(_03265_),
    .A1(_03266_),
    .A2(_03267_),
    .A3(_03268_),
    .S0(net502),
    .S1(net499),
    .X(_03269_));
 sky130_fd_sc_hd__mux4_2 _26529_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net510),
    .S1(net514),
    .X(_03270_));
 sky130_fd_sc_hd__mux4_2 _26530_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net510),
    .S1(net514),
    .X(_03271_));
 sky130_fd_sc_hd__mux4_2 _26531_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net510),
    .S1(net514),
    .X(_03272_));
 sky130_fd_sc_hd__mux4_2 _26532_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net510),
    .S1(net514),
    .X(_03273_));
 sky130_fd_sc_hd__mux4_2 _26533_ (.A0(_03270_),
    .A1(_03271_),
    .A2(_03272_),
    .A3(_03273_),
    .S0(net503),
    .S1(net500),
    .X(_03274_));
 sky130_fd_sc_hd__mux2i_4 _26534_ (.A0(_03269_),
    .A1(_03274_),
    .S(net498),
    .Y(_03275_));
 sky130_fd_sc_hd__xnor2_1 _26535_ (.A(_03264_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__xnor2_2 _26536_ (.A(_02882_),
    .B(_03276_),
    .Y(_11860_));
 sky130_fd_sc_hd__mux4_2 _26537_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net543),
    .S1(net394),
    .X(_03277_));
 sky130_fd_sc_hd__mux4_2 _26538_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net543),
    .S1(net394),
    .X(_03278_));
 sky130_fd_sc_hd__mux4_2 _26539_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net543),
    .S1(net394),
    .X(_03279_));
 sky130_fd_sc_hd__mux4_2 _26540_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net543),
    .S1(net394),
    .X(_03280_));
 sky130_fd_sc_hd__mux4_2 _26541_ (.A0(_03277_),
    .A1(_03278_),
    .A2(_03279_),
    .A3(_03280_),
    .S0(\count7_2[3] ),
    .S1(net383),
    .X(_03281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__mux4_2 _26543_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net393),
    .S1(net394),
    .X(_03283_));
 sky130_fd_sc_hd__mux4_2 _26544_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net393),
    .S1(net394),
    .X(_03284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_61 ();
 sky130_fd_sc_hd__mux4_2 _26546_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net393),
    .S1(net394),
    .X(_03286_));
 sky130_fd_sc_hd__mux4_2 _26547_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net393),
    .S1(net394),
    .X(_03287_));
 sky130_fd_sc_hd__mux4_2 _26548_ (.A0(_03283_),
    .A1(_03284_),
    .A2(_03286_),
    .A3(_03287_),
    .S0(net386),
    .S1(net383),
    .X(_03288_));
 sky130_fd_sc_hd__mux2i_4 _26549_ (.A0(_03281_),
    .A1(_03288_),
    .S(\count7_2[5] ),
    .Y(_11859_));
 sky130_fd_sc_hd__mux4_2 _26550_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net465),
    .S1(net475),
    .X(_03289_));
 sky130_fd_sc_hd__mux4_2 _26551_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net465),
    .S1(net475),
    .X(_03290_));
 sky130_fd_sc_hd__mux4_2 _26552_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net465),
    .S1(net475),
    .X(_03291_));
 sky130_fd_sc_hd__mux4_2 _26553_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net465),
    .S1(net475),
    .X(_03292_));
 sky130_fd_sc_hd__mux4_2 _26554_ (.A0(_03289_),
    .A1(_03290_),
    .A2(_03291_),
    .A3(_03292_),
    .S0(net462),
    .S1(net460),
    .X(_03293_));
 sky130_fd_sc_hd__mux4_2 _26555_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net467),
    .S1(net476),
    .X(_03294_));
 sky130_fd_sc_hd__mux4_2 _26556_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net467),
    .S1(net476),
    .X(_03295_));
 sky130_fd_sc_hd__mux4_2 _26557_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net467),
    .S1(net476),
    .X(_03296_));
 sky130_fd_sc_hd__mux4_2 _26558_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net467),
    .S1(net476),
    .X(_03297_));
 sky130_fd_sc_hd__mux4_2 _26559_ (.A0(_03294_),
    .A1(_03295_),
    .A2(_03296_),
    .A3(_03297_),
    .S0(net463),
    .S1(net459),
    .X(_03298_));
 sky130_fd_sc_hd__mux2i_4 _26560_ (.A0(_03293_),
    .A1(_03298_),
    .S(net458),
    .Y(_11864_));
 sky130_fd_sc_hd__mux4_2 _26561_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net425),
    .S1(net436),
    .X(_03299_));
 sky130_fd_sc_hd__mux4_2 _26562_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net425),
    .S1(net436),
    .X(_03300_));
 sky130_fd_sc_hd__mux4_2 _26563_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net425),
    .S1(net436),
    .X(_03301_));
 sky130_fd_sc_hd__mux4_2 _26564_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net425),
    .S1(net436),
    .X(_03302_));
 sky130_fd_sc_hd__mux4_2 _26565_ (.A0(_03299_),
    .A1(_03300_),
    .A2(_03301_),
    .A3(_03302_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_03303_));
 sky130_fd_sc_hd__mux4_2 _26566_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net424),
    .S1(net435),
    .X(_03304_));
 sky130_fd_sc_hd__mux4_2 _26567_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net424),
    .S1(net435),
    .X(_03305_));
 sky130_fd_sc_hd__mux4_2 _26568_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net425),
    .S1(net435),
    .X(_03306_));
 sky130_fd_sc_hd__mux4_2 _26569_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net425),
    .S1(net435),
    .X(_03307_));
 sky130_fd_sc_hd__mux4_2 _26570_ (.A0(_03304_),
    .A1(_03305_),
    .A2(_03306_),
    .A3(_03307_),
    .S0(net549),
    .S1(net548),
    .X(_03308_));
 sky130_fd_sc_hd__mux2i_4 _26571_ (.A0(_03303_),
    .A1(_03308_),
    .S(\count2_2[5] ),
    .Y(_03309_));
 sky130_fd_sc_hd__mux4_2 _26572_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net425),
    .S1(net436),
    .X(_03310_));
 sky130_fd_sc_hd__mux4_2 _26573_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net425),
    .S1(net436),
    .X(_03311_));
 sky130_fd_sc_hd__mux4_2 _26574_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net425),
    .S1(net436),
    .X(_03312_));
 sky130_fd_sc_hd__mux4_2 _26575_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net425),
    .S1(net436),
    .X(_03313_));
 sky130_fd_sc_hd__mux4_2 _26576_ (.A0(_03310_),
    .A1(_03311_),
    .A2(_03312_),
    .A3(_03313_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_03314_));
 sky130_fd_sc_hd__mux4_2 _26577_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net424),
    .S1(net435),
    .X(_03315_));
 sky130_fd_sc_hd__mux4_2 _26578_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net424),
    .S1(net435),
    .X(_03316_));
 sky130_fd_sc_hd__mux4_2 _26579_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net424),
    .S1(net435),
    .X(_03317_));
 sky130_fd_sc_hd__mux4_2 _26580_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net424),
    .S1(net435),
    .X(_03318_));
 sky130_fd_sc_hd__mux4_2 _26581_ (.A0(_03315_),
    .A1(_03316_),
    .A2(_03317_),
    .A3(_03318_),
    .S0(net549),
    .S1(net548),
    .X(_03319_));
 sky130_fd_sc_hd__mux2i_4 _26582_ (.A0(_03314_),
    .A1(_03319_),
    .S(\count2_2[5] ),
    .Y(_03320_));
 sky130_fd_sc_hd__xnor2_1 _26583_ (.A(_03309_),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_1 _26584_ (.A(_03168_),
    .B(_03321_),
    .Y(_11869_));
 sky130_fd_sc_hd__mux4_2 _26585_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net506),
    .S1(net515),
    .X(_03322_));
 sky130_fd_sc_hd__mux4_2 _26586_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net506),
    .S1(net515),
    .X(_03323_));
 sky130_fd_sc_hd__mux4_2 _26587_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net506),
    .S1(net515),
    .X(_03324_));
 sky130_fd_sc_hd__mux4_2 _26588_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net506),
    .S1(net515),
    .X(_03325_));
 sky130_fd_sc_hd__mux4_2 _26589_ (.A0(_03322_),
    .A1(_03323_),
    .A2(_03324_),
    .A3(_03325_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_03326_));
 sky130_fd_sc_hd__mux4_2 _26590_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net511),
    .S1(net515),
    .X(_03327_));
 sky130_fd_sc_hd__mux4_2 _26591_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net511),
    .S1(net515),
    .X(_03328_));
 sky130_fd_sc_hd__mux4_2 _26592_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net511),
    .S1(net515),
    .X(_03329_));
 sky130_fd_sc_hd__mux4_2 _26593_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net511),
    .S1(net515),
    .X(_03330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_60 ();
 sky130_fd_sc_hd__mux4_2 _26595_ (.A0(_03327_),
    .A1(_03328_),
    .A2(_03329_),
    .A3(_03330_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_03332_));
 sky130_fd_sc_hd__mux2i_4 _26596_ (.A0(_03326_),
    .A1(_03332_),
    .S(net498),
    .Y(_03333_));
 sky130_fd_sc_hd__mux4_2 _26597_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net506),
    .S1(net515),
    .X(_03334_));
 sky130_fd_sc_hd__mux4_2 _26598_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net506),
    .S1(net515),
    .X(_03335_));
 sky130_fd_sc_hd__mux4_2 _26599_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net506),
    .S1(net515),
    .X(_03336_));
 sky130_fd_sc_hd__mux4_2 _26600_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net506),
    .S1(net515),
    .X(_03337_));
 sky130_fd_sc_hd__mux4_2 _26601_ (.A0(_03334_),
    .A1(_03335_),
    .A2(_03336_),
    .A3(_03337_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_03338_));
 sky130_fd_sc_hd__mux4_2 _26602_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net511),
    .S1(net515),
    .X(_03339_));
 sky130_fd_sc_hd__mux4_2 _26603_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net511),
    .S1(net516),
    .X(_03340_));
 sky130_fd_sc_hd__mux4_2 _26604_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net511),
    .S1(net516),
    .X(_03341_));
 sky130_fd_sc_hd__mux4_2 _26605_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net511),
    .S1(net516),
    .X(_03342_));
 sky130_fd_sc_hd__mux4_2 _26606_ (.A0(_03339_),
    .A1(_03340_),
    .A2(_03341_),
    .A3(_03342_),
    .S0(net503),
    .S1(\count15_2[4] ),
    .X(_03343_));
 sky130_fd_sc_hd__mux2i_4 _26607_ (.A0(_03338_),
    .A1(_03343_),
    .S(net498),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_1 _26608_ (.A(_03333_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__xnor2_1 _26609_ (.A(net1132),
    .B(_03345_),
    .Y(_11868_));
 sky130_fd_sc_hd__mux4_2 _26610_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net543),
    .S1(net394),
    .X(_03346_));
 sky130_fd_sc_hd__mux4_2 _26611_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net543),
    .S1(net394),
    .X(_03347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_59 ();
 sky130_fd_sc_hd__mux4_2 _26613_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net543),
    .S1(net394),
    .X(_03349_));
 sky130_fd_sc_hd__mux4_2 _26614_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net543),
    .S1(net394),
    .X(_03350_));
 sky130_fd_sc_hd__mux4_2 _26615_ (.A0(_03346_),
    .A1(_03347_),
    .A2(_03349_),
    .A3(_03350_),
    .S0(\count7_2[3] ),
    .S1(net383),
    .X(_03351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_58 ();
 sky130_fd_sc_hd__mux4_2 _26617_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net389),
    .S1(net394),
    .X(_03353_));
 sky130_fd_sc_hd__mux4_2 _26618_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net389),
    .S1(net394),
    .X(_03354_));
 sky130_fd_sc_hd__mux4_2 _26619_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net389),
    .S1(net394),
    .X(_03355_));
 sky130_fd_sc_hd__mux4_2 _26620_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net389),
    .S1(net394),
    .X(_03356_));
 sky130_fd_sc_hd__mux4_2 _26621_ (.A0(_03353_),
    .A1(_03354_),
    .A2(_03355_),
    .A3(_03356_),
    .S0(net386),
    .S1(net383),
    .X(_03357_));
 sky130_fd_sc_hd__mux2i_4 _26622_ (.A0(_03351_),
    .A1(_03357_),
    .S(net381),
    .Y(_11867_));
 sky130_fd_sc_hd__mux4_2 _26623_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03358_));
 sky130_fd_sc_hd__mux4_2 _26624_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03359_));
 sky130_fd_sc_hd__mux4_2 _26625_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03360_));
 sky130_fd_sc_hd__mux4_2 _26626_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03361_));
 sky130_fd_sc_hd__mux4_2 _26627_ (.A0(_03358_),
    .A1(_03359_),
    .A2(_03360_),
    .A3(_03361_),
    .S0(net464),
    .S1(net461),
    .X(_03362_));
 sky130_fd_sc_hd__mux4_2 _26628_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03363_));
 sky130_fd_sc_hd__mux4_2 _26629_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03364_));
 sky130_fd_sc_hd__mux4_2 _26630_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03365_));
 sky130_fd_sc_hd__mux4_2 _26631_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net468),
    .S1(net475),
    .X(_03366_));
 sky130_fd_sc_hd__mux4_2 _26632_ (.A0(_03363_),
    .A1(_03364_),
    .A2(_03365_),
    .A3(_03366_),
    .S0(net464),
    .S1(net461),
    .X(_03367_));
 sky130_fd_sc_hd__mux2i_4 _26633_ (.A0(_03362_),
    .A1(_03367_),
    .S(\count16_2[5] ),
    .Y(_11872_));
 sky130_fd_sc_hd__mux4_2 _26634_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net426),
    .S1(net431),
    .X(_03368_));
 sky130_fd_sc_hd__mux4_2 _26635_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net426),
    .S1(net431),
    .X(_03369_));
 sky130_fd_sc_hd__mux4_2 _26636_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net426),
    .S1(net431),
    .X(_03370_));
 sky130_fd_sc_hd__mux4_2 _26637_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net426),
    .S1(net431),
    .X(_03371_));
 sky130_fd_sc_hd__mux4_2 _26638_ (.A0(_03368_),
    .A1(_03369_),
    .A2(_03370_),
    .A3(_03371_),
    .S0(net423),
    .S1(net421),
    .X(_03372_));
 sky130_fd_sc_hd__mux4_2 _26639_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net429),
    .S1(net433),
    .X(_03373_));
 sky130_fd_sc_hd__mux4_2 _26640_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net429),
    .S1(net433),
    .X(_03374_));
 sky130_fd_sc_hd__mux4_2 _26641_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net429),
    .S1(net433),
    .X(_03375_));
 sky130_fd_sc_hd__mux4_2 _26642_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net429),
    .S1(net433),
    .X(_03376_));
 sky130_fd_sc_hd__mux4_2 _26643_ (.A0(_03373_),
    .A1(_03374_),
    .A2(_03375_),
    .A3(_03376_),
    .S0(net422),
    .S1(net420),
    .X(_03377_));
 sky130_fd_sc_hd__mux2i_4 _26644_ (.A0(_03372_),
    .A1(_03377_),
    .S(net418),
    .Y(_03378_));
 sky130_fd_sc_hd__mux4_2 _26645_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net427),
    .S1(net432),
    .X(_03379_));
 sky130_fd_sc_hd__mux4_2 _26646_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net427),
    .S1(net432),
    .X(_03380_));
 sky130_fd_sc_hd__mux4_2 _26647_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net427),
    .S1(net432),
    .X(_03381_));
 sky130_fd_sc_hd__mux4_2 _26648_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net427),
    .S1(net432),
    .X(_03382_));
 sky130_fd_sc_hd__mux4_2 _26649_ (.A0(_03379_),
    .A1(_03380_),
    .A2(_03381_),
    .A3(_03382_),
    .S0(net423),
    .S1(net421),
    .X(_03383_));
 sky130_fd_sc_hd__mux4_2 _26650_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net429),
    .S1(net433),
    .X(_03384_));
 sky130_fd_sc_hd__mux4_2 _26651_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net429),
    .S1(net433),
    .X(_03385_));
 sky130_fd_sc_hd__mux4_2 _26652_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net429),
    .S1(net433),
    .X(_03386_));
 sky130_fd_sc_hd__mux4_2 _26653_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net429),
    .S1(net433),
    .X(_03387_));
 sky130_fd_sc_hd__mux4_2 _26654_ (.A0(_03384_),
    .A1(_03385_),
    .A2(_03386_),
    .A3(_03387_),
    .S0(net422),
    .S1(net420),
    .X(_03388_));
 sky130_fd_sc_hd__mux2i_4 _26655_ (.A0(_03383_),
    .A1(_03388_),
    .S(net418),
    .Y(_03389_));
 sky130_fd_sc_hd__xnor2_1 _26656_ (.A(_03378_),
    .B(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__xnor2_1 _26657_ (.A(_03250_),
    .B(_03390_),
    .Y(_11877_));
 sky130_fd_sc_hd__mux4_2 _26658_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net506),
    .S1(net515),
    .X(_03391_));
 sky130_fd_sc_hd__mux4_2 _26659_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net506),
    .S1(net515),
    .X(_03392_));
 sky130_fd_sc_hd__mux4_2 _26660_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net506),
    .S1(net515),
    .X(_03393_));
 sky130_fd_sc_hd__mux4_2 _26661_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net506),
    .S1(net515),
    .X(_03394_));
 sky130_fd_sc_hd__mux4_2 _26662_ (.A0(_03391_),
    .A1(_03392_),
    .A2(_03393_),
    .A3(_03394_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_03395_));
 sky130_fd_sc_hd__mux4_2 _26663_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net511),
    .S1(net515),
    .X(_03396_));
 sky130_fd_sc_hd__mux4_2 _26664_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net511),
    .S1(net515),
    .X(_03397_));
 sky130_fd_sc_hd__mux4_2 _26665_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net511),
    .S1(net515),
    .X(_03398_));
 sky130_fd_sc_hd__mux4_2 _26666_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net511),
    .S1(net515),
    .X(_03399_));
 sky130_fd_sc_hd__mux4_2 _26667_ (.A0(_03396_),
    .A1(_03397_),
    .A2(_03398_),
    .A3(_03399_),
    .S0(net503),
    .S1(\count15_2[4] ),
    .X(_03400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_57 ();
 sky130_fd_sc_hd__mux2i_4 _26669_ (.A0(_03395_),
    .A1(_03400_),
    .S(net498),
    .Y(_03402_));
 sky130_fd_sc_hd__mux4_2 _26670_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03403_));
 sky130_fd_sc_hd__mux4_2 _26671_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03404_));
 sky130_fd_sc_hd__mux4_2 _26672_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03405_));
 sky130_fd_sc_hd__mux4_2 _26673_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03406_));
 sky130_fd_sc_hd__mux4_2 _26674_ (.A0(_03403_),
    .A1(_03404_),
    .A2(_03405_),
    .A3(_03406_),
    .S0(net502),
    .S1(net499),
    .X(_03407_));
 sky130_fd_sc_hd__mux4_2 _26675_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03408_));
 sky130_fd_sc_hd__mux4_2 _26676_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03409_));
 sky130_fd_sc_hd__mux4_2 _26677_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03410_));
 sky130_fd_sc_hd__mux4_2 _26678_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net508),
    .S1(net513),
    .X(_03411_));
 sky130_fd_sc_hd__mux4_2 _26679_ (.A0(_03408_),
    .A1(_03409_),
    .A2(_03410_),
    .A3(_03411_),
    .S0(net502),
    .S1(net499),
    .X(_03412_));
 sky130_fd_sc_hd__mux2i_4 _26680_ (.A0(_03407_),
    .A1(_03412_),
    .S(net497),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_1 _26681_ (.A(_03402_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_1 _26682_ (.A(net1130),
    .B(_03414_),
    .Y(_11876_));
 sky130_fd_sc_hd__mux4_2 _26683_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net543),
    .S1(\count7_2[1] ),
    .X(_03415_));
 sky130_fd_sc_hd__mux4_2 _26684_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net543),
    .S1(\count7_2[1] ),
    .X(_03416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_56 ();
 sky130_fd_sc_hd__mux4_2 _26686_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net543),
    .S1(\count7_2[1] ),
    .X(_03418_));
 sky130_fd_sc_hd__mux4_2 _26687_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net543),
    .S1(net394),
    .X(_03419_));
 sky130_fd_sc_hd__mux4_2 _26688_ (.A0(_03415_),
    .A1(_03416_),
    .A2(_03418_),
    .A3(_03419_),
    .S0(\count7_2[3] ),
    .S1(net383),
    .X(_03420_));
 sky130_fd_sc_hd__mux4_2 _26689_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net393),
    .S1(net544),
    .X(_03421_));
 sky130_fd_sc_hd__mux4_2 _26690_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net393),
    .S1(net544),
    .X(_03422_));
 sky130_fd_sc_hd__mux4_2 _26691_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net393),
    .S1(net544),
    .X(_03423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_55 ();
 sky130_fd_sc_hd__mux4_2 _26693_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net393),
    .S1(net544),
    .X(_03425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_54 ();
 sky130_fd_sc_hd__mux4_2 _26695_ (.A0(_03421_),
    .A1(_03422_),
    .A2(_03423_),
    .A3(_03425_),
    .S0(net386),
    .S1(net383),
    .X(_03427_));
 sky130_fd_sc_hd__mux2i_4 _26696_ (.A0(_03420_),
    .A1(_03427_),
    .S(net381),
    .Y(_11875_));
 sky130_fd_sc_hd__mux4_2 _26697_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03428_));
 sky130_fd_sc_hd__mux4_2 _26698_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03429_));
 sky130_fd_sc_hd__mux4_2 _26699_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03430_));
 sky130_fd_sc_hd__mux4_2 _26700_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03431_));
 sky130_fd_sc_hd__mux4_2 _26701_ (.A0(_03428_),
    .A1(_03429_),
    .A2(_03430_),
    .A3(_03431_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_03432_));
 sky130_fd_sc_hd__mux4_2 _26702_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_03433_));
 sky130_fd_sc_hd__mux4_2 _26703_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_03434_));
 sky130_fd_sc_hd__mux4_2 _26704_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_03435_));
 sky130_fd_sc_hd__mux4_2 _26705_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(\count16_2[2] ),
    .S1(net477),
    .X(_03436_));
 sky130_fd_sc_hd__mux4_2 _26706_ (.A0(_03433_),
    .A1(_03434_),
    .A2(_03435_),
    .A3(_03436_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_03437_));
 sky130_fd_sc_hd__mux2i_2 _26707_ (.A0(_03432_),
    .A1(_03437_),
    .S(\count16_2[5] ),
    .Y(_11880_));
 sky130_fd_sc_hd__mux4_2 _26708_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net425),
    .S1(net436),
    .X(_03438_));
 sky130_fd_sc_hd__mux4_2 _26709_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net425),
    .S1(net436),
    .X(_03439_));
 sky130_fd_sc_hd__mux4_2 _26710_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net425),
    .S1(net436),
    .X(_03440_));
 sky130_fd_sc_hd__mux4_2 _26711_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net425),
    .S1(net436),
    .X(_03441_));
 sky130_fd_sc_hd__mux4_2 _26712_ (.A0(_03438_),
    .A1(_03439_),
    .A2(_03440_),
    .A3(_03441_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_03442_));
 sky130_fd_sc_hd__mux4_2 _26713_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net429),
    .S1(net433),
    .X(_03443_));
 sky130_fd_sc_hd__mux4_2 _26714_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net430),
    .S1(net433),
    .X(_03444_));
 sky130_fd_sc_hd__mux4_2 _26715_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net430),
    .S1(net433),
    .X(_03445_));
 sky130_fd_sc_hd__mux4_2 _26716_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net430),
    .S1(net433),
    .X(_03446_));
 sky130_fd_sc_hd__mux4_2 _26717_ (.A0(_03443_),
    .A1(_03444_),
    .A2(_03445_),
    .A3(_03446_),
    .S0(net423),
    .S1(net548),
    .X(_03447_));
 sky130_fd_sc_hd__mux2i_4 _26718_ (.A0(_03442_),
    .A1(_03447_),
    .S(net419),
    .Y(_03448_));
 sky130_fd_sc_hd__xnor2_1 _26719_ (.A(_03320_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__xnor2_2 _26720_ (.A(_02788_),
    .B(_03449_),
    .Y(_11885_));
 sky130_fd_sc_hd__mux4_2 _26721_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net506),
    .S1(net515),
    .X(_03450_));
 sky130_fd_sc_hd__mux4_2 _26722_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net506),
    .S1(net515),
    .X(_03451_));
 sky130_fd_sc_hd__mux4_2 _26723_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net506),
    .S1(net515),
    .X(_03452_));
 sky130_fd_sc_hd__mux4_2 _26724_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net506),
    .S1(net515),
    .X(_03453_));
 sky130_fd_sc_hd__mux4_2 _26725_ (.A0(_03450_),
    .A1(_03451_),
    .A2(_03452_),
    .A3(_03453_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_03454_));
 sky130_fd_sc_hd__mux4_2 _26726_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net510),
    .S1(net514),
    .X(_03455_));
 sky130_fd_sc_hd__mux4_2 _26727_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net510),
    .S1(net516),
    .X(_03456_));
 sky130_fd_sc_hd__mux4_2 _26728_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net510),
    .S1(net516),
    .X(_03457_));
 sky130_fd_sc_hd__mux4_2 _26729_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net510),
    .S1(net516),
    .X(_03458_));
 sky130_fd_sc_hd__mux4_2 _26730_ (.A0(_03455_),
    .A1(_03456_),
    .A2(_03457_),
    .A3(_03458_),
    .S0(net503),
    .S1(net500),
    .X(_03459_));
 sky130_fd_sc_hd__mux2i_4 _26731_ (.A0(_03454_),
    .A1(_03459_),
    .S(net497),
    .Y(_03460_));
 sky130_fd_sc_hd__mux4_2 _26732_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03461_));
 sky130_fd_sc_hd__mux4_2 _26733_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03462_));
 sky130_fd_sc_hd__mux4_2 _26734_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03463_));
 sky130_fd_sc_hd__mux4_2 _26735_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03464_));
 sky130_fd_sc_hd__mux4_2 _26736_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(net502),
    .S1(net499),
    .X(_03465_));
 sky130_fd_sc_hd__mux4_2 _26737_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03466_));
 sky130_fd_sc_hd__mux4_2 _26738_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03467_));
 sky130_fd_sc_hd__mux4_2 _26739_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03468_));
 sky130_fd_sc_hd__mux4_2 _26740_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net508),
    .S1(net513),
    .X(_03469_));
 sky130_fd_sc_hd__mux4_2 _26741_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(net502),
    .S1(net499),
    .X(_03470_));
 sky130_fd_sc_hd__mux2i_4 _26742_ (.A0(_03465_),
    .A1(_03470_),
    .S(net497),
    .Y(_03471_));
 sky130_fd_sc_hd__xnor2_1 _26743_ (.A(_03460_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__xnor2_1 _26744_ (.A(_03205_),
    .B(_03472_),
    .Y(_11884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_53 ();
 sky130_fd_sc_hd__mux4_2 _26746_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net388),
    .S1(net398),
    .X(_03474_));
 sky130_fd_sc_hd__mux4_2 _26747_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net388),
    .S1(net398),
    .X(_03475_));
 sky130_fd_sc_hd__mux4_2 _26748_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net388),
    .S1(net398),
    .X(_03476_));
 sky130_fd_sc_hd__mux4_2 _26749_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net388),
    .S1(net398),
    .X(_03477_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_52 ();
 sky130_fd_sc_hd__mux4_2 _26751_ (.A0(_03474_),
    .A1(_03475_),
    .A2(_03476_),
    .A3(_03477_),
    .S0(net386),
    .S1(net383),
    .X(_03479_));
 sky130_fd_sc_hd__mux4_2 _26752_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net392),
    .S1(net544),
    .X(_03480_));
 sky130_fd_sc_hd__mux4_2 _26753_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net392),
    .S1(net544),
    .X(_03481_));
 sky130_fd_sc_hd__mux4_2 _26754_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net392),
    .S1(net544),
    .X(_03482_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_51 ();
 sky130_fd_sc_hd__mux4_2 _26756_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net392),
    .S1(net544),
    .X(_03484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_50 ();
 sky130_fd_sc_hd__mux4_2 _26758_ (.A0(_03480_),
    .A1(_03481_),
    .A2(_03482_),
    .A3(_03484_),
    .S0(net385),
    .S1(\count7_2[4] ),
    .X(_03486_));
 sky130_fd_sc_hd__mux2i_4 _26759_ (.A0(_03479_),
    .A1(_03486_),
    .S(net381),
    .Y(_11883_));
 sky130_fd_sc_hd__mux4_2 _26760_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03487_));
 sky130_fd_sc_hd__mux4_2 _26761_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03488_));
 sky130_fd_sc_hd__mux4_2 _26762_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03489_));
 sky130_fd_sc_hd__mux4_2 _26763_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(\count16_2[2] ),
    .S1(net553),
    .X(_03490_));
 sky130_fd_sc_hd__mux4_2 _26764_ (.A0(_03487_),
    .A1(_03488_),
    .A2(_03489_),
    .A3(_03490_),
    .S0(net464),
    .S1(\count16_2[4] ),
    .X(_03491_));
 sky130_fd_sc_hd__mux4_2 _26765_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net471),
    .S1(net477),
    .X(_03492_));
 sky130_fd_sc_hd__mux4_2 _26766_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net471),
    .S1(net477),
    .X(_03493_));
 sky130_fd_sc_hd__mux4_2 _26767_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net471),
    .S1(net477),
    .X(_03494_));
 sky130_fd_sc_hd__mux4_2 _26768_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net471),
    .S1(net477),
    .X(_03495_));
 sky130_fd_sc_hd__mux4_2 _26769_ (.A0(_03492_),
    .A1(_03493_),
    .A2(_03494_),
    .A3(_03495_),
    .S0(net463),
    .S1(net461),
    .X(_03496_));
 sky130_fd_sc_hd__mux2i_2 _26770_ (.A0(_03491_),
    .A1(_03496_),
    .S(net458),
    .Y(_11888_));
 sky130_fd_sc_hd__mux4_2 _26771_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net426),
    .S1(net431),
    .X(_03497_));
 sky130_fd_sc_hd__mux4_2 _26772_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net426),
    .S1(net431),
    .X(_03498_));
 sky130_fd_sc_hd__mux4_2 _26773_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net426),
    .S1(net431),
    .X(_03499_));
 sky130_fd_sc_hd__mux4_2 _26774_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net426),
    .S1(net431),
    .X(_03500_));
 sky130_fd_sc_hd__mux4_2 _26775_ (.A0(_03497_),
    .A1(_03498_),
    .A2(_03499_),
    .A3(_03500_),
    .S0(net423),
    .S1(net421),
    .X(_03501_));
 sky130_fd_sc_hd__mux4_2 _26776_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net429),
    .S1(net432),
    .X(_03502_));
 sky130_fd_sc_hd__mux4_2 _26777_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net429),
    .S1(net432),
    .X(_03503_));
 sky130_fd_sc_hd__mux4_2 _26778_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net429),
    .S1(net432),
    .X(_03504_));
 sky130_fd_sc_hd__mux4_2 _26779_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net429),
    .S1(net433),
    .X(_03505_));
 sky130_fd_sc_hd__mux4_2 _26780_ (.A0(_03502_),
    .A1(_03503_),
    .A2(_03504_),
    .A3(_03505_),
    .S0(net423),
    .S1(net421),
    .X(_03506_));
 sky130_fd_sc_hd__mux2i_4 _26781_ (.A0(_03501_),
    .A1(_03506_),
    .S(net419),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_1 _26782_ (.A(_03389_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__xnor2_1 _26783_ (.A(_02964_),
    .B(_03508_),
    .Y(_11893_));
 sky130_fd_sc_hd__mux4_2 _26784_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net505),
    .S1(net517),
    .X(_03509_));
 sky130_fd_sc_hd__mux4_2 _26785_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net505),
    .S1(net517),
    .X(_03510_));
 sky130_fd_sc_hd__mux4_2 _26786_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03511_));
 sky130_fd_sc_hd__mux4_2 _26787_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03512_));
 sky130_fd_sc_hd__mux4_2 _26788_ (.A0(_03509_),
    .A1(_03510_),
    .A2(_03511_),
    .A3(_03512_),
    .S0(net504),
    .S1(net501),
    .X(_03513_));
 sky130_fd_sc_hd__mux4_2 _26789_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03514_));
 sky130_fd_sc_hd__mux4_2 _26790_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03515_));
 sky130_fd_sc_hd__mux4_2 _26791_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03516_));
 sky130_fd_sc_hd__mux4_2 _26792_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03517_));
 sky130_fd_sc_hd__mux4_2 _26793_ (.A0(_03514_),
    .A1(_03515_),
    .A2(_03516_),
    .A3(_03517_),
    .S0(net504),
    .S1(net501),
    .X(_03518_));
 sky130_fd_sc_hd__mux2i_4 _26794_ (.A0(_03513_),
    .A1(_03518_),
    .S(\count15_2[5] ),
    .Y(_03519_));
 sky130_fd_sc_hd__mux4_2 _26795_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03520_));
 sky130_fd_sc_hd__mux4_2 _26796_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03521_));
 sky130_fd_sc_hd__mux4_2 _26797_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03522_));
 sky130_fd_sc_hd__mux4_2 _26798_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03523_));
 sky130_fd_sc_hd__mux4_2 _26799_ (.A0(_03520_),
    .A1(_03521_),
    .A2(_03522_),
    .A3(_03523_),
    .S0(net502),
    .S1(net499),
    .X(_03524_));
 sky130_fd_sc_hd__mux4_2 _26800_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03525_));
 sky130_fd_sc_hd__mux4_2 _26801_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03526_));
 sky130_fd_sc_hd__mux4_2 _26802_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03527_));
 sky130_fd_sc_hd__mux4_2 _26803_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net508),
    .S1(net513),
    .X(_03528_));
 sky130_fd_sc_hd__mux4_2 _26804_ (.A0(_03525_),
    .A1(_03526_),
    .A2(_03527_),
    .A3(_03528_),
    .S0(net502),
    .S1(net499),
    .X(_03529_));
 sky130_fd_sc_hd__mux2i_4 _26805_ (.A0(_03524_),
    .A1(_03529_),
    .S(net497),
    .Y(_03530_));
 sky130_fd_sc_hd__xnor2_1 _26806_ (.A(_03519_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__xnor2_1 _26807_ (.A(_03275_),
    .B(_03531_),
    .Y(_11892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_49 ();
 sky130_fd_sc_hd__mux4_2 _26809_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net390),
    .S1(net396),
    .X(_03533_));
 sky130_fd_sc_hd__mux4_2 _26810_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net390),
    .S1(net396),
    .X(_03534_));
 sky130_fd_sc_hd__mux4_2 _26811_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net390),
    .S1(net396),
    .X(_03535_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_48 ();
 sky130_fd_sc_hd__mux4_2 _26813_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net390),
    .S1(net396),
    .X(_03537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__mux4_2 _26815_ (.A0(_03533_),
    .A1(_03534_),
    .A2(_03535_),
    .A3(_03537_),
    .S0(net384),
    .S1(net542),
    .X(_03539_));
 sky130_fd_sc_hd__mux4_2 _26816_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net390),
    .S1(net395),
    .X(_03540_));
 sky130_fd_sc_hd__mux4_2 _26817_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net390),
    .S1(net395),
    .X(_03541_));
 sky130_fd_sc_hd__mux4_2 _26818_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net390),
    .S1(net395),
    .X(_03542_));
 sky130_fd_sc_hd__mux4_2 _26819_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net390),
    .S1(net395),
    .X(_03543_));
 sky130_fd_sc_hd__mux4_2 _26820_ (.A0(_03540_),
    .A1(_03541_),
    .A2(_03542_),
    .A3(_03543_),
    .S0(net385),
    .S1(net382),
    .X(_03544_));
 sky130_fd_sc_hd__mux2i_4 _26821_ (.A0(_03539_),
    .A1(_03544_),
    .S(net380),
    .Y(_11891_));
 sky130_fd_sc_hd__mux4_2 _26822_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net466),
    .S1(net474),
    .X(_03545_));
 sky130_fd_sc_hd__mux4_2 _26823_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net466),
    .S1(net474),
    .X(_03546_));
 sky130_fd_sc_hd__mux4_2 _26824_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net466),
    .S1(net474),
    .X(_03547_));
 sky130_fd_sc_hd__mux4_2 _26825_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net466),
    .S1(net474),
    .X(_03548_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_46 ();
 sky130_fd_sc_hd__mux4_2 _26827_ (.A0(_03545_),
    .A1(_03546_),
    .A2(_03547_),
    .A3(_03548_),
    .S0(net462),
    .S1(net460),
    .X(_03550_));
 sky130_fd_sc_hd__mux4_2 _26828_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net469),
    .S1(net473),
    .X(_03551_));
 sky130_fd_sc_hd__mux4_2 _26829_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net469),
    .S1(net473),
    .X(_03552_));
 sky130_fd_sc_hd__mux4_2 _26830_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net469),
    .S1(net473),
    .X(_03553_));
 sky130_fd_sc_hd__mux4_2 _26831_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net469),
    .S1(net473),
    .X(_03554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_45 ();
 sky130_fd_sc_hd__mux4_2 _26833_ (.A0(_03551_),
    .A1(_03552_),
    .A2(_03553_),
    .A3(_03554_),
    .S0(net463),
    .S1(net460),
    .X(_03556_));
 sky130_fd_sc_hd__mux2i_4 _26834_ (.A0(_03550_),
    .A1(_03556_),
    .S(net457),
    .Y(_11896_));
 sky130_fd_sc_hd__mux4_2 _26835_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net425),
    .S1(net436),
    .X(_03557_));
 sky130_fd_sc_hd__mux4_2 _26836_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net425),
    .S1(net436),
    .X(_03558_));
 sky130_fd_sc_hd__mux4_2 _26837_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net425),
    .S1(net436),
    .X(_03559_));
 sky130_fd_sc_hd__mux4_2 _26838_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net425),
    .S1(net436),
    .X(_03560_));
 sky130_fd_sc_hd__mux4_2 _26839_ (.A0(_03557_),
    .A1(_03558_),
    .A2(_03559_),
    .A3(_03560_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_03561_));
 sky130_fd_sc_hd__mux4_2 _26840_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net424),
    .S1(net435),
    .X(_03562_));
 sky130_fd_sc_hd__mux4_2 _26841_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net424),
    .S1(net435),
    .X(_03563_));
 sky130_fd_sc_hd__mux4_2 _26842_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net424),
    .S1(net435),
    .X(_03564_));
 sky130_fd_sc_hd__mux4_2 _26843_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net424),
    .S1(net435),
    .X(_03565_));
 sky130_fd_sc_hd__mux4_2 _26844_ (.A0(_03562_),
    .A1(_03563_),
    .A2(_03564_),
    .A3(_03565_),
    .S0(net549),
    .S1(net548),
    .X(_03566_));
 sky130_fd_sc_hd__mux2i_4 _26845_ (.A0(_03561_),
    .A1(_03566_),
    .S(\count2_2[5] ),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_1 _26846_ (.A(_03448_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__xnor2_2 _26847_ (.A(_02770_),
    .B(_03568_),
    .Y(_11901_));
 sky130_fd_sc_hd__mux4_2 _26848_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03569_));
 sky130_fd_sc_hd__mux4_2 _26849_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03570_));
 sky130_fd_sc_hd__mux4_2 _26850_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03571_));
 sky130_fd_sc_hd__mux4_2 _26851_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net557),
    .S1(\count15_2[1] ),
    .X(_03572_));
 sky130_fd_sc_hd__mux4_2 _26852_ (.A0(_03569_),
    .A1(_03570_),
    .A2(_03571_),
    .A3(_03572_),
    .S0(net504),
    .S1(net501),
    .X(_03573_));
 sky130_fd_sc_hd__mux4_2 _26853_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net511),
    .S1(net516),
    .X(_03574_));
 sky130_fd_sc_hd__mux4_2 _26854_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net511),
    .S1(net516),
    .X(_03575_));
 sky130_fd_sc_hd__mux4_2 _26855_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net511),
    .S1(net516),
    .X(_03576_));
 sky130_fd_sc_hd__mux4_2 _26856_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net511),
    .S1(net516),
    .X(_03577_));
 sky130_fd_sc_hd__mux4_2 _26857_ (.A0(_03574_),
    .A1(_03575_),
    .A2(_03576_),
    .A3(_03577_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03578_));
 sky130_fd_sc_hd__mux2i_4 _26858_ (.A0(_03573_),
    .A1(_03578_),
    .S(net498),
    .Y(_03579_));
 sky130_fd_sc_hd__mux4_2 _26859_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03580_));
 sky130_fd_sc_hd__mux4_2 _26860_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03581_));
 sky130_fd_sc_hd__mux4_2 _26861_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03582_));
 sky130_fd_sc_hd__mux4_2 _26862_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03583_));
 sky130_fd_sc_hd__mux4_2 _26863_ (.A0(_03580_),
    .A1(_03581_),
    .A2(_03582_),
    .A3(_03583_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_03584_));
 sky130_fd_sc_hd__mux4_2 _26864_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03585_));
 sky130_fd_sc_hd__mux4_2 _26865_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03586_));
 sky130_fd_sc_hd__mux4_2 _26866_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03587_));
 sky130_fd_sc_hd__mux4_2 _26867_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net506),
    .S1(net515),
    .X(_03588_));
 sky130_fd_sc_hd__mux4_2 _26868_ (.A0(_03585_),
    .A1(_03586_),
    .A2(_03587_),
    .A3(_03588_),
    .S0(net504),
    .S1(\count15_2[4] ),
    .X(_03589_));
 sky130_fd_sc_hd__mux2i_4 _26869_ (.A0(_03584_),
    .A1(_03589_),
    .S(net498),
    .Y(_03590_));
 sky130_fd_sc_hd__xnor2_1 _26870_ (.A(_03579_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__xnor2_1 _26871_ (.A(_03344_),
    .B(_03591_),
    .Y(_11900_));
 sky130_fd_sc_hd__mux4_2 _26872_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03592_));
 sky130_fd_sc_hd__mux4_2 _26873_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03593_));
 sky130_fd_sc_hd__mux4_2 _26874_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03594_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_44 ();
 sky130_fd_sc_hd__mux4_2 _26876_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03596_));
 sky130_fd_sc_hd__mux4_2 _26877_ (.A0(_03592_),
    .A1(_03593_),
    .A2(_03594_),
    .A3(_03596_),
    .S0(net384),
    .S1(net542),
    .X(_03597_));
 sky130_fd_sc_hd__mux4_2 _26878_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03598_));
 sky130_fd_sc_hd__mux4_2 _26879_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03599_));
 sky130_fd_sc_hd__mux4_2 _26880_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03600_));
 sky130_fd_sc_hd__mux4_2 _26881_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net390),
    .S1(net395),
    .X(_03601_));
 sky130_fd_sc_hd__mux4_2 _26882_ (.A0(_03598_),
    .A1(_03599_),
    .A2(_03600_),
    .A3(_03601_),
    .S0(net384),
    .S1(net542),
    .X(_03602_));
 sky130_fd_sc_hd__mux2i_4 _26883_ (.A0(_03597_),
    .A1(_03602_),
    .S(net380),
    .Y(_11899_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__mux4_2 _26885_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03604_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__mux4_2 _26887_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_41 ();
 sky130_fd_sc_hd__mux4_2 _26889_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03608_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_40 ();
 sky130_fd_sc_hd__mux4_2 _26891_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__mux4_2 _26893_ (.A0(_03604_),
    .A1(_03606_),
    .A2(_03608_),
    .A3(_03610_),
    .S0(\count16_2[3] ),
    .S1(net461),
    .X(_03612_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__mux4_2 _26895_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__mux4_2 _26897_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__mux4_2 _26899_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03618_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__mux4_2 _26901_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net472),
    .S1(net477),
    .X(_03620_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__mux4_2 _26903_ (.A0(_03614_),
    .A1(_03616_),
    .A2(_03618_),
    .A3(_03620_),
    .S0(\count16_2[3] ),
    .S1(net461),
    .X(_03622_));
 sky130_fd_sc_hd__mux2i_2 _26904_ (.A0(_03612_),
    .A1(_03622_),
    .S(net458),
    .Y(_11904_));
 sky130_fd_sc_hd__mux4_2 _26905_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net425),
    .S1(net436),
    .X(_03623_));
 sky130_fd_sc_hd__mux4_2 _26906_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net425),
    .S1(net436),
    .X(_03624_));
 sky130_fd_sc_hd__mux4_2 _26907_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net425),
    .S1(net436),
    .X(_03625_));
 sky130_fd_sc_hd__mux4_2 _26908_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net425),
    .S1(net436),
    .X(_03626_));
 sky130_fd_sc_hd__mux4_2 _26909_ (.A0(_03623_),
    .A1(_03624_),
    .A2(_03625_),
    .A3(_03626_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_03627_));
 sky130_fd_sc_hd__mux4_2 _26910_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net424),
    .S1(net435),
    .X(_03628_));
 sky130_fd_sc_hd__mux4_2 _26911_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net424),
    .S1(net435),
    .X(_03629_));
 sky130_fd_sc_hd__mux4_2 _26912_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net424),
    .S1(net435),
    .X(_03630_));
 sky130_fd_sc_hd__mux4_2 _26913_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net424),
    .S1(net435),
    .X(_03631_));
 sky130_fd_sc_hd__mux4_2 _26914_ (.A0(_03628_),
    .A1(_03629_),
    .A2(_03630_),
    .A3(_03631_),
    .S0(net549),
    .S1(net548),
    .X(_03632_));
 sky130_fd_sc_hd__mux2i_4 _26915_ (.A0(_03627_),
    .A1(_03632_),
    .S(\count2_2[5] ),
    .Y(_03633_));
 sky130_fd_sc_hd__xnor2_1 _26916_ (.A(_03507_),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__xnor2_2 _26917_ (.A(_02953_),
    .B(_03634_),
    .Y(_11909_));
 sky130_fd_sc_hd__mux4_2 _26918_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net506),
    .S1(net515),
    .X(_03635_));
 sky130_fd_sc_hd__mux4_2 _26919_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net506),
    .S1(net515),
    .X(_03636_));
 sky130_fd_sc_hd__mux4_2 _26920_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net506),
    .S1(net515),
    .X(_03637_));
 sky130_fd_sc_hd__mux4_2 _26921_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net506),
    .S1(net515),
    .X(_03638_));
 sky130_fd_sc_hd__mux4_2 _26922_ (.A0(_03635_),
    .A1(_03636_),
    .A2(_03637_),
    .A3(_03638_),
    .S0(net502),
    .S1(net499),
    .X(_03639_));
 sky130_fd_sc_hd__mux4_2 _26923_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net510),
    .S1(net514),
    .X(_03640_));
 sky130_fd_sc_hd__mux4_2 _26924_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net509),
    .S1(net514),
    .X(_03641_));
 sky130_fd_sc_hd__mux4_2 _26925_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net509),
    .S1(net514),
    .X(_03642_));
 sky130_fd_sc_hd__mux4_2 _26926_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net509),
    .S1(net514),
    .X(_03643_));
 sky130_fd_sc_hd__mux4_2 _26927_ (.A0(_03640_),
    .A1(_03641_),
    .A2(_03642_),
    .A3(_03643_),
    .S0(net503),
    .S1(net500),
    .X(_03644_));
 sky130_fd_sc_hd__mux2i_4 _26928_ (.A0(_03639_),
    .A1(_03644_),
    .S(net497),
    .Y(_03645_));
 sky130_fd_sc_hd__mux4_2 _26929_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03646_));
 sky130_fd_sc_hd__mux4_2 _26930_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03647_));
 sky130_fd_sc_hd__mux4_2 _26931_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03648_));
 sky130_fd_sc_hd__mux4_2 _26932_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03649_));
 sky130_fd_sc_hd__mux4_2 _26933_ (.A0(_03646_),
    .A1(_03647_),
    .A2(_03648_),
    .A3(_03649_),
    .S0(net502),
    .S1(net499),
    .X(_03650_));
 sky130_fd_sc_hd__mux4_2 _26934_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03651_));
 sky130_fd_sc_hd__mux4_2 _26935_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03652_));
 sky130_fd_sc_hd__mux4_2 _26936_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03653_));
 sky130_fd_sc_hd__mux4_2 _26937_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net510),
    .S1(net516),
    .X(_03654_));
 sky130_fd_sc_hd__mux4_2 _26938_ (.A0(_03651_),
    .A1(_03652_),
    .A2(_03653_),
    .A3(_03654_),
    .S0(net502),
    .S1(net499),
    .X(_03655_));
 sky130_fd_sc_hd__mux2i_4 _26939_ (.A0(_03650_),
    .A1(_03655_),
    .S(net497),
    .Y(_03656_));
 sky130_fd_sc_hd__xnor2_1 _26940_ (.A(_03645_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__xnor2_1 _26941_ (.A(_03402_),
    .B(_03657_),
    .Y(_11908_));
 sky130_fd_sc_hd__mux4_2 _26942_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net390),
    .S1(net395),
    .X(_03658_));
 sky130_fd_sc_hd__mux4_2 _26943_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net390),
    .S1(net395),
    .X(_03659_));
 sky130_fd_sc_hd__mux4_2 _26944_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net390),
    .S1(net395),
    .X(_03660_));
 sky130_fd_sc_hd__mux4_2 _26945_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net390),
    .S1(net395),
    .X(_03661_));
 sky130_fd_sc_hd__mux4_2 _26946_ (.A0(_03658_),
    .A1(_03659_),
    .A2(_03660_),
    .A3(_03661_),
    .S0(net384),
    .S1(net542),
    .X(_03662_));
 sky130_fd_sc_hd__mux4_2 _26947_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net391),
    .S1(net397),
    .X(_03663_));
 sky130_fd_sc_hd__mux4_2 _26948_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net391),
    .S1(net397),
    .X(_03664_));
 sky130_fd_sc_hd__mux4_2 _26949_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net391),
    .S1(net397),
    .X(_03665_));
 sky130_fd_sc_hd__mux4_2 _26950_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net391),
    .S1(net397),
    .X(_03666_));
 sky130_fd_sc_hd__mux4_2 _26951_ (.A0(_03663_),
    .A1(_03664_),
    .A2(_03665_),
    .A3(_03666_),
    .S0(net384),
    .S1(net542),
    .X(_03667_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__mux2i_4 _26953_ (.A0(_03662_),
    .A1(_03667_),
    .S(net380),
    .Y(_11907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__mux4_2 _26955_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net470),
    .S1(net473),
    .X(_03670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__mux4_2 _26957_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net470),
    .S1(net473),
    .X(_03672_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__mux4_2 _26959_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net470),
    .S1(net473),
    .X(_03674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__mux4_2 _26961_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net470),
    .S1(net473),
    .X(_03676_));
 sky130_fd_sc_hd__mux4_2 _26962_ (.A0(_03670_),
    .A1(_03672_),
    .A2(_03674_),
    .A3(_03676_),
    .S0(\count16_2[3] ),
    .S1(net459),
    .X(_03677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__mux4_2 _26964_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net470),
    .S1(net477),
    .X(_03679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__mux4_2 _26966_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net470),
    .S1(net477),
    .X(_03681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__mux4_2 _26968_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net470),
    .S1(net477),
    .X(_03683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__mux4_2 _26970_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net470),
    .S1(net477),
    .X(_03685_));
 sky130_fd_sc_hd__mux4_2 _26971_ (.A0(_03679_),
    .A1(_03681_),
    .A2(_03683_),
    .A3(_03685_),
    .S0(\count16_2[3] ),
    .S1(net460),
    .X(_03686_));
 sky130_fd_sc_hd__mux2i_4 _26972_ (.A0(_03677_),
    .A1(_03686_),
    .S(net457),
    .Y(_11912_));
 sky130_fd_sc_hd__mux4_2 _26973_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_03687_));
 sky130_fd_sc_hd__mux4_2 _26974_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_03688_));
 sky130_fd_sc_hd__mux4_2 _26975_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_03689_));
 sky130_fd_sc_hd__mux4_2 _26976_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(\count2_2[2] ),
    .S1(net436),
    .X(_03690_));
 sky130_fd_sc_hd__mux4_2 _26977_ (.A0(_03687_),
    .A1(_03688_),
    .A2(_03689_),
    .A3(_03690_),
    .S0(\count2_2[3] ),
    .S1(net548),
    .X(_03691_));
 sky130_fd_sc_hd__mux4_2 _26978_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_03692_));
 sky130_fd_sc_hd__mux4_2 _26979_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_03693_));
 sky130_fd_sc_hd__mux4_2 _26980_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_03694_));
 sky130_fd_sc_hd__mux4_2 _26981_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net430),
    .S1(\count2_2[1] ),
    .X(_03695_));
 sky130_fd_sc_hd__mux4_2 _26982_ (.A0(_03692_),
    .A1(_03693_),
    .A2(_03694_),
    .A3(_03695_),
    .S0(net423),
    .S1(\count2_2[4] ),
    .X(_03696_));
 sky130_fd_sc_hd__mux2i_2 _26983_ (.A0(_03691_),
    .A1(_03696_),
    .S(net419),
    .Y(_03697_));
 sky130_fd_sc_hd__xnor2_1 _26984_ (.A(_03567_),
    .B(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__xnor2_2 _26985_ (.A(_03086_),
    .B(_03698_),
    .Y(_11917_));
 sky130_fd_sc_hd__mux4_2 _26986_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03699_));
 sky130_fd_sc_hd__mux4_2 _26987_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03700_));
 sky130_fd_sc_hd__mux4_2 _26988_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03701_));
 sky130_fd_sc_hd__mux4_2 _26989_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03702_));
 sky130_fd_sc_hd__mux4_2 _26990_ (.A0(_03699_),
    .A1(_03700_),
    .A2(_03701_),
    .A3(_03702_),
    .S0(net504),
    .S1(net501),
    .X(_03703_));
 sky130_fd_sc_hd__mux4_2 _26991_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03704_));
 sky130_fd_sc_hd__mux4_2 _26992_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03705_));
 sky130_fd_sc_hd__mux4_2 _26993_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03706_));
 sky130_fd_sc_hd__mux4_2 _26994_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net505),
    .S1(net517),
    .X(_03707_));
 sky130_fd_sc_hd__mux4_2 _26995_ (.A0(_03704_),
    .A1(_03705_),
    .A2(_03706_),
    .A3(_03707_),
    .S0(net504),
    .S1(net501),
    .X(_03708_));
 sky130_fd_sc_hd__mux2i_4 _26996_ (.A0(_03703_),
    .A1(_03708_),
    .S(\count15_2[5] ),
    .Y(_03709_));
 sky130_fd_sc_hd__xnor2_1 _26997_ (.A(_03460_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__xnor2_1 _26998_ (.A(_02853_),
    .B(_03710_),
    .Y(_11916_));
 sky130_fd_sc_hd__mux4_2 _26999_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net388),
    .S1(net398),
    .X(_03711_));
 sky130_fd_sc_hd__mux4_2 _27000_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net388),
    .S1(net398),
    .X(_03712_));
 sky130_fd_sc_hd__mux4_2 _27001_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net388),
    .S1(net398),
    .X(_03713_));
 sky130_fd_sc_hd__mux4_2 _27002_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net388),
    .S1(net398),
    .X(_03714_));
 sky130_fd_sc_hd__mux4_2 _27003_ (.A0(_03711_),
    .A1(_03712_),
    .A2(_03713_),
    .A3(_03714_),
    .S0(net386),
    .S1(net382),
    .X(_03715_));
 sky130_fd_sc_hd__mux4_2 _27004_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net391),
    .S1(net397),
    .X(_03716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__mux4_2 _27006_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net391),
    .S1(net397),
    .X(_03718_));
 sky130_fd_sc_hd__mux4_2 _27007_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net391),
    .S1(net397),
    .X(_03719_));
 sky130_fd_sc_hd__mux4_2 _27008_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net391),
    .S1(net397),
    .X(_03720_));
 sky130_fd_sc_hd__mux4_2 _27009_ (.A0(_03716_),
    .A1(_03718_),
    .A2(_03719_),
    .A3(_03720_),
    .S0(net384),
    .S1(net542),
    .X(_03721_));
 sky130_fd_sc_hd__mux2i_4 _27010_ (.A0(_03715_),
    .A1(_03721_),
    .S(net380),
    .Y(_11915_));
 sky130_fd_sc_hd__mux4_2 _27011_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net466),
    .S1(net474),
    .X(_03722_));
 sky130_fd_sc_hd__mux4_2 _27012_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net466),
    .S1(net474),
    .X(_03723_));
 sky130_fd_sc_hd__mux4_2 _27013_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net466),
    .S1(net474),
    .X(_03724_));
 sky130_fd_sc_hd__mux4_2 _27014_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net466),
    .S1(net474),
    .X(_03725_));
 sky130_fd_sc_hd__mux4_2 _27015_ (.A0(_03722_),
    .A1(_03723_),
    .A2(_03724_),
    .A3(_03725_),
    .S0(net463),
    .S1(net459),
    .X(_03726_));
 sky130_fd_sc_hd__mux4_2 _27016_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net470),
    .S1(net477),
    .X(_03727_));
 sky130_fd_sc_hd__mux4_2 _27017_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net470),
    .S1(net477),
    .X(_03728_));
 sky130_fd_sc_hd__mux4_2 _27018_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net470),
    .S1(net477),
    .X(_03729_));
 sky130_fd_sc_hd__mux4_2 _27019_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net470),
    .S1(net477),
    .X(_03730_));
 sky130_fd_sc_hd__mux4_2 _27020_ (.A0(_03727_),
    .A1(_03728_),
    .A2(_03729_),
    .A3(_03730_),
    .S0(\count16_2[3] ),
    .S1(net461),
    .X(_03731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__mux2i_4 _27022_ (.A0(_03726_),
    .A1(_03731_),
    .S(net457),
    .Y(_11920_));
 sky130_fd_sc_hd__mux4_2 _27023_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net424),
    .S1(net435),
    .X(_03733_));
 sky130_fd_sc_hd__mux4_2 _27024_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net424),
    .S1(net435),
    .X(_03734_));
 sky130_fd_sc_hd__mux4_2 _27025_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net424),
    .S1(net435),
    .X(_03735_));
 sky130_fd_sc_hd__mux4_2 _27026_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net424),
    .S1(net435),
    .X(_03736_));
 sky130_fd_sc_hd__mux4_2 _27027_ (.A0(_03733_),
    .A1(_03734_),
    .A2(_03735_),
    .A3(_03736_),
    .S0(net549),
    .S1(net421),
    .X(_03737_));
 sky130_fd_sc_hd__mux4_2 _27028_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net426),
    .S1(net431),
    .X(_03738_));
 sky130_fd_sc_hd__mux4_2 _27029_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net426),
    .S1(net431),
    .X(_03739_));
 sky130_fd_sc_hd__mux4_2 _27030_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net426),
    .S1(net431),
    .X(_03740_));
 sky130_fd_sc_hd__mux4_2 _27031_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net426),
    .S1(net431),
    .X(_03741_));
 sky130_fd_sc_hd__mux4_2 _27032_ (.A0(_03738_),
    .A1(_03739_),
    .A2(_03740_),
    .A3(_03741_),
    .S0(net549),
    .S1(net421),
    .X(_03742_));
 sky130_fd_sc_hd__mux2i_4 _27033_ (.A0(_03737_),
    .A1(_03742_),
    .S(\count2_2[5] ),
    .Y(_03743_));
 sky130_fd_sc_hd__xnor2_1 _27034_ (.A(_03633_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__xnor2_1 _27035_ (.A(_03168_),
    .B(_03744_),
    .Y(_11925_));
 sky130_fd_sc_hd__mux4_2 _27036_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03745_));
 sky130_fd_sc_hd__mux4_2 _27037_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03746_));
 sky130_fd_sc_hd__mux4_2 _27038_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03747_));
 sky130_fd_sc_hd__mux4_2 _27039_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03748_));
 sky130_fd_sc_hd__mux4_2 _27040_ (.A0(_03745_),
    .A1(_03746_),
    .A2(_03747_),
    .A3(_03748_),
    .S0(net504),
    .S1(net501),
    .X(_03749_));
 sky130_fd_sc_hd__mux4_2 _27041_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03750_));
 sky130_fd_sc_hd__mux4_2 _27042_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03751_));
 sky130_fd_sc_hd__mux4_2 _27043_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03752_));
 sky130_fd_sc_hd__mux4_2 _27044_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net505),
    .S1(net517),
    .X(_03753_));
 sky130_fd_sc_hd__mux4_2 _27045_ (.A0(_03750_),
    .A1(_03751_),
    .A2(_03752_),
    .A3(_03753_),
    .S0(net504),
    .S1(net501),
    .X(_03754_));
 sky130_fd_sc_hd__mux2i_4 _27046_ (.A0(_03749_),
    .A1(_03754_),
    .S(\count15_2[5] ),
    .Y(_03755_));
 sky130_fd_sc_hd__xnor2_1 _27047_ (.A(_03519_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__xnor2_1 _27048_ (.A(net1141),
    .B(_03756_),
    .Y(_11924_));
 sky130_fd_sc_hd__mux4_2 _27049_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net389),
    .S1(net398),
    .X(_03757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__mux4_2 _27051_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net389),
    .S1(net398),
    .X(_03759_));
 sky130_fd_sc_hd__mux4_2 _27052_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net389),
    .S1(net398),
    .X(_03760_));
 sky130_fd_sc_hd__mux4_2 _27053_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net389),
    .S1(net398),
    .X(_03761_));
 sky130_fd_sc_hd__mux4_2 _27054_ (.A0(_03757_),
    .A1(_03759_),
    .A2(_03760_),
    .A3(_03761_),
    .S0(net386),
    .S1(net383),
    .X(_03762_));
 sky130_fd_sc_hd__mux4_2 _27055_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net392),
    .S1(net398),
    .X(_03763_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__mux4_2 _27057_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net392),
    .S1(net544),
    .X(_03765_));
 sky130_fd_sc_hd__mux4_2 _27058_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net392),
    .S1(net544),
    .X(_03766_));
 sky130_fd_sc_hd__mux4_2 _27059_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net392),
    .S1(net544),
    .X(_03767_));
 sky130_fd_sc_hd__mux4_2 _27060_ (.A0(_03763_),
    .A1(_03765_),
    .A2(_03766_),
    .A3(_03767_),
    .S0(net385),
    .S1(\count7_2[4] ),
    .X(_03768_));
 sky130_fd_sc_hd__mux2i_4 _27061_ (.A0(_03762_),
    .A1(_03768_),
    .S(net381),
    .Y(_11923_));
 sky130_fd_sc_hd__mux4_2 _27062_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net466),
    .S1(net474),
    .X(_03769_));
 sky130_fd_sc_hd__mux4_2 _27063_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net466),
    .S1(net474),
    .X(_03770_));
 sky130_fd_sc_hd__mux4_2 _27064_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net466),
    .S1(net474),
    .X(_03771_));
 sky130_fd_sc_hd__mux4_2 _27065_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net466),
    .S1(net474),
    .X(_03772_));
 sky130_fd_sc_hd__mux4_2 _27066_ (.A0(_03769_),
    .A1(_03770_),
    .A2(_03771_),
    .A3(_03772_),
    .S0(net463),
    .S1(net459),
    .X(_03773_));
 sky130_fd_sc_hd__mux4_2 _27067_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net469),
    .S1(net473),
    .X(_03774_));
 sky130_fd_sc_hd__mux4_2 _27068_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net469),
    .S1(net473),
    .X(_03775_));
 sky130_fd_sc_hd__mux4_2 _27069_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net469),
    .S1(net473),
    .X(_03776_));
 sky130_fd_sc_hd__mux4_2 _27070_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net469),
    .S1(net473),
    .X(_03777_));
 sky130_fd_sc_hd__mux4_2 _27071_ (.A0(_03774_),
    .A1(_03775_),
    .A2(_03776_),
    .A3(_03777_),
    .S0(net463),
    .S1(net460),
    .X(_03778_));
 sky130_fd_sc_hd__mux2i_4 _27072_ (.A0(_03773_),
    .A1(_03778_),
    .S(net457),
    .Y(_11928_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__mux4_2 _27075_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__mux4_2 _27078_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__mux4_2 _27081_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03787_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__mux4_2 _27084_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03790_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__mux4_2 _27087_ (.A0(_03781_),
    .A1(_03784_),
    .A2(_03787_),
    .A3(_03790_),
    .S0(net423),
    .S1(net421),
    .X(_03793_));
 sky130_fd_sc_hd__mux4_2 _27088_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03794_));
 sky130_fd_sc_hd__mux4_2 _27089_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03795_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__mux4_2 _27092_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03798_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__mux4_2 _27095_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net426),
    .S1(net431),
    .X(_03801_));
 sky130_fd_sc_hd__mux4_2 _27096_ (.A0(_03794_),
    .A1(_03795_),
    .A2(_03798_),
    .A3(_03801_),
    .S0(net423),
    .S1(net421),
    .X(_03802_));
 sky130_fd_sc_hd__mux2i_4 _27097_ (.A0(_03793_),
    .A1(_03802_),
    .S(net419),
    .Y(_03803_));
 sky130_fd_sc_hd__xnor2_1 _27098_ (.A(_03697_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__xnor2_1 _27099_ (.A(_03250_),
    .B(_03804_),
    .Y(_11933_));
 sky130_fd_sc_hd__mux4_2 _27100_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net510),
    .S1(net516),
    .X(_03805_));
 sky130_fd_sc_hd__mux4_2 _27101_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net510),
    .S1(net516),
    .X(_03806_));
 sky130_fd_sc_hd__mux4_2 _27102_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net510),
    .S1(net516),
    .X(_03807_));
 sky130_fd_sc_hd__mux4_2 _27103_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net510),
    .S1(net516),
    .X(_03808_));
 sky130_fd_sc_hd__mux4_2 _27104_ (.A0(_03805_),
    .A1(_03806_),
    .A2(_03807_),
    .A3(_03808_),
    .S0(net502),
    .S1(net499),
    .X(_03809_));
 sky130_fd_sc_hd__mux4_2 _27105_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net510),
    .S1(net514),
    .X(_03810_));
 sky130_fd_sc_hd__mux4_2 _27106_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net510),
    .S1(net514),
    .X(_03811_));
 sky130_fd_sc_hd__mux4_2 _27107_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net510),
    .S1(net514),
    .X(_03812_));
 sky130_fd_sc_hd__mux4_2 _27108_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net510),
    .S1(net514),
    .X(_03813_));
 sky130_fd_sc_hd__mux4_2 _27109_ (.A0(_03810_),
    .A1(_03811_),
    .A2(_03812_),
    .A3(_03813_),
    .S0(net503),
    .S1(net500),
    .X(_03814_));
 sky130_fd_sc_hd__mux2i_4 _27110_ (.A0(_03809_),
    .A1(_03814_),
    .S(net498),
    .Y(_03815_));
 sky130_fd_sc_hd__xnor2_1 _27111_ (.A(_03579_),
    .B(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__xnor2_1 _27112_ (.A(_03109_),
    .B(_03816_),
    .Y(_11932_));
 sky130_fd_sc_hd__mux4_2 _27113_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net389),
    .S1(net398),
    .X(_03817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__mux4_2 _27115_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net389),
    .S1(net398),
    .X(_03819_));
 sky130_fd_sc_hd__mux4_2 _27116_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net389),
    .S1(net398),
    .X(_03820_));
 sky130_fd_sc_hd__mux4_2 _27117_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net389),
    .S1(net398),
    .X(_03821_));
 sky130_fd_sc_hd__mux4_2 _27118_ (.A0(_03817_),
    .A1(_03819_),
    .A2(_03820_),
    .A3(_03821_),
    .S0(net386),
    .S1(net383),
    .X(_03822_));
 sky130_fd_sc_hd__mux4_2 _27119_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net392),
    .S1(net398),
    .X(_03823_));
 sky130_fd_sc_hd__mux4_2 _27120_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net392),
    .S1(net398),
    .X(_03824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__mux4_2 _27122_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net392),
    .S1(net398),
    .X(_03826_));
 sky130_fd_sc_hd__mux4_2 _27123_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net392),
    .S1(net398),
    .X(_03827_));
 sky130_fd_sc_hd__mux4_2 _27124_ (.A0(_03823_),
    .A1(_03824_),
    .A2(_03826_),
    .A3(_03827_),
    .S0(net385),
    .S1(\count7_2[4] ),
    .X(_03828_));
 sky130_fd_sc_hd__mux2i_4 _27125_ (.A0(_03822_),
    .A1(_03828_),
    .S(net381),
    .Y(_11931_));
 sky130_fd_sc_hd__mux4_2 _27126_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net470),
    .S1(net473),
    .X(_03829_));
 sky130_fd_sc_hd__mux4_2 _27127_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net470),
    .S1(net473),
    .X(_03830_));
 sky130_fd_sc_hd__mux4_2 _27128_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net470),
    .S1(net473),
    .X(_03831_));
 sky130_fd_sc_hd__mux4_2 _27129_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net470),
    .S1(net473),
    .X(_03832_));
 sky130_fd_sc_hd__mux4_2 _27130_ (.A0(_03829_),
    .A1(_03830_),
    .A2(_03831_),
    .A3(_03832_),
    .S0(\count16_2[3] ),
    .S1(net459),
    .X(_03833_));
 sky130_fd_sc_hd__mux4_2 _27131_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net470),
    .S1(net477),
    .X(_03834_));
 sky130_fd_sc_hd__mux4_2 _27132_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net470),
    .S1(net477),
    .X(_03835_));
 sky130_fd_sc_hd__mux4_2 _27133_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net470),
    .S1(net477),
    .X(_03836_));
 sky130_fd_sc_hd__mux4_2 _27134_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net470),
    .S1(net477),
    .X(_03837_));
 sky130_fd_sc_hd__mux4_2 _27135_ (.A0(_03834_),
    .A1(_03835_),
    .A2(_03836_),
    .A3(_03837_),
    .S0(\count16_2[3] ),
    .S1(net461),
    .X(_03838_));
 sky130_fd_sc_hd__mux2i_4 _27136_ (.A0(_03833_),
    .A1(_03838_),
    .S(net457),
    .Y(_11936_));
 sky130_fd_sc_hd__mux4_2 _27137_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03839_));
 sky130_fd_sc_hd__mux4_2 _27138_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03840_));
 sky130_fd_sc_hd__mux4_2 _27139_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03841_));
 sky130_fd_sc_hd__mux4_2 _27140_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03842_));
 sky130_fd_sc_hd__mux4_2 _27141_ (.A0(_03839_),
    .A1(_03840_),
    .A2(_03841_),
    .A3(_03842_),
    .S0(net423),
    .S1(net421),
    .X(_03843_));
 sky130_fd_sc_hd__mux4_2 _27142_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03844_));
 sky130_fd_sc_hd__mux4_2 _27143_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03845_));
 sky130_fd_sc_hd__mux4_2 _27144_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03846_));
 sky130_fd_sc_hd__mux4_2 _27145_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net426),
    .S1(net431),
    .X(_03847_));
 sky130_fd_sc_hd__mux4_2 _27146_ (.A0(_03844_),
    .A1(_03845_),
    .A2(_03846_),
    .A3(_03847_),
    .S0(net423),
    .S1(net421),
    .X(_03848_));
 sky130_fd_sc_hd__mux2i_4 _27147_ (.A0(_03843_),
    .A1(_03848_),
    .S(\count2_2[5] ),
    .Y(_03849_));
 sky130_fd_sc_hd__xnor2_1 _27148_ (.A(_03743_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _27149_ (.A(_03320_),
    .B(_03850_),
    .Y(_11941_));
 sky130_fd_sc_hd__mux4_2 _27150_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__mux4_2 _27152_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__mux4_2 _27155_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03856_));
 sky130_fd_sc_hd__mux4_2 _27156_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03857_));
 sky130_fd_sc_hd__mux4_2 _27157_ (.A0(_03851_),
    .A1(_03853_),
    .A2(_03856_),
    .A3(_03857_),
    .S0(net502),
    .S1(net499),
    .X(_03858_));
 sky130_fd_sc_hd__mux4_2 _27158_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03859_));
 sky130_fd_sc_hd__mux4_2 _27159_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03860_));
 sky130_fd_sc_hd__mux4_2 _27160_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03861_));
 sky130_fd_sc_hd__mux4_2 _27161_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net507),
    .S1(net512),
    .X(_03862_));
 sky130_fd_sc_hd__mux4_2 _27162_ (.A0(_03859_),
    .A1(_03860_),
    .A2(_03861_),
    .A3(_03862_),
    .S0(net503),
    .S1(net500),
    .X(_03863_));
 sky130_fd_sc_hd__mux2i_4 _27163_ (.A0(_03858_),
    .A1(_03863_),
    .S(net497),
    .Y(_03864_));
 sky130_fd_sc_hd__xnor2_1 _27164_ (.A(_03656_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__xnor2_2 _27165_ (.A(_03181_),
    .B(_03865_),
    .Y(_11940_));
 sky130_fd_sc_hd__mux4_2 _27166_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net388),
    .S1(net398),
    .X(_03866_));
 sky130_fd_sc_hd__mux4_2 _27167_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net388),
    .S1(net398),
    .X(_03867_));
 sky130_fd_sc_hd__mux4_2 _27168_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net388),
    .S1(net398),
    .X(_03868_));
 sky130_fd_sc_hd__mux4_2 _27169_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net388),
    .S1(net398),
    .X(_03869_));
 sky130_fd_sc_hd__mux4_2 _27170_ (.A0(_03866_),
    .A1(_03867_),
    .A2(_03868_),
    .A3(_03869_),
    .S0(net386),
    .S1(net383),
    .X(_03870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__mux4_2 _27172_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net392),
    .S1(net397),
    .X(_03872_));
 sky130_fd_sc_hd__mux4_2 _27173_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net392),
    .S1(net544),
    .X(_03873_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__mux4_2 _27175_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net392),
    .S1(net544),
    .X(_03875_));
 sky130_fd_sc_hd__mux4_2 _27176_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net392),
    .S1(net544),
    .X(_03876_));
 sky130_fd_sc_hd__mux4_2 _27177_ (.A0(_03872_),
    .A1(_03873_),
    .A2(_03875_),
    .A3(_03876_),
    .S0(net385),
    .S1(net382),
    .X(_03877_));
 sky130_fd_sc_hd__mux2i_4 _27178_ (.A0(_03870_),
    .A1(_03877_),
    .S(net381),
    .Y(_11939_));
 sky130_fd_sc_hd__mux4_2 _27179_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03878_));
 sky130_fd_sc_hd__mux4_2 _27180_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03879_));
 sky130_fd_sc_hd__mux4_2 _27181_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03880_));
 sky130_fd_sc_hd__mux4_2 _27182_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net466),
    .S1(net474),
    .X(_03881_));
 sky130_fd_sc_hd__mux4_2 _27183_ (.A0(_03878_),
    .A1(_03879_),
    .A2(_03880_),
    .A3(_03881_),
    .S0(net462),
    .S1(net460),
    .X(_03882_));
 sky130_fd_sc_hd__fa_1 _27184_ (.A(_11579_),
    .B(_11580_),
    .CIN(_11581_),
    .COUT(_11582_),
    .SUM(_11583_));
 sky130_fd_sc_hd__fa_1 _27185_ (.A(_11584_),
    .B(_11585_),
    .CIN(_11586_),
    .COUT(_11587_),
    .SUM(_11588_));
 sky130_fd_sc_hd__fa_1 _27186_ (.A(_11589_),
    .B(_11582_),
    .CIN(_11588_),
    .COUT(_11590_),
    .SUM(_11591_));
 sky130_fd_sc_hd__fa_1 _27187_ (.A(_11592_),
    .B(_11593_),
    .CIN(_11594_),
    .COUT(_11595_),
    .SUM(_11596_));
 sky130_fd_sc_hd__fa_1 _27188_ (.A(_11597_),
    .B(_11587_),
    .CIN(_11596_),
    .COUT(_11598_),
    .SUM(_11599_));
 sky130_fd_sc_hd__fa_1 _27189_ (.A(_11600_),
    .B(_11590_),
    .CIN(_11599_),
    .COUT(_11601_),
    .SUM(_11602_));
 sky130_fd_sc_hd__fa_1 _27190_ (.A(_11603_),
    .B(_11604_),
    .CIN(_11605_),
    .COUT(_11606_),
    .SUM(_11607_));
 sky130_fd_sc_hd__fa_1 _27191_ (.A(_11608_),
    .B(_11595_),
    .CIN(_11607_),
    .COUT(_11609_),
    .SUM(_11610_));
 sky130_fd_sc_hd__fa_1 _27192_ (.A(_11611_),
    .B(_11612_),
    .CIN(_11613_),
    .COUT(_11614_),
    .SUM(_11615_));
 sky130_fd_sc_hd__fa_1 _27193_ (.A(_11616_),
    .B(_11606_),
    .CIN(_11615_),
    .COUT(_11617_),
    .SUM(_11618_));
 sky130_fd_sc_hd__fa_1 _27194_ (.A(_11619_),
    .B(_11620_),
    .CIN(_11621_),
    .COUT(_11622_),
    .SUM(_11623_));
 sky130_fd_sc_hd__fa_1 _27195_ (.A(_11624_),
    .B(_11614_),
    .CIN(_11623_),
    .COUT(_11625_),
    .SUM(_11626_));
 sky130_fd_sc_hd__fa_1 _27196_ (.A(_11627_),
    .B(_11628_),
    .CIN(_11629_),
    .COUT(_11630_),
    .SUM(_11631_));
 sky130_fd_sc_hd__fa_1 _27197_ (.A(_11632_),
    .B(_11622_),
    .CIN(_11631_),
    .COUT(_11633_),
    .SUM(_11634_));
 sky130_fd_sc_hd__fa_1 _27198_ (.A(_11635_),
    .B(_11636_),
    .CIN(_11637_),
    .COUT(_11638_),
    .SUM(_11639_));
 sky130_fd_sc_hd__fa_1 _27199_ (.A(_11640_),
    .B(_11630_),
    .CIN(_11639_),
    .COUT(_11641_),
    .SUM(_11642_));
 sky130_fd_sc_hd__fa_1 _27200_ (.A(_11643_),
    .B(_11644_),
    .CIN(_11645_),
    .COUT(_11646_),
    .SUM(_11647_));
 sky130_fd_sc_hd__fa_1 _27201_ (.A(_11648_),
    .B(_11638_),
    .CIN(_11647_),
    .COUT(_11649_),
    .SUM(_11650_));
 sky130_fd_sc_hd__fa_1 _27202_ (.A(_11651_),
    .B(_11652_),
    .CIN(_11653_),
    .COUT(_11654_),
    .SUM(_11655_));
 sky130_fd_sc_hd__fa_1 _27203_ (.A(_11656_),
    .B(_11646_),
    .CIN(_11655_),
    .COUT(_11657_),
    .SUM(_11658_));
 sky130_fd_sc_hd__fa_1 _27204_ (.A(_11659_),
    .B(_11660_),
    .CIN(_11661_),
    .COUT(_11662_),
    .SUM(_11663_));
 sky130_fd_sc_hd__fa_1 _27205_ (.A(_11664_),
    .B(_11654_),
    .CIN(_11663_),
    .COUT(_11665_),
    .SUM(_11666_));
 sky130_fd_sc_hd__fa_1 _27206_ (.A(_11667_),
    .B(_11668_),
    .CIN(_11669_),
    .COUT(_11670_),
    .SUM(_11671_));
 sky130_fd_sc_hd__fa_1 _27207_ (.A(_11672_),
    .B(_11662_),
    .CIN(_11671_),
    .COUT(_11673_),
    .SUM(_11674_));
 sky130_fd_sc_hd__fa_1 _27208_ (.A(_11675_),
    .B(_11676_),
    .CIN(_11677_),
    .COUT(_11678_),
    .SUM(_11679_));
 sky130_fd_sc_hd__fa_1 _27209_ (.A(_11680_),
    .B(_11670_),
    .CIN(_11679_),
    .COUT(_11681_),
    .SUM(_11682_));
 sky130_fd_sc_hd__fa_1 _27210_ (.A(_11683_),
    .B(_11684_),
    .CIN(_11685_),
    .COUT(_11686_),
    .SUM(_11687_));
 sky130_fd_sc_hd__fa_1 _27211_ (.A(_11688_),
    .B(_11678_),
    .CIN(_11687_),
    .COUT(_11689_),
    .SUM(_11690_));
 sky130_fd_sc_hd__fa_1 _27212_ (.A(_11691_),
    .B(_11692_),
    .CIN(_11693_),
    .COUT(_11694_),
    .SUM(_11695_));
 sky130_fd_sc_hd__fa_1 _27213_ (.A(_11696_),
    .B(_11686_),
    .CIN(_11695_),
    .COUT(_11697_),
    .SUM(_11698_));
 sky130_fd_sc_hd__fa_1 _27214_ (.A(_11699_),
    .B(_11700_),
    .CIN(_11701_),
    .COUT(_11702_),
    .SUM(_11703_));
 sky130_fd_sc_hd__fa_1 _27215_ (.A(_11704_),
    .B(_11694_),
    .CIN(_11703_),
    .COUT(_11705_),
    .SUM(_11706_));
 sky130_fd_sc_hd__fa_1 _27216_ (.A(_11707_),
    .B(_11708_),
    .CIN(_11709_),
    .COUT(_11710_),
    .SUM(_11711_));
 sky130_fd_sc_hd__fa_1 _27217_ (.A(_11712_),
    .B(_11702_),
    .CIN(_11711_),
    .COUT(_11713_),
    .SUM(_11714_));
 sky130_fd_sc_hd__fa_1 _27218_ (.A(_11715_),
    .B(_11716_),
    .CIN(_11717_),
    .COUT(_11718_),
    .SUM(_11719_));
 sky130_fd_sc_hd__fa_1 _27219_ (.A(_11720_),
    .B(_11710_),
    .CIN(_11719_),
    .COUT(_11721_),
    .SUM(_11722_));
 sky130_fd_sc_hd__fa_1 _27220_ (.A(_11723_),
    .B(_11724_),
    .CIN(_11725_),
    .COUT(_11726_),
    .SUM(_11727_));
 sky130_fd_sc_hd__fa_1 _27221_ (.A(_11728_),
    .B(_11718_),
    .CIN(_11727_),
    .COUT(_11729_),
    .SUM(_11730_));
 sky130_fd_sc_hd__fa_1 _27222_ (.A(_11731_),
    .B(_11732_),
    .CIN(_11733_),
    .COUT(_11734_),
    .SUM(_11735_));
 sky130_fd_sc_hd__fa_1 _27223_ (.A(_11736_),
    .B(_11726_),
    .CIN(_11735_),
    .COUT(_11737_),
    .SUM(_11738_));
 sky130_fd_sc_hd__fa_1 _27224_ (.A(_11739_),
    .B(_11740_),
    .CIN(_11741_),
    .COUT(_11742_),
    .SUM(_11743_));
 sky130_fd_sc_hd__fa_1 _27225_ (.A(_11744_),
    .B(_11734_),
    .CIN(_11743_),
    .COUT(_11745_),
    .SUM(_11746_));
 sky130_fd_sc_hd__fa_1 _27226_ (.A(_11747_),
    .B(_11748_),
    .CIN(_11749_),
    .COUT(_11750_),
    .SUM(_11751_));
 sky130_fd_sc_hd__fa_1 _27227_ (.A(_11752_),
    .B(_11742_),
    .CIN(_11751_),
    .COUT(_11753_),
    .SUM(_11754_));
 sky130_fd_sc_hd__fa_1 _27228_ (.A(_11755_),
    .B(_11756_),
    .CIN(_11757_),
    .COUT(_11758_),
    .SUM(_11759_));
 sky130_fd_sc_hd__fa_1 _27229_ (.A(_11760_),
    .B(_11750_),
    .CIN(_11759_),
    .COUT(_11761_),
    .SUM(_11762_));
 sky130_fd_sc_hd__fa_1 _27230_ (.A(_11763_),
    .B(_11764_),
    .CIN(_11765_),
    .COUT(_11766_),
    .SUM(_11767_));
 sky130_fd_sc_hd__fa_1 _27231_ (.A(_11768_),
    .B(_11758_),
    .CIN(_11767_),
    .COUT(_11769_),
    .SUM(_11770_));
 sky130_fd_sc_hd__fa_1 _27232_ (.A(_11771_),
    .B(_11772_),
    .CIN(_11773_),
    .COUT(_11774_),
    .SUM(_11775_));
 sky130_fd_sc_hd__fa_1 _27233_ (.A(_11776_),
    .B(_11766_),
    .CIN(_11775_),
    .COUT(_11777_),
    .SUM(_11778_));
 sky130_fd_sc_hd__fa_1 _27234_ (.A(_11779_),
    .B(_11780_),
    .CIN(_11781_),
    .COUT(_11782_),
    .SUM(_11783_));
 sky130_fd_sc_hd__fa_1 _27235_ (.A(_11784_),
    .B(_11774_),
    .CIN(_11783_),
    .COUT(_11785_),
    .SUM(_11786_));
 sky130_fd_sc_hd__fa_1 _27236_ (.A(_11787_),
    .B(_11788_),
    .CIN(_11789_),
    .COUT(_11790_),
    .SUM(_11791_));
 sky130_fd_sc_hd__fa_1 _27237_ (.A(_11792_),
    .B(_11782_),
    .CIN(_11791_),
    .COUT(_11793_),
    .SUM(_11794_));
 sky130_fd_sc_hd__fa_1 _27238_ (.A(_11795_),
    .B(_11796_),
    .CIN(_11797_),
    .COUT(_11798_),
    .SUM(_11799_));
 sky130_fd_sc_hd__fa_1 _27239_ (.A(_11800_),
    .B(_11790_),
    .CIN(_11799_),
    .COUT(_11801_),
    .SUM(_11802_));
 sky130_fd_sc_hd__fa_1 _27240_ (.A(_11803_),
    .B(_11804_),
    .CIN(_11805_),
    .COUT(_11806_),
    .SUM(_11807_));
 sky130_fd_sc_hd__fa_1 _27241_ (.A(_11808_),
    .B(_11798_),
    .CIN(_11807_),
    .COUT(_11809_),
    .SUM(_11810_));
 sky130_fd_sc_hd__fa_1 _27242_ (.A(_11811_),
    .B(_11812_),
    .CIN(_11813_),
    .COUT(_11814_),
    .SUM(_11815_));
 sky130_fd_sc_hd__fa_1 _27243_ (.A(_11816_),
    .B(_11806_),
    .CIN(_11815_),
    .COUT(_11817_),
    .SUM(_11818_));
 sky130_fd_sc_hd__fa_1 _27244_ (.A(_11819_),
    .B(_11820_),
    .CIN(_11821_),
    .COUT(_11822_),
    .SUM(_11823_));
 sky130_fd_sc_hd__fa_1 _27245_ (.A(_11824_),
    .B(_11814_),
    .CIN(_11823_),
    .COUT(_11825_),
    .SUM(_11826_));
 sky130_fd_sc_hd__fa_1 _27246_ (.A(_11827_),
    .B(_11828_),
    .CIN(_11829_),
    .COUT(_11830_),
    .SUM(_11831_));
 sky130_fd_sc_hd__fa_1 _27247_ (.A(_11832_),
    .B(_11833_),
    .CIN(_11834_),
    .COUT(_11835_),
    .SUM(_11836_));
 sky130_fd_sc_hd__fa_1 _27248_ (.A(_11837_),
    .B(_11830_),
    .CIN(_11836_),
    .COUT(_11838_),
    .SUM(_11839_));
 sky130_fd_sc_hd__fa_1 _27249_ (.A(_11840_),
    .B(_11841_),
    .CIN(_11842_),
    .COUT(_11843_),
    .SUM(_11844_));
 sky130_fd_sc_hd__fa_1 _27250_ (.A(_11845_),
    .B(_11835_),
    .CIN(_11844_),
    .COUT(_11846_),
    .SUM(_11847_));
 sky130_fd_sc_hd__fa_1 _27251_ (.A(_11848_),
    .B(_11838_),
    .CIN(_11847_),
    .COUT(_11849_),
    .SUM(_11850_));
 sky130_fd_sc_hd__fa_1 _27252_ (.A(_11851_),
    .B(_11852_),
    .CIN(_11853_),
    .COUT(_11854_),
    .SUM(_11855_));
 sky130_fd_sc_hd__fa_1 _27253_ (.A(_11856_),
    .B(_11843_),
    .CIN(_11855_),
    .COUT(_11857_),
    .SUM(_11858_));
 sky130_fd_sc_hd__fa_1 _27254_ (.A(_11859_),
    .B(_11860_),
    .CIN(_11861_),
    .COUT(_11862_),
    .SUM(_11863_));
 sky130_fd_sc_hd__fa_1 _27255_ (.A(_11864_),
    .B(_11854_),
    .CIN(_11863_),
    .COUT(_11865_),
    .SUM(_11866_));
 sky130_fd_sc_hd__fa_1 _27256_ (.A(_11867_),
    .B(_11868_),
    .CIN(_11869_),
    .COUT(_11870_),
    .SUM(_11871_));
 sky130_fd_sc_hd__fa_1 _27257_ (.A(_11872_),
    .B(_11862_),
    .CIN(_11871_),
    .COUT(_11873_),
    .SUM(_11874_));
 sky130_fd_sc_hd__fa_1 _27258_ (.A(_11875_),
    .B(_11876_),
    .CIN(_11877_),
    .COUT(_11878_),
    .SUM(_11879_));
 sky130_fd_sc_hd__fa_1 _27259_ (.A(_11880_),
    .B(_11870_),
    .CIN(_11879_),
    .COUT(_11881_),
    .SUM(_11882_));
 sky130_fd_sc_hd__fa_1 _27260_ (.A(_11883_),
    .B(_11884_),
    .CIN(_11885_),
    .COUT(_11886_),
    .SUM(_11887_));
 sky130_fd_sc_hd__fa_1 _27261_ (.A(_11888_),
    .B(_11878_),
    .CIN(_11887_),
    .COUT(_11889_),
    .SUM(_11890_));
 sky130_fd_sc_hd__fa_1 _27262_ (.A(_11891_),
    .B(_11892_),
    .CIN(_11893_),
    .COUT(_11894_),
    .SUM(_11895_));
 sky130_fd_sc_hd__fa_1 _27263_ (.A(_11896_),
    .B(_11886_),
    .CIN(_11895_),
    .COUT(_11897_),
    .SUM(_11898_));
 sky130_fd_sc_hd__fa_1 _27264_ (.A(_11899_),
    .B(_11900_),
    .CIN(_11901_),
    .COUT(_11902_),
    .SUM(_11903_));
 sky130_fd_sc_hd__fa_1 _27265_ (.A(_11904_),
    .B(_11894_),
    .CIN(_11903_),
    .COUT(_11905_),
    .SUM(_11906_));
 sky130_fd_sc_hd__fa_1 _27266_ (.A(_11907_),
    .B(_11908_),
    .CIN(_11909_),
    .COUT(_11910_),
    .SUM(_11911_));
 sky130_fd_sc_hd__fa_1 _27267_ (.A(_11912_),
    .B(_11902_),
    .CIN(_11911_),
    .COUT(_11913_),
    .SUM(_11914_));
 sky130_fd_sc_hd__fa_1 _27268_ (.A(_11915_),
    .B(_11916_),
    .CIN(_11917_),
    .COUT(_11918_),
    .SUM(_11919_));
 sky130_fd_sc_hd__fa_1 _27269_ (.A(_11920_),
    .B(_11910_),
    .CIN(_11919_),
    .COUT(_11921_),
    .SUM(_11922_));
 sky130_fd_sc_hd__fa_1 _27270_ (.A(_11923_),
    .B(_11924_),
    .CIN(_11925_),
    .COUT(_11926_),
    .SUM(_11927_));
 sky130_fd_sc_hd__fa_1 _27271_ (.A(_11928_),
    .B(_11918_),
    .CIN(_11927_),
    .COUT(_11929_),
    .SUM(_11930_));
 sky130_fd_sc_hd__fa_1 _27272_ (.A(_11931_),
    .B(_11932_),
    .CIN(_11933_),
    .COUT(_11934_),
    .SUM(_11935_));
 sky130_fd_sc_hd__fa_1 _27273_ (.A(_11936_),
    .B(_11926_),
    .CIN(_11935_),
    .COUT(_11937_),
    .SUM(_11938_));
 sky130_fd_sc_hd__fa_1 _27274_ (.A(_11939_),
    .B(_11940_),
    .CIN(_11941_),
    .COUT(_11942_),
    .SUM(_11943_));
 sky130_fd_sc_hd__fa_1 _27275_ (.A(_11944_),
    .B(_11934_),
    .CIN(_11943_),
    .COUT(_11945_),
    .SUM(_11946_));
 sky130_fd_sc_hd__fa_1 _27276_ (.A(_11947_),
    .B(_11948_),
    .CIN(_11949_),
    .COUT(_11950_),
    .SUM(_11951_));
 sky130_fd_sc_hd__fa_1 _27277_ (.A(_11952_),
    .B(_11942_),
    .CIN(_11951_),
    .COUT(_11953_),
    .SUM(_11954_));
 sky130_fd_sc_hd__fa_1 _27278_ (.A(_11955_),
    .B(_11956_),
    .CIN(_11957_),
    .COUT(_11958_),
    .SUM(_11959_));
 sky130_fd_sc_hd__fa_1 _27279_ (.A(_11960_),
    .B(_11950_),
    .CIN(_11959_),
    .COUT(_11961_),
    .SUM(_11962_));
 sky130_fd_sc_hd__fa_1 _27280_ (.A(_11963_),
    .B(_11964_),
    .CIN(_11965_),
    .COUT(_11966_),
    .SUM(_11967_));
 sky130_fd_sc_hd__fa_1 _27281_ (.A(_11968_),
    .B(_11958_),
    .CIN(_11967_),
    .COUT(_11969_),
    .SUM(_11970_));
 sky130_fd_sc_hd__fa_1 _27282_ (.A(_11971_),
    .B(_11972_),
    .CIN(_11973_),
    .COUT(_11974_),
    .SUM(_11975_));
 sky130_fd_sc_hd__fa_1 _27283_ (.A(_11976_),
    .B(_11966_),
    .CIN(_11975_),
    .COUT(_11977_),
    .SUM(_11978_));
 sky130_fd_sc_hd__fa_1 _27284_ (.A(_11979_),
    .B(_11980_),
    .CIN(_11981_),
    .COUT(_11982_),
    .SUM(_11983_));
 sky130_fd_sc_hd__fa_1 _27285_ (.A(_11984_),
    .B(_11974_),
    .CIN(_11983_),
    .COUT(_11985_),
    .SUM(_11986_));
 sky130_fd_sc_hd__fa_1 _27286_ (.A(_11987_),
    .B(_11988_),
    .CIN(_11989_),
    .COUT(_11990_),
    .SUM(_11991_));
 sky130_fd_sc_hd__fa_1 _27287_ (.A(_11992_),
    .B(_11982_),
    .CIN(_11991_),
    .COUT(_11993_),
    .SUM(_11994_));
 sky130_fd_sc_hd__fa_1 _27288_ (.A(_11995_),
    .B(_11996_),
    .CIN(_11997_),
    .COUT(_11998_),
    .SUM(_11999_));
 sky130_fd_sc_hd__fa_1 _27289_ (.A(_12000_),
    .B(_11990_),
    .CIN(_11999_),
    .COUT(_12001_),
    .SUM(_12002_));
 sky130_fd_sc_hd__fa_1 _27290_ (.A(_12003_),
    .B(_12004_),
    .CIN(_12005_),
    .COUT(_12006_),
    .SUM(_12007_));
 sky130_fd_sc_hd__fa_1 _27291_ (.A(_12008_),
    .B(_11998_),
    .CIN(_12007_),
    .COUT(_12009_),
    .SUM(_12010_));
 sky130_fd_sc_hd__fa_1 _27292_ (.A(_12011_),
    .B(_12012_),
    .CIN(_12013_),
    .COUT(_12014_),
    .SUM(_12015_));
 sky130_fd_sc_hd__fa_1 _27293_ (.A(_12016_),
    .B(_12006_),
    .CIN(_12015_),
    .COUT(_12017_),
    .SUM(_12018_));
 sky130_fd_sc_hd__fa_1 _27294_ (.A(_12019_),
    .B(_12020_),
    .CIN(_12021_),
    .COUT(_12022_),
    .SUM(_12023_));
 sky130_fd_sc_hd__fa_1 _27295_ (.A(_12024_),
    .B(_12014_),
    .CIN(_12023_),
    .COUT(_12025_),
    .SUM(_12026_));
 sky130_fd_sc_hd__fa_1 _27296_ (.A(_12027_),
    .B(_12028_),
    .CIN(_12029_),
    .COUT(_12030_),
    .SUM(_12031_));
 sky130_fd_sc_hd__fa_1 _27297_ (.A(_12032_),
    .B(_12022_),
    .CIN(_12031_),
    .COUT(_12033_),
    .SUM(_12034_));
 sky130_fd_sc_hd__fa_1 _27298_ (.A(_12035_),
    .B(_12036_),
    .CIN(_12037_),
    .COUT(_12038_),
    .SUM(_12039_));
 sky130_fd_sc_hd__fa_1 _27299_ (.A(_12040_),
    .B(_12030_),
    .CIN(_12039_),
    .COUT(_12041_),
    .SUM(_12042_));
 sky130_fd_sc_hd__fa_1 _27300_ (.A(_12043_),
    .B(_12044_),
    .CIN(_12045_),
    .COUT(_12046_),
    .SUM(_12047_));
 sky130_fd_sc_hd__fa_1 _27301_ (.A(_12048_),
    .B(_12038_),
    .CIN(_12047_),
    .COUT(_12049_),
    .SUM(_12050_));
 sky130_fd_sc_hd__fa_1 _27302_ (.A(_12051_),
    .B(_12052_),
    .CIN(_12053_),
    .COUT(_12054_),
    .SUM(_12055_));
 sky130_fd_sc_hd__fa_1 _27303_ (.A(_12056_),
    .B(_12046_),
    .CIN(_12055_),
    .COUT(_12057_),
    .SUM(_12058_));
 sky130_fd_sc_hd__fa_1 _27304_ (.A(_12059_),
    .B(_12060_),
    .CIN(_12061_),
    .COUT(_12062_),
    .SUM(_12063_));
 sky130_fd_sc_hd__fa_1 _27305_ (.A(_12064_),
    .B(_12054_),
    .CIN(_12063_),
    .COUT(_12065_),
    .SUM(_12066_));
 sky130_fd_sc_hd__fa_1 _27306_ (.A(_12067_),
    .B(_12068_),
    .CIN(_12069_),
    .COUT(_12070_),
    .SUM(_12071_));
 sky130_fd_sc_hd__fa_1 _27307_ (.A(_12072_),
    .B(_12062_),
    .CIN(_12071_),
    .COUT(_12073_),
    .SUM(_12074_));
 sky130_fd_sc_hd__fa_1 _27308_ (.A(_12075_),
    .B(_12076_),
    .CIN(_12077_),
    .COUT(_12078_),
    .SUM(_12079_));
 sky130_fd_sc_hd__fa_4 _27309_ (.A(\hash.CA2.p1[1] ),
    .B(_12080_),
    .CIN(\hash.CA2.p3[1] ),
    .COUT(_12081_),
    .SUM(_12082_));
 sky130_fd_sc_hd__fa_2 _27310_ (.A(_12083_),
    .B(_12084_),
    .CIN(_12085_),
    .COUT(_12086_),
    .SUM(_12087_));
 sky130_fd_sc_hd__fa_1 _27311_ (.A(_12088_),
    .B(_12087_),
    .CIN(_12089_),
    .COUT(_12090_),
    .SUM(_12091_));
 sky130_fd_sc_hd__fa_1 _27312_ (.A(\hash.CA2.p4[1] ),
    .B(_12092_),
    .CIN(_12093_),
    .COUT(_12094_),
    .SUM(_12095_));
 sky130_fd_sc_hd__fa_1 _27313_ (.A(_12096_),
    .B(_12097_),
    .CIN(_12098_),
    .COUT(_12099_),
    .SUM(_12100_));
 sky130_fd_sc_hd__fa_1 _27314_ (.A(\hash.CA2.p4[2] ),
    .B(_12101_),
    .CIN(_12102_),
    .COUT(_12103_),
    .SUM(_12104_));
 sky130_fd_sc_hd__fa_1 _27315_ (.A(_12105_),
    .B(_12106_),
    .CIN(_12107_),
    .COUT(_12108_),
    .SUM(_12109_));
 sky130_fd_sc_hd__fa_1 _27316_ (.A(_12110_),
    .B(_12111_),
    .CIN(_12112_),
    .COUT(_12113_),
    .SUM(_12114_));
 sky130_fd_sc_hd__fa_1 _27317_ (.A(\hash.CA2.p4[3] ),
    .B(_12115_),
    .CIN(_12116_),
    .COUT(_12117_),
    .SUM(_12118_));
 sky130_fd_sc_hd__fa_1 _27318_ (.A(_12119_),
    .B(_12120_),
    .CIN(_12121_),
    .COUT(_12122_),
    .SUM(_12123_));
 sky130_fd_sc_hd__fa_1 _27319_ (.A(\hash.CA2.p4[4] ),
    .B(_12124_),
    .CIN(_12125_),
    .COUT(_12126_),
    .SUM(_12127_));
 sky130_fd_sc_hd__fa_1 _27320_ (.A(_12128_),
    .B(_12129_),
    .CIN(_12130_),
    .COUT(_12131_),
    .SUM(_12132_));
 sky130_fd_sc_hd__fa_1 _27321_ (.A(\hash.CA2.p4[5] ),
    .B(_12133_),
    .CIN(_12134_),
    .COUT(_12135_),
    .SUM(_12136_));
 sky130_fd_sc_hd__fa_1 _27322_ (.A(_12137_),
    .B(_12138_),
    .CIN(_12139_),
    .COUT(_12140_),
    .SUM(_12141_));
 sky130_fd_sc_hd__fa_1 _27323_ (.A(\hash.CA2.p4[6] ),
    .B(_12142_),
    .CIN(_12143_),
    .COUT(_12144_),
    .SUM(_12145_));
 sky130_fd_sc_hd__fa_1 _27324_ (.A(_12146_),
    .B(_12147_),
    .CIN(_12148_),
    .COUT(_12149_),
    .SUM(_12150_));
 sky130_fd_sc_hd__fa_1 _27325_ (.A(\hash.CA2.p4[7] ),
    .B(_12151_),
    .CIN(_12152_),
    .COUT(_12153_),
    .SUM(_12154_));
 sky130_fd_sc_hd__fa_1 _27326_ (.A(_12157_),
    .B(_12156_),
    .CIN(_12155_),
    .COUT(_12158_),
    .SUM(_12159_));
 sky130_fd_sc_hd__fa_2 _27327_ (.A(\hash.CA2.p4[8] ),
    .B(_12161_),
    .CIN(_12160_),
    .COUT(_12162_),
    .SUM(_12163_));
 sky130_fd_sc_hd__fa_1 _27328_ (.A(_12164_),
    .B(_12165_),
    .CIN(_12166_),
    .COUT(_12167_),
    .SUM(_12168_));
 sky130_fd_sc_hd__fa_1 _27329_ (.A(\hash.CA2.p4[9] ),
    .B(_12169_),
    .CIN(_12170_),
    .COUT(_12171_),
    .SUM(_12172_));
 sky130_fd_sc_hd__fa_1 _27330_ (.A(_12173_),
    .B(_12174_),
    .CIN(_12175_),
    .COUT(_12176_),
    .SUM(_12177_));
 sky130_fd_sc_hd__fa_1 _27331_ (.A(\hash.CA2.p4[10] ),
    .B(_12178_),
    .CIN(_12179_),
    .COUT(_12180_),
    .SUM(_12181_));
 sky130_fd_sc_hd__fa_1 _27332_ (.A(_12182_),
    .B(_12183_),
    .CIN(_12184_),
    .COUT(_12185_),
    .SUM(_12186_));
 sky130_fd_sc_hd__fa_1 _27333_ (.A(\hash.CA2.p4[11] ),
    .B(_12187_),
    .CIN(_12188_),
    .COUT(_12189_),
    .SUM(_12190_));
 sky130_fd_sc_hd__fa_1 _27334_ (.A(_12191_),
    .B(_12192_),
    .CIN(_12193_),
    .COUT(_12194_),
    .SUM(_12195_));
 sky130_fd_sc_hd__fa_1 _27335_ (.A(\hash.CA2.p4[12] ),
    .B(_12196_),
    .CIN(_12197_),
    .COUT(_12198_),
    .SUM(_12199_));
 sky130_fd_sc_hd__fa_1 _27336_ (.A(_12200_),
    .B(_12201_),
    .CIN(_12202_),
    .COUT(_12203_),
    .SUM(_12204_));
 sky130_fd_sc_hd__fa_1 _27337_ (.A(\hash.CA2.p4[13] ),
    .B(_12205_),
    .CIN(_12206_),
    .COUT(_12207_),
    .SUM(_12208_));
 sky130_fd_sc_hd__fa_1 _27338_ (.A(_12209_),
    .B(_12210_),
    .CIN(_12211_),
    .COUT(_12212_),
    .SUM(_12213_));
 sky130_fd_sc_hd__fa_1 _27339_ (.A(\hash.CA2.p4[14] ),
    .B(_12214_),
    .CIN(_12215_),
    .COUT(_12216_),
    .SUM(_12217_));
 sky130_fd_sc_hd__fa_1 _27340_ (.A(_12218_),
    .B(_12219_),
    .CIN(_12220_),
    .COUT(_12221_),
    .SUM(_12222_));
 sky130_fd_sc_hd__fa_1 _27341_ (.A(\hash.CA2.p4[15] ),
    .B(_12223_),
    .CIN(_12224_),
    .COUT(_12225_),
    .SUM(_12226_));
 sky130_fd_sc_hd__fa_1 _27342_ (.A(_12227_),
    .B(_12228_),
    .CIN(_12229_),
    .COUT(_12230_),
    .SUM(_12231_));
 sky130_fd_sc_hd__fa_1 _27343_ (.A(\hash.CA2.p4[16] ),
    .B(_12232_),
    .CIN(_12233_),
    .COUT(_12234_),
    .SUM(_12235_));
 sky130_fd_sc_hd__fa_1 _27344_ (.A(_12238_),
    .B(_12237_),
    .CIN(_12236_),
    .COUT(_12239_),
    .SUM(_12240_));
 sky130_fd_sc_hd__fa_1 _27345_ (.A(\hash.CA2.p4[17] ),
    .B(_12242_),
    .CIN(_12241_),
    .COUT(_12243_),
    .SUM(_12244_));
 sky130_fd_sc_hd__fa_1 _27346_ (.A(_12245_),
    .B(_12246_),
    .CIN(_12247_),
    .COUT(_12248_),
    .SUM(_12249_));
 sky130_fd_sc_hd__fa_1 _27347_ (.A(\hash.CA2.p4[18] ),
    .B(_12250_),
    .CIN(_12251_),
    .COUT(_12252_),
    .SUM(_12253_));
 sky130_fd_sc_hd__fa_1 _27348_ (.A(_12254_),
    .B(_12255_),
    .CIN(_12256_),
    .COUT(_12257_),
    .SUM(_12258_));
 sky130_fd_sc_hd__fa_1 _27349_ (.A(\hash.CA2.p4[19] ),
    .B(_12259_),
    .CIN(_12260_),
    .COUT(_12261_),
    .SUM(_12262_));
 sky130_fd_sc_hd__fa_1 _27350_ (.A(_12263_),
    .B(_12264_),
    .CIN(_12265_),
    .COUT(_12266_),
    .SUM(_12267_));
 sky130_fd_sc_hd__fa_1 _27351_ (.A(\hash.CA2.p4[20] ),
    .B(_12268_),
    .CIN(_12269_),
    .COUT(_12270_),
    .SUM(_12271_));
 sky130_fd_sc_hd__fa_1 _27352_ (.A(_12272_),
    .B(_12273_),
    .CIN(_12274_),
    .COUT(_12275_),
    .SUM(_12276_));
 sky130_fd_sc_hd__fa_1 _27353_ (.A(\hash.CA2.p4[21] ),
    .B(_12277_),
    .CIN(_12278_),
    .COUT(_12279_),
    .SUM(_12280_));
 sky130_fd_sc_hd__fa_1 _27354_ (.A(_12281_),
    .B(_12282_),
    .CIN(_12283_),
    .COUT(_12284_),
    .SUM(_12285_));
 sky130_fd_sc_hd__fa_1 _27355_ (.A(\hash.CA2.p4[22] ),
    .B(_12286_),
    .CIN(_12287_),
    .COUT(_12288_),
    .SUM(_12289_));
 sky130_fd_sc_hd__fa_1 _27356_ (.A(_12290_),
    .B(_12291_),
    .CIN(_12292_),
    .COUT(_12293_),
    .SUM(_12294_));
 sky130_fd_sc_hd__fa_1 _27357_ (.A(\hash.CA2.p4[23] ),
    .B(_12295_),
    .CIN(_12296_),
    .COUT(_12297_),
    .SUM(_12298_));
 sky130_fd_sc_hd__fa_1 _27358_ (.A(_12299_),
    .B(_12300_),
    .CIN(_12301_),
    .COUT(_12302_),
    .SUM(_12303_));
 sky130_fd_sc_hd__fa_1 _27359_ (.A(\hash.CA2.p4[24] ),
    .B(_12304_),
    .CIN(_12305_),
    .COUT(_12306_),
    .SUM(_12307_));
 sky130_fd_sc_hd__fa_1 _27360_ (.A(_12308_),
    .B(_12309_),
    .CIN(_12310_),
    .COUT(_12311_),
    .SUM(_12312_));
 sky130_fd_sc_hd__fa_1 _27361_ (.A(\hash.CA2.p4[25] ),
    .B(_12313_),
    .CIN(_12314_),
    .COUT(_12315_),
    .SUM(_12316_));
 sky130_fd_sc_hd__fa_1 _27362_ (.A(_12317_),
    .B(_12318_),
    .CIN(_12319_),
    .COUT(_12320_),
    .SUM(_12321_));
 sky130_fd_sc_hd__fa_1 _27363_ (.A(\hash.CA2.p4[26] ),
    .B(_12322_),
    .CIN(_12323_),
    .COUT(_12324_),
    .SUM(_12325_));
 sky130_fd_sc_hd__fa_1 _27364_ (.A(_12326_),
    .B(_12327_),
    .CIN(_12328_),
    .COUT(_12329_),
    .SUM(_12330_));
 sky130_fd_sc_hd__fa_1 _27365_ (.A(\hash.CA2.p4[27] ),
    .B(_12331_),
    .CIN(_12332_),
    .COUT(_12333_),
    .SUM(_12334_));
 sky130_fd_sc_hd__fa_1 _27366_ (.A(_12335_),
    .B(_12336_),
    .CIN(_12337_),
    .COUT(_12338_),
    .SUM(_12339_));
 sky130_fd_sc_hd__fa_1 _27367_ (.A(\hash.CA2.p4[28] ),
    .B(_12340_),
    .CIN(_12341_),
    .COUT(_12342_),
    .SUM(_12343_));
 sky130_fd_sc_hd__fa_1 _27368_ (.A(_12344_),
    .B(_12345_),
    .CIN(_12346_),
    .COUT(_12347_),
    .SUM(_12348_));
 sky130_fd_sc_hd__fa_1 _27369_ (.A(\hash.CA2.p4[29] ),
    .B(_12349_),
    .CIN(_12350_),
    .COUT(_12351_),
    .SUM(_12352_));
 sky130_fd_sc_hd__fa_1 _27370_ (.A(_12353_),
    .B(_12354_),
    .CIN(_12355_),
    .COUT(_12356_),
    .SUM(_12357_));
 sky130_fd_sc_hd__fa_1 _27371_ (.A(\hash.CA2.p4[30] ),
    .B(_12358_),
    .CIN(_12359_),
    .COUT(_12360_),
    .SUM(_12361_));
 sky130_fd_sc_hd__fa_2 _27372_ (.A(\hash.CA2.p5[1] ),
    .B(_12362_),
    .CIN(_12363_),
    .COUT(_12364_),
    .SUM(_12365_));
 sky130_fd_sc_hd__fa_1 _27373_ (.A(_12366_),
    .B(_12367_),
    .CIN(_12368_),
    .COUT(_12369_),
    .SUM(_12370_));
 sky130_fd_sc_hd__fa_1 _27374_ (.A(_12371_),
    .B(_12372_),
    .CIN(_00843_),
    .COUT(_12373_),
    .SUM(_12374_));
 sky130_fd_sc_hd__fa_1 _27375_ (.A(\hash.CA1.k_i2[2] ),
    .B(\hash.CA1.w_i2[2] ),
    .CIN(_12375_),
    .COUT(_12376_),
    .SUM(_12377_));
 sky130_fd_sc_hd__fa_1 _27376_ (.A(_12378_),
    .B(_12379_),
    .CIN(_12377_),
    .COUT(_12380_),
    .SUM(\hash.CA1.p4[2] ));
 sky130_fd_sc_hd__fa_1 _27377_ (.A(_12381_),
    .B(_12382_),
    .CIN(_12383_),
    .COUT(_12384_),
    .SUM(_12385_));
 sky130_fd_sc_hd__fa_1 _27378_ (.A(\hash.CA1.k_i2[4] ),
    .B(\hash.CA1.w_i2[4] ),
    .CIN(_12386_),
    .COUT(_12387_),
    .SUM(_12388_));
 sky130_fd_sc_hd__fa_1 _27379_ (.A(_12389_),
    .B(_12390_),
    .CIN(_12391_),
    .COUT(_12392_),
    .SUM(_12393_));
 sky130_fd_sc_hd__fa_1 _27380_ (.A(\hash.CA1.k_i2[6] ),
    .B(\hash.CA1.w_i2[6] ),
    .CIN(_12394_),
    .COUT(_12395_),
    .SUM(_12396_));
 sky130_fd_sc_hd__fa_1 _27381_ (.A(_12397_),
    .B(_12398_),
    .CIN(_12399_),
    .COUT(_12400_),
    .SUM(_12401_));
 sky130_fd_sc_hd__fa_1 _27382_ (.A(_12402_),
    .B(_12403_),
    .CIN(_12404_),
    .COUT(_12405_),
    .SUM(_12406_));
 sky130_fd_sc_hd__fa_2 _27383_ (.A(\hash.CA1.k_i2[9] ),
    .B(\hash.CA1.w_i2[9] ),
    .CIN(_12407_),
    .COUT(_12408_),
    .SUM(_12409_));
 sky130_fd_sc_hd__fa_1 _27384_ (.A(\hash.CA1.k_i2[10] ),
    .B(\hash.CA1.w_i2[10] ),
    .CIN(_12410_),
    .COUT(_12411_),
    .SUM(_12412_));
 sky130_fd_sc_hd__fa_1 _27385_ (.A(_12413_),
    .B(_12414_),
    .CIN(_12415_),
    .COUT(_12416_),
    .SUM(_12417_));
 sky130_fd_sc_hd__fa_1 _27386_ (.A(_12418_),
    .B(_12419_),
    .CIN(_12420_),
    .COUT(_12421_),
    .SUM(_12422_));
 sky130_fd_sc_hd__fa_1 _27387_ (.A(\hash.CA1.k_i2[13] ),
    .B(\hash.CA1.w_i2[13] ),
    .CIN(_12423_),
    .COUT(_12424_),
    .SUM(_12425_));
 sky130_fd_sc_hd__fa_1 _27388_ (.A(_12426_),
    .B(_12427_),
    .CIN(_12428_),
    .COUT(_12429_),
    .SUM(_12430_));
 sky130_fd_sc_hd__fa_1 _27389_ (.A(_12431_),
    .B(_12432_),
    .CIN(_12433_),
    .COUT(_12434_),
    .SUM(_12435_));
 sky130_fd_sc_hd__fa_1 _27390_ (.A(_12436_),
    .B(_12437_),
    .CIN(_12438_),
    .COUT(_12439_),
    .SUM(_12440_));
 sky130_fd_sc_hd__fa_1 _27391_ (.A(_12441_),
    .B(_12442_),
    .CIN(_12443_),
    .COUT(_12444_),
    .SUM(_12445_));
 sky130_fd_sc_hd__fa_1 _27392_ (.A(\hash.CA1.k_i2[18] ),
    .B(\hash.CA1.w_i2[18] ),
    .CIN(_12446_),
    .COUT(_12447_),
    .SUM(_12448_));
 sky130_fd_sc_hd__fa_1 _27393_ (.A(\hash.CA1.k_i2[19] ),
    .B(\hash.CA1.w_i2[19] ),
    .CIN(_12449_),
    .COUT(_12450_),
    .SUM(_12451_));
 sky130_fd_sc_hd__fa_1 _27394_ (.A(\hash.CA1.k_i2[20] ),
    .B(\hash.CA1.w_i2[20] ),
    .CIN(_12452_),
    .COUT(_12453_),
    .SUM(_12454_));
 sky130_fd_sc_hd__fa_1 _27395_ (.A(\hash.CA1.k_i2[21] ),
    .B(\hash.CA1.w_i2[21] ),
    .CIN(_12455_),
    .COUT(_12456_),
    .SUM(_12457_));
 sky130_fd_sc_hd__fa_1 _27396_ (.A(\hash.CA1.k_i2[22] ),
    .B(\hash.CA1.w_i2[22] ),
    .CIN(_12458_),
    .COUT(_12459_),
    .SUM(_12460_));
 sky130_fd_sc_hd__fa_1 _27397_ (.A(_12461_),
    .B(_12462_),
    .CIN(_12463_),
    .COUT(_12464_),
    .SUM(_12465_));
 sky130_fd_sc_hd__fa_1 _27398_ (.A(_12466_),
    .B(_12467_),
    .CIN(_12468_),
    .COUT(_12469_),
    .SUM(_12470_));
 sky130_fd_sc_hd__fa_1 _27399_ (.A(_12471_),
    .B(_12472_),
    .CIN(_12473_),
    .COUT(_12474_),
    .SUM(_12475_));
 sky130_fd_sc_hd__fa_1 _27400_ (.A(_12476_),
    .B(_12477_),
    .CIN(_12478_),
    .COUT(_12479_),
    .SUM(_12480_));
 sky130_fd_sc_hd__fa_1 _27401_ (.A(_12481_),
    .B(_12482_),
    .CIN(_12483_),
    .COUT(_12484_),
    .SUM(_12485_));
 sky130_fd_sc_hd__fa_1 _27402_ (.A(_12486_),
    .B(_12487_),
    .CIN(_12488_),
    .COUT(_12489_),
    .SUM(_12490_));
 sky130_fd_sc_hd__fa_1 _27403_ (.A(\hash.CA1.k_i2[29] ),
    .B(\hash.CA1.w_i2[29] ),
    .CIN(_12491_),
    .COUT(_12492_),
    .SUM(_12493_));
 sky130_fd_sc_hd__fa_1 _27404_ (.A(\hash.CA1.k_i2[30] ),
    .B(\hash.CA1.w_i2[30] ),
    .CIN(_12494_),
    .COUT(_12495_),
    .SUM(_12496_));
 sky130_fd_sc_hd__fa_1 _27405_ (.A(\hash.CA1.k_i1[1] ),
    .B(\hash.CA1.w_i1[1] ),
    .CIN(_12497_),
    .COUT(_12498_),
    .SUM(_12499_));
 sky130_fd_sc_hd__fa_2 _27406_ (.A(_12500_),
    .B(_12501_),
    .CIN(_12502_),
    .COUT(_12503_),
    .SUM(_12504_));
 sky130_fd_sc_hd__fa_1 _27407_ (.A(_12504_),
    .B(_12499_),
    .CIN(_12505_),
    .COUT(_12506_),
    .SUM(_12507_));
 sky130_fd_sc_hd__fa_1 _27408_ (.A(_12508_),
    .B(_12509_),
    .CIN(_12510_),
    .COUT(_12511_),
    .SUM(_12512_));
 sky130_fd_sc_hd__fa_1 _27409_ (.A(_12513_),
    .B(_12514_),
    .CIN(_12515_),
    .COUT(_12516_),
    .SUM(_12517_));
 sky130_fd_sc_hd__fa_1 _27410_ (.A(_12518_),
    .B(_12519_),
    .CIN(_12520_),
    .COUT(_12521_),
    .SUM(_12522_));
 sky130_fd_sc_hd__fa_1 _27411_ (.A(_12523_),
    .B(_12524_),
    .CIN(_12525_),
    .COUT(_12526_),
    .SUM(_12527_));
 sky130_fd_sc_hd__fa_1 _27412_ (.A(_12528_),
    .B(_12529_),
    .CIN(_12530_),
    .COUT(_12531_),
    .SUM(_12532_));
 sky130_fd_sc_hd__fa_1 _27413_ (.A(_12533_),
    .B(_12534_),
    .CIN(_12535_),
    .COUT(_12536_),
    .SUM(_12537_));
 sky130_fd_sc_hd__fa_1 _27414_ (.A(_12538_),
    .B(_12539_),
    .CIN(_12540_),
    .COUT(_12541_),
    .SUM(_12542_));
 sky130_fd_sc_hd__fa_1 _27415_ (.A(_12543_),
    .B(_12544_),
    .CIN(_12545_),
    .COUT(_12546_),
    .SUM(_12547_));
 sky130_fd_sc_hd__fa_1 _27416_ (.A(_12548_),
    .B(_12549_),
    .CIN(_12550_),
    .COUT(_12551_),
    .SUM(_12552_));
 sky130_fd_sc_hd__fa_1 _27417_ (.A(_12553_),
    .B(_12554_),
    .CIN(_12555_),
    .COUT(_12556_),
    .SUM(_12557_));
 sky130_fd_sc_hd__fa_1 _27418_ (.A(_12558_),
    .B(_12559_),
    .CIN(_12560_),
    .COUT(_12561_),
    .SUM(_12562_));
 sky130_fd_sc_hd__fa_1 _27419_ (.A(_12563_),
    .B(_12564_),
    .CIN(_12565_),
    .COUT(_12566_),
    .SUM(_12567_));
 sky130_fd_sc_hd__fa_1 _27420_ (.A(_12568_),
    .B(_12569_),
    .CIN(_12570_),
    .COUT(_12571_),
    .SUM(_12572_));
 sky130_fd_sc_hd__fa_1 _27421_ (.A(_12573_),
    .B(_12574_),
    .CIN(_12575_),
    .COUT(_12576_),
    .SUM(_12577_));
 sky130_fd_sc_hd__fa_1 _27422_ (.A(_12578_),
    .B(_12579_),
    .CIN(_12580_),
    .COUT(_12581_),
    .SUM(_12582_));
 sky130_fd_sc_hd__fa_1 _27423_ (.A(_12583_),
    .B(_12584_),
    .CIN(_12585_),
    .COUT(_12586_),
    .SUM(_12587_));
 sky130_fd_sc_hd__fa_1 _27424_ (.A(_12588_),
    .B(_12589_),
    .CIN(_06325_),
    .COUT(_12591_),
    .SUM(_12592_));
 sky130_fd_sc_hd__fa_1 _27425_ (.A(_12593_),
    .B(_12594_),
    .CIN(_12595_),
    .COUT(_12596_),
    .SUM(_12597_));
 sky130_fd_sc_hd__fa_1 _27426_ (.A(_12598_),
    .B(_12599_),
    .CIN(_12600_),
    .COUT(_12601_),
    .SUM(_12602_));
 sky130_fd_sc_hd__fa_1 _27427_ (.A(_12603_),
    .B(_12604_),
    .CIN(_12605_),
    .COUT(_12606_),
    .SUM(_12607_));
 sky130_fd_sc_hd__fa_1 _27428_ (.A(_12608_),
    .B(_12609_),
    .CIN(_12610_),
    .COUT(_12611_),
    .SUM(_12612_));
 sky130_fd_sc_hd__fa_1 _27429_ (.A(_12613_),
    .B(_12614_),
    .CIN(_12615_),
    .COUT(_12616_),
    .SUM(_12617_));
 sky130_fd_sc_hd__fa_1 _27430_ (.A(_12618_),
    .B(_12619_),
    .CIN(_12620_),
    .COUT(_12621_),
    .SUM(_12622_));
 sky130_fd_sc_hd__fa_1 _27431_ (.A(_12623_),
    .B(_12624_),
    .CIN(_12625_),
    .COUT(_12626_),
    .SUM(_12627_));
 sky130_fd_sc_hd__fa_1 _27432_ (.A(_12628_),
    .B(_12629_),
    .CIN(_12630_),
    .COUT(_12631_),
    .SUM(_12632_));
 sky130_fd_sc_hd__fa_1 _27433_ (.A(_12633_),
    .B(_12634_),
    .CIN(_12635_),
    .COUT(_12636_),
    .SUM(_12637_));
 sky130_fd_sc_hd__fa_1 _27434_ (.A(_12638_),
    .B(_12639_),
    .CIN(_12640_),
    .COUT(_12641_),
    .SUM(_12642_));
 sky130_fd_sc_hd__fa_1 _27435_ (.A(_12643_),
    .B(_12644_),
    .CIN(_12645_),
    .COUT(_12646_),
    .SUM(_12647_));
 sky130_fd_sc_hd__fa_1 _27436_ (.A(_12648_),
    .B(_12649_),
    .CIN(_12650_),
    .COUT(_12651_),
    .SUM(_12652_));
 sky130_fd_sc_hd__fa_1 _27437_ (.A(\hash.CA1.d[0] ),
    .B(_12653_),
    .CIN(_12654_),
    .COUT(_12655_),
    .SUM(_12656_));
 sky130_fd_sc_hd__fa_1 _27438_ (.A(_12657_),
    .B(_12499_),
    .CIN(_12505_),
    .COUT(_12658_),
    .SUM(_12659_));
 sky130_fd_sc_hd__fa_1 _27439_ (.A(_12660_),
    .B(_12661_),
    .CIN(_12662_),
    .COUT(_12663_),
    .SUM(_12664_));
 sky130_fd_sc_hd__fa_1 _27440_ (.A(_12665_),
    .B(_12666_),
    .CIN(_12667_),
    .COUT(_12668_),
    .SUM(_12669_));
 sky130_fd_sc_hd__fa_1 _27441_ (.A(_12670_),
    .B(_12669_),
    .CIN(_12671_),
    .COUT(_12672_),
    .SUM(_12673_));
 sky130_fd_sc_hd__fa_1 _27442_ (.A(_12514_),
    .B(_12674_),
    .CIN(_12515_),
    .COUT(_12675_),
    .SUM(_12676_));
 sky130_fd_sc_hd__fa_1 _27443_ (.A(_12668_),
    .B(_12676_),
    .CIN(_12513_),
    .COUT(_12677_),
    .SUM(_12678_));
 sky130_fd_sc_hd__fa_1 _27444_ (.A(_12519_),
    .B(_12679_),
    .CIN(_12520_),
    .COUT(_12680_),
    .SUM(_12681_));
 sky130_fd_sc_hd__fa_1 _27445_ (.A(_12675_),
    .B(_12681_),
    .CIN(_12518_),
    .COUT(_12682_),
    .SUM(_12683_));
 sky130_fd_sc_hd__fa_1 _27446_ (.A(_12524_),
    .B(_12684_),
    .CIN(_12525_),
    .COUT(_12685_),
    .SUM(_12686_));
 sky130_fd_sc_hd__fa_1 _27447_ (.A(_12680_),
    .B(_12687_),
    .CIN(_12688_),
    .COUT(_12689_),
    .SUM(_12690_));
 sky130_fd_sc_hd__fa_1 _27448_ (.A(_12691_),
    .B(_12692_),
    .CIN(_12693_),
    .COUT(_12694_),
    .SUM(_12695_));
 sky130_fd_sc_hd__fa_1 _27449_ (.A(_12696_),
    .B(_12695_),
    .CIN(_12697_),
    .COUT(_12698_),
    .SUM(_12699_));
 sky130_fd_sc_hd__fa_1 _27450_ (.A(_12700_),
    .B(_12701_),
    .CIN(_12702_),
    .COUT(_12703_),
    .SUM(_12704_));
 sky130_fd_sc_hd__fa_1 _27451_ (.A(_12694_),
    .B(_12704_),
    .CIN(_12705_),
    .COUT(_12706_),
    .SUM(_12707_));
 sky130_fd_sc_hd__fa_1 _27452_ (.A(_12539_),
    .B(_12708_),
    .CIN(_12540_),
    .COUT(_12709_),
    .SUM(_12710_));
 sky130_fd_sc_hd__fa_1 _27453_ (.A(_12703_),
    .B(_12710_),
    .CIN(_12538_),
    .COUT(_12711_),
    .SUM(_12712_));
 sky130_fd_sc_hd__fa_1 _27454_ (.A(_12713_),
    .B(_12714_),
    .CIN(_12715_),
    .COUT(_12716_),
    .SUM(_12717_));
 sky130_fd_sc_hd__fa_1 _27455_ (.A(_12720_),
    .B(_12719_),
    .CIN(_12718_),
    .COUT(_12721_),
    .SUM(_12722_));
 sky130_fd_sc_hd__fa_1 _27456_ (.A(_12549_),
    .B(_12723_),
    .CIN(_12550_),
    .COUT(_12724_),
    .SUM(_12725_));
 sky130_fd_sc_hd__fa_1 _27457_ (.A(_12726_),
    .B(_12728_),
    .CIN(_12727_),
    .COUT(_12729_),
    .SUM(_12730_));
 sky130_fd_sc_hd__fa_1 _27458_ (.A(_12731_),
    .B(_12732_),
    .CIN(_12733_),
    .COUT(_12734_),
    .SUM(_12735_));
 sky130_fd_sc_hd__fa_1 _27459_ (.A(_12736_),
    .B(_12735_),
    .CIN(_12737_),
    .COUT(_12738_),
    .SUM(_12739_));
 sky130_fd_sc_hd__fa_1 _27460_ (.A(_12559_),
    .B(_06747_),
    .CIN(_12560_),
    .COUT(_12741_),
    .SUM(_12742_));
 sky130_fd_sc_hd__fa_1 _27461_ (.A(_12734_),
    .B(_12742_),
    .CIN(_12743_),
    .COUT(_12744_),
    .SUM(_12745_));
 sky130_fd_sc_hd__fa_1 _27462_ (.A(_12564_),
    .B(_12746_),
    .CIN(_12565_),
    .COUT(_12747_),
    .SUM(_12748_));
 sky130_fd_sc_hd__fa_1 _27463_ (.A(_12741_),
    .B(_12748_),
    .CIN(_12749_),
    .COUT(_12750_),
    .SUM(_12751_));
 sky130_fd_sc_hd__fa_1 _27464_ (.A(_12569_),
    .B(_12752_),
    .CIN(_12570_),
    .COUT(_12753_),
    .SUM(_12754_));
 sky130_fd_sc_hd__fa_1 _27465_ (.A(_12747_),
    .B(_12755_),
    .CIN(_12756_),
    .COUT(_12757_),
    .SUM(_12758_));
 sky130_fd_sc_hd__fa_1 _27466_ (.A(_12574_),
    .B(_12759_),
    .CIN(_12575_),
    .COUT(_12760_),
    .SUM(_12761_));
 sky130_fd_sc_hd__fa_1 _27467_ (.A(_12762_),
    .B(_12763_),
    .CIN(_12764_),
    .COUT(_12765_),
    .SUM(_12766_));
 sky130_fd_sc_hd__fa_1 _27468_ (.A(_12579_),
    .B(_12767_),
    .CIN(_12580_),
    .COUT(_12768_),
    .SUM(_12769_));
 sky130_fd_sc_hd__fa_1 _27469_ (.A(_12770_),
    .B(_12769_),
    .CIN(_12771_),
    .COUT(_12772_),
    .SUM(_12773_));
 sky130_fd_sc_hd__fa_1 _27470_ (.A(_12584_),
    .B(_12774_),
    .CIN(_12585_),
    .COUT(_12775_),
    .SUM(_12776_));
 sky130_fd_sc_hd__fa_1 _27471_ (.A(_12768_),
    .B(_12776_),
    .CIN(_12777_),
    .COUT(_12778_),
    .SUM(_12779_));
 sky130_fd_sc_hd__fa_1 _27472_ (.A(_12589_),
    .B(_12780_),
    .CIN(_06325_),
    .COUT(_12781_),
    .SUM(_12782_));
 sky130_fd_sc_hd__fa_1 _27473_ (.A(_12775_),
    .B(_12782_),
    .CIN(_12783_),
    .COUT(_12784_),
    .SUM(_12785_));
 sky130_fd_sc_hd__fa_1 _27474_ (.A(_12594_),
    .B(_12786_),
    .CIN(_12595_),
    .COUT(_12787_),
    .SUM(_12788_));
 sky130_fd_sc_hd__fa_1 _27475_ (.A(_12781_),
    .B(_12788_),
    .CIN(_12789_),
    .COUT(_12790_),
    .SUM(_12791_));
 sky130_fd_sc_hd__fa_1 _27476_ (.A(_12792_),
    .B(_12793_),
    .CIN(_12794_),
    .COUT(_12795_),
    .SUM(_12796_));
 sky130_fd_sc_hd__fa_1 _27477_ (.A(_12787_),
    .B(_12797_),
    .CIN(_12798_),
    .COUT(_12799_),
    .SUM(_12800_));
 sky130_fd_sc_hd__fa_1 _27478_ (.A(_12801_),
    .B(_12802_),
    .CIN(_12803_),
    .COUT(_12804_),
    .SUM(_12805_));
 sky130_fd_sc_hd__fa_1 _27479_ (.A(_12806_),
    .B(_12805_),
    .CIN(_12807_),
    .COUT(_12808_),
    .SUM(_12809_));
 sky130_fd_sc_hd__fa_1 _27480_ (.A(_12609_),
    .B(_12810_),
    .CIN(_12610_),
    .COUT(_12811_),
    .SUM(_12812_));
 sky130_fd_sc_hd__fa_1 _27481_ (.A(_12804_),
    .B(_12813_),
    .CIN(_12814_),
    .COUT(_12815_),
    .SUM(_12816_));
 sky130_fd_sc_hd__fa_1 _27482_ (.A(_12817_),
    .B(_12818_),
    .CIN(_12819_),
    .COUT(_12820_),
    .SUM(_12821_));
 sky130_fd_sc_hd__fa_1 _27483_ (.A(_12822_),
    .B(_12821_),
    .CIN(_12823_),
    .COUT(_12824_),
    .SUM(_12825_));
 sky130_fd_sc_hd__fa_1 _27484_ (.A(_12619_),
    .B(_12826_),
    .CIN(_12620_),
    .COUT(_12827_),
    .SUM(_12828_));
 sky130_fd_sc_hd__fa_1 _27485_ (.A(_12820_),
    .B(_12829_),
    .CIN(_12830_),
    .COUT(_12831_),
    .SUM(_12832_));
 sky130_fd_sc_hd__fa_1 _27486_ (.A(_12833_),
    .B(_12834_),
    .CIN(_12835_),
    .COUT(_12836_),
    .SUM(_12837_));
 sky130_fd_sc_hd__fa_1 _27487_ (.A(_12838_),
    .B(_12837_),
    .CIN(_12839_),
    .COUT(_12840_),
    .SUM(_12841_));
 sky130_fd_sc_hd__fa_1 _27488_ (.A(_12629_),
    .B(_12842_),
    .CIN(_12630_),
    .COUT(_12843_),
    .SUM(_12844_));
 sky130_fd_sc_hd__fa_1 _27489_ (.A(_12836_),
    .B(_12844_),
    .CIN(_12845_),
    .COUT(_12846_),
    .SUM(_12847_));
 sky130_fd_sc_hd__fa_1 _27490_ (.A(_12848_),
    .B(_12849_),
    .CIN(_12850_),
    .COUT(_12851_),
    .SUM(_12852_));
 sky130_fd_sc_hd__fa_1 _27491_ (.A(_12843_),
    .B(_12852_),
    .CIN(_12853_),
    .COUT(_12854_),
    .SUM(_12855_));
 sky130_fd_sc_hd__fa_1 _27492_ (.A(_12856_),
    .B(_12857_),
    .CIN(_12858_),
    .COUT(_12859_),
    .SUM(_12860_));
 sky130_fd_sc_hd__fa_1 _27493_ (.A(_12851_),
    .B(_12860_),
    .CIN(_12861_),
    .COUT(_12862_),
    .SUM(_12863_));
 sky130_fd_sc_hd__fa_1 _27494_ (.A(_12644_),
    .B(_12864_),
    .CIN(_12645_),
    .COUT(_12865_),
    .SUM(_12866_));
 sky130_fd_sc_hd__fa_1 _27495_ (.A(_12859_),
    .B(_12866_),
    .CIN(_12867_),
    .COUT(_12868_),
    .SUM(_12869_));
 sky130_fd_sc_hd__fa_1 _27496_ (.A(_12870_),
    .B(_12871_),
    .CIN(_12872_),
    .COUT(_12873_),
    .SUM(_12874_));
 sky130_fd_sc_hd__fa_1 _27497_ (.A(_12875_),
    .B(_12876_),
    .CIN(_12648_),
    .COUT(_12877_),
    .SUM(_12878_));
 sky130_fd_sc_hd__fa_2 _27498_ (.A(_12881_),
    .B(_12880_),
    .CIN(_12879_),
    .COUT(_12882_),
    .SUM(_12883_));
 sky130_fd_sc_hd__fa_1 _27499_ (.A(_12884_),
    .B(_12663_),
    .CIN(_12673_),
    .COUT(_12885_),
    .SUM(_12886_));
 sky130_fd_sc_hd__fa_1 _27500_ (.A(_12653_),
    .B(_12887_),
    .CIN(_12654_),
    .COUT(_12888_),
    .SUM(\hash.CA1.p3[0] ));
 sky130_fd_sc_hd__fa_1 _27501_ (.A(_12889_),
    .B(_12890_),
    .CIN(_12891_),
    .COUT(_12892_),
    .SUM(_12893_));
 sky130_fd_sc_hd__fa_1 _27502_ (.A(_00721_),
    .B(_12894_),
    .CIN(_12895_),
    .COUT(_12896_),
    .SUM(_12897_));
 sky130_fd_sc_hd__ha_4 _27503_ (.A(_00656_),
    .B(_12900_),
    .COUT(_12901_),
    .SUM(_00657_));
 sky130_fd_sc_hd__ha_4 _27504_ (.A(_00656_),
    .B(\count_hash2[2] ),
    .COUT(_12902_),
    .SUM(_12903_));
 sky130_fd_sc_hd__ha_4 _27505_ (.A(\count_hash2[1] ),
    .B(_12900_),
    .COUT(_12904_),
    .SUM(_12905_));
 sky130_fd_sc_hd__ha_4 _27506_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_12906_),
    .SUM(_12907_));
 sky130_fd_sc_hd__ha_4 _27507_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_12908_),
    .SUM(_12909_));
 sky130_fd_sc_hd__ha_4 _27508_ (.A(_00654_),
    .B(_12910_),
    .COUT(_12911_),
    .SUM(_00655_));
 sky130_fd_sc_hd__ha_4 _27509_ (.A(_00654_),
    .B(\count_hash1[2] ),
    .COUT(_12912_),
    .SUM(_12913_));
 sky130_fd_sc_hd__ha_1 _27510_ (.A(_00654_),
    .B(\count_hash1[2] ),
    .COUT(_12914_),
    .SUM(_12915_));
 sky130_fd_sc_hd__ha_4 _27511_ (.A(\count_hash1[1] ),
    .B(_12910_),
    .COUT(_12916_),
    .SUM(_12917_));
 sky130_fd_sc_hd__ha_4 _27512_ (.A(\count_hash1[1] ),
    .B(\count_hash1[2] ),
    .COUT(_12918_),
    .SUM(_12919_));
 sky130_fd_sc_hd__ha_4 _27513_ (.A(\count_hash1[1] ),
    .B(\count_hash1[2] ),
    .COUT(_12920_),
    .SUM(_12921_));
 sky130_fd_sc_hd__ha_4 _27514_ (.A(\hash.CA2.p3[0] ),
    .B(\hash.CA2.p1[0] ),
    .COUT(_12080_),
    .SUM(_12922_));
 sky130_fd_sc_hd__ha_4 _27515_ (.A(\hash.CA2.p1[2] ),
    .B(\hash.CA2.p3[2] ),
    .COUT(_12923_),
    .SUM(_12924_));
 sky130_fd_sc_hd__ha_1 _27516_ (.A(\hash.CA2.p1[1] ),
    .B(\hash.CA2.p3[1] ),
    .COUT(_12925_),
    .SUM(_12926_));
 sky130_fd_sc_hd__ha_4 _27517_ (.A(\hash.CA2.p1[7] ),
    .B(\hash.CA2.p3[7] ),
    .COUT(_12927_),
    .SUM(_12928_));
 sky130_fd_sc_hd__ha_2 _27518_ (.A(\hash.CA2.p1[6] ),
    .B(\hash.CA2.p3[6] ),
    .COUT(_12929_),
    .SUM(_12930_));
 sky130_fd_sc_hd__ha_1 _27519_ (.A(\hash.CA2.p1[5] ),
    .B(\hash.CA2.p3[5] ),
    .COUT(_12931_),
    .SUM(_12932_));
 sky130_fd_sc_hd__ha_1 _27520_ (.A(\hash.CA2.p1[4] ),
    .B(\hash.CA2.p3[4] ),
    .COUT(_12933_),
    .SUM(_12934_));
 sky130_fd_sc_hd__ha_4 _27521_ (.A(\hash.CA2.p1[3] ),
    .B(\hash.CA2.p3[3] ),
    .COUT(_12935_),
    .SUM(_12936_));
 sky130_fd_sc_hd__ha_1 _27522_ (.A(\hash.CA2.p1[9] ),
    .B(\hash.CA2.p3[9] ),
    .COUT(_12937_),
    .SUM(_12938_));
 sky130_fd_sc_hd__ha_4 _27523_ (.A(\hash.CA2.p1[8] ),
    .B(\hash.CA2.p3[8] ),
    .COUT(_12939_),
    .SUM(_12940_));
 sky130_fd_sc_hd__ha_1 _27524_ (.A(\hash.CA2.p1[10] ),
    .B(\hash.CA2.p3[10] ),
    .COUT(_12941_),
    .SUM(_12942_));
 sky130_fd_sc_hd__ha_4 _27525_ (.A(\hash.CA2.p1[11] ),
    .B(\hash.CA2.p3[11] ),
    .COUT(_12943_),
    .SUM(_12944_));
 sky130_fd_sc_hd__ha_4 _27526_ (.A(\hash.CA2.p1[13] ),
    .B(\hash.CA2.p3[13] ),
    .COUT(_12945_),
    .SUM(_12946_));
 sky130_fd_sc_hd__ha_4 _27527_ (.A(\hash.CA2.p1[12] ),
    .B(\hash.CA2.p3[12] ),
    .COUT(_12947_),
    .SUM(_12948_));
 sky130_fd_sc_hd__ha_1 _27528_ (.A(\hash.CA2.p1[15] ),
    .B(\hash.CA2.p3[15] ),
    .COUT(_12949_),
    .SUM(_12950_));
 sky130_fd_sc_hd__ha_1 _27529_ (.A(\hash.CA2.p1[14] ),
    .B(\hash.CA2.p3[14] ),
    .COUT(_12951_),
    .SUM(_12952_));
 sky130_fd_sc_hd__ha_4 _27530_ (.A(\hash.CA2.p1[16] ),
    .B(\hash.CA2.p3[16] ),
    .COUT(_12953_),
    .SUM(_12954_));
 sky130_fd_sc_hd__ha_2 _27531_ (.A(\hash.CA2.p1[17] ),
    .B(\hash.CA2.p3[17] ),
    .COUT(_12955_),
    .SUM(_12956_));
 sky130_fd_sc_hd__ha_1 _27532_ (.A(\hash.CA2.p1[18] ),
    .B(\hash.CA2.p3[18] ),
    .COUT(_12957_),
    .SUM(_12958_));
 sky130_fd_sc_hd__ha_4 _27533_ (.A(\hash.CA2.p1[21] ),
    .B(\hash.CA2.p3[21] ),
    .COUT(_12959_),
    .SUM(_12960_));
 sky130_fd_sc_hd__ha_4 _27534_ (.A(\hash.CA2.p1[20] ),
    .B(\hash.CA2.p3[20] ),
    .COUT(_12961_),
    .SUM(_12962_));
 sky130_fd_sc_hd__ha_4 _27535_ (.A(\hash.CA2.p1[19] ),
    .B(\hash.CA2.p3[19] ),
    .COUT(_12963_),
    .SUM(_12964_));
 sky130_fd_sc_hd__ha_4 _27536_ (.A(\hash.CA2.p1[22] ),
    .B(\hash.CA2.p3[22] ),
    .COUT(_12965_),
    .SUM(_12966_));
 sky130_fd_sc_hd__ha_2 _27537_ (.A(\hash.CA2.p1[24] ),
    .B(\hash.CA2.p3[24] ),
    .COUT(_12967_),
    .SUM(_12968_));
 sky130_fd_sc_hd__ha_4 _27538_ (.A(\hash.CA2.p1[23] ),
    .B(\hash.CA2.p3[23] ),
    .COUT(_12969_),
    .SUM(_12970_));
 sky130_fd_sc_hd__ha_4 _27539_ (.A(\hash.CA2.p1[25] ),
    .B(\hash.CA2.p3[25] ),
    .COUT(_12971_),
    .SUM(_12972_));
 sky130_fd_sc_hd__ha_4 _27540_ (.A(\hash.CA2.p1[27] ),
    .B(\hash.CA2.p3[27] ),
    .COUT(_12973_),
    .SUM(_12974_));
 sky130_fd_sc_hd__ha_4 _27541_ (.A(\hash.CA2.p1[26] ),
    .B(\hash.CA2.p3[26] ),
    .COUT(_12975_),
    .SUM(_12976_));
 sky130_fd_sc_hd__ha_4 _27542_ (.A(\hash.CA2.p1[28] ),
    .B(\hash.CA2.p3[28] ),
    .COUT(_12977_),
    .SUM(_12978_));
 sky130_fd_sc_hd__ha_4 _27543_ (.A(\hash.CA2.p1[29] ),
    .B(\hash.CA2.p3[29] ),
    .COUT(_12979_),
    .SUM(_12980_));
 sky130_fd_sc_hd__ha_1 _27544_ (.A(\hash.CA2.p1[30] ),
    .B(\hash.CA2.p3[30] ),
    .COUT(_12981_),
    .SUM(_12982_));
 sky130_fd_sc_hd__ha_1 _27545_ (.A(_12983_),
    .B(_12984_),
    .COUT(_12985_),
    .SUM(_12986_));
 sky130_fd_sc_hd__ha_1 _27546_ (.A(_12985_),
    .B(_12987_),
    .COUT(_12988_),
    .SUM(_12989_));
 sky130_fd_sc_hd__ha_1 _27547_ (.A(_12990_),
    .B(_12991_),
    .COUT(_12992_),
    .SUM(_12993_));
 sky130_fd_sc_hd__ha_1 _27548_ (.A(_12994_),
    .B(_12995_),
    .COUT(_12996_),
    .SUM(_12997_));
 sky130_fd_sc_hd__ha_1 _27549_ (.A(_12998_),
    .B(_12999_),
    .COUT(_13000_),
    .SUM(_13001_));
 sky130_fd_sc_hd__ha_1 _27550_ (.A(_13002_),
    .B(_13003_),
    .COUT(_13004_),
    .SUM(_13005_));
 sky130_fd_sc_hd__ha_1 _27551_ (.A(_13006_),
    .B(_13007_),
    .COUT(_13008_),
    .SUM(_13009_));
 sky130_fd_sc_hd__ha_4 _27552_ (.A(_13010_),
    .B(_13011_),
    .COUT(_13012_),
    .SUM(_13013_));
 sky130_fd_sc_hd__ha_4 _27553_ (.A(_13014_),
    .B(_13015_),
    .COUT(_13016_),
    .SUM(_13017_));
 sky130_fd_sc_hd__ha_4 _27554_ (.A(_13018_),
    .B(_13019_),
    .COUT(_13020_),
    .SUM(_13021_));
 sky130_fd_sc_hd__ha_4 _27555_ (.A(_13022_),
    .B(_13023_),
    .COUT(_13024_),
    .SUM(_13025_));
 sky130_fd_sc_hd__ha_4 _27556_ (.A(_13026_),
    .B(_13027_),
    .COUT(_13028_),
    .SUM(_13029_));
 sky130_fd_sc_hd__ha_1 _27557_ (.A(_13030_),
    .B(_13031_),
    .COUT(_13032_),
    .SUM(_13033_));
 sky130_fd_sc_hd__ha_1 _27558_ (.A(_13034_),
    .B(_13035_),
    .COUT(_13036_),
    .SUM(_13037_));
 sky130_fd_sc_hd__ha_1 _27559_ (.A(_13038_),
    .B(_13039_),
    .COUT(_13040_),
    .SUM(_13041_));
 sky130_fd_sc_hd__ha_1 _27560_ (.A(_13042_),
    .B(_13043_),
    .COUT(_13044_),
    .SUM(_13045_));
 sky130_fd_sc_hd__ha_1 _27561_ (.A(_13046_),
    .B(_13047_),
    .COUT(_13048_),
    .SUM(_13049_));
 sky130_fd_sc_hd__ha_1 _27562_ (.A(_13050_),
    .B(_13051_),
    .COUT(_13052_),
    .SUM(_13053_));
 sky130_fd_sc_hd__ha_1 _27563_ (.A(_13054_),
    .B(_13055_),
    .COUT(_13056_),
    .SUM(_13057_));
 sky130_fd_sc_hd__ha_1 _27564_ (.A(_13058_),
    .B(_13059_),
    .COUT(_13060_),
    .SUM(_13061_));
 sky130_fd_sc_hd__ha_4 _27565_ (.A(_13062_),
    .B(_13063_),
    .COUT(_13064_),
    .SUM(_13065_));
 sky130_fd_sc_hd__ha_1 _27566_ (.A(_13066_),
    .B(_13067_),
    .COUT(_13068_),
    .SUM(_13069_));
 sky130_fd_sc_hd__ha_4 _27567_ (.A(_13070_),
    .B(_13071_),
    .COUT(_13072_),
    .SUM(_13073_));
 sky130_fd_sc_hd__ha_2 _27568_ (.A(_13074_),
    .B(_13075_),
    .COUT(_13076_),
    .SUM(_13077_));
 sky130_fd_sc_hd__ha_1 _27569_ (.A(_13078_),
    .B(_13079_),
    .COUT(_13080_),
    .SUM(_13081_));
 sky130_fd_sc_hd__ha_4 _27570_ (.A(_13082_),
    .B(_13083_),
    .COUT(_13084_),
    .SUM(_13085_));
 sky130_fd_sc_hd__ha_4 _27571_ (.A(_13086_),
    .B(_13087_),
    .COUT(_13088_),
    .SUM(_13089_));
 sky130_fd_sc_hd__ha_4 _27572_ (.A(_13090_),
    .B(_13091_),
    .COUT(_13092_),
    .SUM(_13093_));
 sky130_fd_sc_hd__ha_4 _27573_ (.A(_13094_),
    .B(_13095_),
    .COUT(_13096_),
    .SUM(_13097_));
 sky130_fd_sc_hd__ha_4 _27574_ (.A(_13098_),
    .B(_13099_),
    .COUT(_13100_),
    .SUM(_13101_));
 sky130_fd_sc_hd__ha_4 _27575_ (.A(_13102_),
    .B(_13103_),
    .COUT(_13104_),
    .SUM(_13105_));
 sky130_fd_sc_hd__ha_1 _27576_ (.A(_13106_),
    .B(_13107_),
    .COUT(_13108_),
    .SUM(_13109_));
 sky130_fd_sc_hd__ha_2 _27577_ (.A(_13108_),
    .B(_13110_),
    .COUT(_13111_),
    .SUM(_13112_));
 sky130_fd_sc_hd__ha_1 _27578_ (.A(_13113_),
    .B(_13114_),
    .COUT(_13115_),
    .SUM(_13116_));
 sky130_fd_sc_hd__ha_2 _27579_ (.A(_13117_),
    .B(_13118_),
    .COUT(_13119_),
    .SUM(_13120_));
 sky130_fd_sc_hd__ha_1 _27580_ (.A(_13121_),
    .B(_13122_),
    .COUT(_13123_),
    .SUM(_13124_));
 sky130_fd_sc_hd__ha_2 _27581_ (.A(_13125_),
    .B(_13126_),
    .COUT(_13127_),
    .SUM(_13128_));
 sky130_fd_sc_hd__ha_1 _27582_ (.A(_13129_),
    .B(_13130_),
    .COUT(_13131_),
    .SUM(_13132_));
 sky130_fd_sc_hd__ha_4 _27583_ (.A(_13133_),
    .B(_13134_),
    .COUT(_13135_),
    .SUM(_13136_));
 sky130_fd_sc_hd__ha_4 _27584_ (.A(_13137_),
    .B(_13138_),
    .COUT(_13139_),
    .SUM(_13140_));
 sky130_fd_sc_hd__ha_4 _27585_ (.A(_13141_),
    .B(_13142_),
    .COUT(_13143_),
    .SUM(_13144_));
 sky130_fd_sc_hd__ha_4 _27586_ (.A(_13145_),
    .B(_13146_),
    .COUT(_13147_),
    .SUM(_13148_));
 sky130_fd_sc_hd__ha_4 _27587_ (.A(_13149_),
    .B(_13150_),
    .COUT(_13151_),
    .SUM(_13152_));
 sky130_fd_sc_hd__ha_4 _27588_ (.A(_13153_),
    .B(_13154_),
    .COUT(_13155_),
    .SUM(_13156_));
 sky130_fd_sc_hd__ha_1 _27589_ (.A(_13157_),
    .B(_13158_),
    .COUT(_13159_),
    .SUM(_13160_));
 sky130_fd_sc_hd__ha_1 _27590_ (.A(_13161_),
    .B(_13162_),
    .COUT(_13163_),
    .SUM(_13164_));
 sky130_fd_sc_hd__ha_1 _27591_ (.A(_13165_),
    .B(_13166_),
    .COUT(_13167_),
    .SUM(_13168_));
 sky130_fd_sc_hd__ha_1 _27592_ (.A(_13169_),
    .B(_13170_),
    .COUT(_13171_),
    .SUM(_13172_));
 sky130_fd_sc_hd__ha_4 _27593_ (.A(_13173_),
    .B(_13174_),
    .COUT(_13175_),
    .SUM(_13176_));
 sky130_fd_sc_hd__ha_4 _27594_ (.A(_13177_),
    .B(_13178_),
    .COUT(_13179_),
    .SUM(_13180_));
 sky130_fd_sc_hd__ha_4 _27595_ (.A(_13181_),
    .B(_13182_),
    .COUT(_13183_),
    .SUM(_13184_));
 sky130_fd_sc_hd__ha_1 _27596_ (.A(_13185_),
    .B(_13186_),
    .COUT(_13187_),
    .SUM(_13188_));
 sky130_fd_sc_hd__ha_1 _27597_ (.A(_13189_),
    .B(_13190_),
    .COUT(_13191_),
    .SUM(_13192_));
 sky130_fd_sc_hd__ha_4 _27598_ (.A(_13193_),
    .B(_13194_),
    .COUT(_13195_),
    .SUM(_13196_));
 sky130_fd_sc_hd__ha_4 _27599_ (.A(_13197_),
    .B(_13198_),
    .COUT(_13199_),
    .SUM(_13200_));
 sky130_fd_sc_hd__ha_1 _27600_ (.A(_13201_),
    .B(_13202_),
    .COUT(_13203_),
    .SUM(_13204_));
 sky130_fd_sc_hd__ha_1 _27601_ (.A(_13205_),
    .B(_13206_),
    .COUT(_13207_),
    .SUM(_13208_));
 sky130_fd_sc_hd__ha_4 _27602_ (.A(_13209_),
    .B(_13210_),
    .COUT(_13211_),
    .SUM(_13212_));
 sky130_fd_sc_hd__ha_4 _27603_ (.A(_13213_),
    .B(_13214_),
    .COUT(_13215_),
    .SUM(_13216_));
 sky130_fd_sc_hd__ha_1 _27604_ (.A(_13217_),
    .B(_13218_),
    .COUT(_13219_),
    .SUM(_13220_));
 sky130_fd_sc_hd__ha_1 _27605_ (.A(_13221_),
    .B(_13222_),
    .COUT(_13223_),
    .SUM(_13224_));
 sky130_fd_sc_hd__ha_1 _27606_ (.A(_13225_),
    .B(_13226_),
    .COUT(_13227_),
    .SUM(_13228_));
 sky130_fd_sc_hd__ha_4 _27607_ (.A(_13229_),
    .B(_13230_),
    .COUT(_13231_),
    .SUM(_13232_));
 sky130_fd_sc_hd__ha_1 _27608_ (.A(\hash.CA2.p4[0] ),
    .B(_13233_),
    .COUT(_13234_),
    .SUM(_13235_));
 sky130_fd_sc_hd__ha_1 _27609_ (.A(_13237_),
    .B(_13236_),
    .COUT(_13238_),
    .SUM(_13239_));
 sky130_fd_sc_hd__ha_1 _27610_ (.A(_13234_),
    .B(_12095_),
    .COUT(_13240_),
    .SUM(_13241_));
 sky130_fd_sc_hd__ha_4 _27611_ (.A(_13242_),
    .B(_13243_),
    .COUT(_13244_),
    .SUM(_13245_));
 sky130_fd_sc_hd__ha_1 _27612_ (.A(_12094_),
    .B(_12104_),
    .COUT(_13247_),
    .SUM(_13248_));
 sky130_fd_sc_hd__ha_1 _27613_ (.A(_13249_),
    .B(_13250_),
    .COUT(_13251_),
    .SUM(_13252_));
 sky130_fd_sc_hd__ha_1 _27614_ (.A(_12103_),
    .B(_12118_),
    .COUT(_13254_),
    .SUM(_13255_));
 sky130_fd_sc_hd__ha_1 _27615_ (.A(_13256_),
    .B(_13257_),
    .COUT(_13258_),
    .SUM(_13259_));
 sky130_fd_sc_hd__ha_4 _27616_ (.A(_12117_),
    .B(_12127_),
    .COUT(_13261_),
    .SUM(_13262_));
 sky130_fd_sc_hd__ha_4 _27617_ (.A(_13263_),
    .B(_13264_),
    .COUT(_13265_),
    .SUM(_13266_));
 sky130_fd_sc_hd__ha_1 _27618_ (.A(_12126_),
    .B(_12136_),
    .COUT(_13268_),
    .SUM(_13269_));
 sky130_fd_sc_hd__ha_1 _27619_ (.A(_13270_),
    .B(_13271_),
    .COUT(_13272_),
    .SUM(_13273_));
 sky130_fd_sc_hd__ha_2 _27620_ (.A(_12135_),
    .B(_12145_),
    .COUT(_13275_),
    .SUM(_13276_));
 sky130_fd_sc_hd__ha_1 _27621_ (.A(_13277_),
    .B(_13278_),
    .COUT(_13279_),
    .SUM(_13280_));
 sky130_fd_sc_hd__ha_4 _27622_ (.A(_12144_),
    .B(_12154_),
    .COUT(_13282_),
    .SUM(_13283_));
 sky130_fd_sc_hd__ha_1 _27623_ (.A(_13284_),
    .B(_13285_),
    .COUT(_13286_),
    .SUM(_13287_));
 sky130_fd_sc_hd__ha_4 _27624_ (.A(_12163_),
    .B(_12153_),
    .COUT(_13289_),
    .SUM(_13290_));
 sky130_fd_sc_hd__ha_1 _27625_ (.A(_13291_),
    .B(_13292_),
    .COUT(_13293_),
    .SUM(_13294_));
 sky130_fd_sc_hd__ha_4 _27626_ (.A(_12162_),
    .B(_12172_),
    .COUT(_13296_),
    .SUM(_13297_));
 sky130_fd_sc_hd__ha_4 _27627_ (.A(_13298_),
    .B(_13299_),
    .COUT(_13300_),
    .SUM(_13301_));
 sky130_fd_sc_hd__ha_1 _27628_ (.A(_12171_),
    .B(_12181_),
    .COUT(_13303_),
    .SUM(_13304_));
 sky130_fd_sc_hd__ha_4 _27629_ (.A(_13305_),
    .B(_13306_),
    .COUT(_13307_),
    .SUM(_13308_));
 sky130_fd_sc_hd__ha_4 _27630_ (.A(_12180_),
    .B(_12190_),
    .COUT(_13310_),
    .SUM(_13311_));
 sky130_fd_sc_hd__ha_1 _27631_ (.A(_13312_),
    .B(_13313_),
    .COUT(_13314_),
    .SUM(_13315_));
 sky130_fd_sc_hd__ha_4 _27632_ (.A(_12189_),
    .B(_12199_),
    .COUT(_13317_),
    .SUM(_13318_));
 sky130_fd_sc_hd__ha_2 _27633_ (.A(_13319_),
    .B(_13320_),
    .COUT(_13321_),
    .SUM(_13322_));
 sky130_fd_sc_hd__ha_4 _27634_ (.A(_12198_),
    .B(_12208_),
    .COUT(_13324_),
    .SUM(_13325_));
 sky130_fd_sc_hd__ha_4 _27635_ (.A(_13326_),
    .B(_13327_),
    .COUT(_13328_),
    .SUM(_13329_));
 sky130_fd_sc_hd__ha_4 _27636_ (.A(_12207_),
    .B(_12217_),
    .COUT(_13331_),
    .SUM(_13332_));
 sky130_fd_sc_hd__ha_2 _27637_ (.A(_13333_),
    .B(_13334_),
    .COUT(_13335_),
    .SUM(_13336_));
 sky130_fd_sc_hd__ha_4 _27638_ (.A(_12216_),
    .B(_12226_),
    .COUT(_13338_),
    .SUM(_13339_));
 sky130_fd_sc_hd__ha_2 _27639_ (.A(_13340_),
    .B(_13341_),
    .COUT(_13342_),
    .SUM(_13343_));
 sky130_fd_sc_hd__ha_4 _27640_ (.A(_12225_),
    .B(_12235_),
    .COUT(_13345_),
    .SUM(_13346_));
 sky130_fd_sc_hd__ha_1 _27641_ (.A(_13347_),
    .B(_13348_),
    .COUT(_13349_),
    .SUM(_13350_));
 sky130_fd_sc_hd__ha_4 _27642_ (.A(_12234_),
    .B(_12244_),
    .COUT(_13352_),
    .SUM(_13353_));
 sky130_fd_sc_hd__ha_1 _27643_ (.A(_13354_),
    .B(_13355_),
    .COUT(_13356_),
    .SUM(_13357_));
 sky130_fd_sc_hd__ha_4 _27644_ (.A(_12243_),
    .B(_12253_),
    .COUT(_13359_),
    .SUM(_13360_));
 sky130_fd_sc_hd__ha_4 _27645_ (.A(_13361_),
    .B(_13362_),
    .COUT(_13363_),
    .SUM(_13364_));
 sky130_fd_sc_hd__ha_1 _27646_ (.A(_12252_),
    .B(_12262_),
    .COUT(_13366_),
    .SUM(_13367_));
 sky130_fd_sc_hd__ha_4 _27647_ (.A(_13368_),
    .B(_13369_),
    .COUT(_13370_),
    .SUM(_13371_));
 sky130_fd_sc_hd__ha_4 _27648_ (.A(_12261_),
    .B(_12271_),
    .COUT(_13373_),
    .SUM(_13374_));
 sky130_fd_sc_hd__ha_1 _27649_ (.A(_13375_),
    .B(_13376_),
    .COUT(_13377_),
    .SUM(_13378_));
 sky130_fd_sc_hd__ha_4 _27650_ (.A(_12270_),
    .B(_12280_),
    .COUT(_13380_),
    .SUM(_13381_));
 sky130_fd_sc_hd__ha_2 _27651_ (.A(_13382_),
    .B(_13383_),
    .COUT(_13384_),
    .SUM(_13385_));
 sky130_fd_sc_hd__ha_4 _27652_ (.A(_12279_),
    .B(_12289_),
    .COUT(_13387_),
    .SUM(_13388_));
 sky130_fd_sc_hd__ha_1 _27653_ (.A(_13389_),
    .B(_13390_),
    .COUT(_13391_),
    .SUM(_13392_));
 sky130_fd_sc_hd__ha_4 _27654_ (.A(_12288_),
    .B(_12298_),
    .COUT(_13394_),
    .SUM(_13395_));
 sky130_fd_sc_hd__ha_1 _27655_ (.A(_13396_),
    .B(_13397_),
    .COUT(_13398_),
    .SUM(_13399_));
 sky130_fd_sc_hd__ha_4 _27656_ (.A(_12297_),
    .B(_12307_),
    .COUT(_13401_),
    .SUM(_13402_));
 sky130_fd_sc_hd__ha_1 _27657_ (.A(_13403_),
    .B(_13404_),
    .COUT(_13405_),
    .SUM(_13406_));
 sky130_fd_sc_hd__ha_1 _27658_ (.A(_12306_),
    .B(_12316_),
    .COUT(_13408_),
    .SUM(_13409_));
 sky130_fd_sc_hd__ha_4 _27659_ (.A(_13410_),
    .B(_13411_),
    .COUT(_13412_),
    .SUM(_13413_));
 sky130_fd_sc_hd__ha_4 _27660_ (.A(_12315_),
    .B(_12325_),
    .COUT(_13415_),
    .SUM(_13416_));
 sky130_fd_sc_hd__ha_1 _27661_ (.A(_13417_),
    .B(_13418_),
    .COUT(_13419_),
    .SUM(_13420_));
 sky130_fd_sc_hd__ha_4 _27662_ (.A(_12324_),
    .B(_12334_),
    .COUT(_13422_),
    .SUM(_13423_));
 sky130_fd_sc_hd__ha_1 _27663_ (.A(_13424_),
    .B(_13425_),
    .COUT(_13426_),
    .SUM(_13427_));
 sky130_fd_sc_hd__ha_1 _27664_ (.A(_12333_),
    .B(_12343_),
    .COUT(_13429_),
    .SUM(_13430_));
 sky130_fd_sc_hd__ha_1 _27665_ (.A(_13431_),
    .B(_13432_),
    .COUT(_13433_),
    .SUM(_13434_));
 sky130_fd_sc_hd__ha_4 _27666_ (.A(_12342_),
    .B(_12352_),
    .COUT(_13436_),
    .SUM(_13437_));
 sky130_fd_sc_hd__ha_1 _27667_ (.A(_13438_),
    .B(_13439_),
    .COUT(_13440_),
    .SUM(_13441_));
 sky130_fd_sc_hd__ha_4 _27668_ (.A(_12351_),
    .B(_12361_),
    .COUT(_13443_),
    .SUM(_13444_));
 sky130_fd_sc_hd__ha_4 _27669_ (.A(\hash.CA2.p5[0] ),
    .B(_13232_),
    .COUT(_12362_),
    .SUM(_13445_));
 sky130_fd_sc_hd__ha_1 _27670_ (.A(\hash.CA2.p5[1] ),
    .B(_12363_),
    .COUT(_13446_),
    .SUM(_13447_));
 sky130_fd_sc_hd__ha_4 _27671_ (.A(\hash.CA2.p5[2] ),
    .B(_13246_),
    .COUT(_13448_),
    .SUM(_13449_));
 sky130_fd_sc_hd__ha_4 _27672_ (.A(\hash.CA2.p5[3] ),
    .B(_13253_),
    .COUT(_13450_),
    .SUM(_13451_));
 sky130_fd_sc_hd__ha_4 _27673_ (.A(\hash.CA2.p5[4] ),
    .B(_13260_),
    .COUT(_13452_),
    .SUM(_13453_));
 sky130_fd_sc_hd__ha_4 _27674_ (.A(\hash.CA2.p5[5] ),
    .B(_13267_),
    .COUT(_13454_),
    .SUM(_13455_));
 sky130_fd_sc_hd__ha_4 _27675_ (.A(\hash.CA2.p5[6] ),
    .B(_13274_),
    .COUT(_13456_),
    .SUM(_13457_));
 sky130_fd_sc_hd__ha_1 _27676_ (.A(\hash.CA2.p5[7] ),
    .B(_13281_),
    .COUT(_13458_),
    .SUM(_13459_));
 sky130_fd_sc_hd__ha_4 _27677_ (.A(_13288_),
    .B(\hash.CA2.p5[8] ),
    .COUT(_13460_),
    .SUM(_13461_));
 sky130_fd_sc_hd__ha_4 _27678_ (.A(\hash.CA2.p5[9] ),
    .B(_13295_),
    .COUT(_13462_),
    .SUM(_13463_));
 sky130_fd_sc_hd__ha_2 _27679_ (.A(\hash.CA2.p5[10] ),
    .B(_13302_),
    .COUT(_13464_),
    .SUM(_13465_));
 sky130_fd_sc_hd__ha_1 _27680_ (.A(\hash.CA2.p5[11] ),
    .B(_13309_),
    .COUT(_13466_),
    .SUM(_13467_));
 sky130_fd_sc_hd__ha_4 _27681_ (.A(_13316_),
    .B(\hash.CA2.p5[12] ),
    .COUT(_13468_),
    .SUM(_13469_));
 sky130_fd_sc_hd__ha_1 _27682_ (.A(\hash.CA2.p5[13] ),
    .B(_13323_),
    .COUT(_13470_),
    .SUM(_13471_));
 sky130_fd_sc_hd__ha_4 _27683_ (.A(\hash.CA2.p5[14] ),
    .B(_13330_),
    .COUT(_13472_),
    .SUM(_13473_));
 sky130_fd_sc_hd__ha_4 _27684_ (.A(\hash.CA2.p5[15] ),
    .B(_13337_),
    .COUT(_13474_),
    .SUM(_13475_));
 sky130_fd_sc_hd__ha_4 _27685_ (.A(\hash.CA2.p5[16] ),
    .B(_13344_),
    .COUT(_13476_),
    .SUM(_13477_));
 sky130_fd_sc_hd__ha_4 _27686_ (.A(\hash.CA2.p5[17] ),
    .B(_13351_),
    .COUT(_13478_),
    .SUM(_13479_));
 sky130_fd_sc_hd__ha_1 _27687_ (.A(\hash.CA2.p5[16] ),
    .B(_13344_),
    .COUT(_13480_),
    .SUM(_13481_));
 sky130_fd_sc_hd__ha_1 _27688_ (.A(\hash.CA2.p5[18] ),
    .B(_13358_),
    .COUT(_13482_),
    .SUM(_13483_));
 sky130_fd_sc_hd__ha_1 _27689_ (.A(\hash.CA2.p5[19] ),
    .B(_13365_),
    .COUT(_13484_),
    .SUM(_13485_));
 sky130_fd_sc_hd__ha_1 _27690_ (.A(\hash.CA2.p5[20] ),
    .B(_13372_),
    .COUT(_13486_),
    .SUM(_13487_));
 sky130_fd_sc_hd__ha_1 _27691_ (.A(\hash.CA2.p5[21] ),
    .B(_13379_),
    .COUT(_13488_),
    .SUM(_13489_));
 sky130_fd_sc_hd__ha_1 _27692_ (.A(\hash.CA2.p5[20] ),
    .B(_13372_),
    .COUT(_13490_),
    .SUM(_13491_));
 sky130_fd_sc_hd__ha_1 _27693_ (.A(\hash.CA2.p5[22] ),
    .B(_13386_),
    .COUT(_13492_),
    .SUM(_13493_));
 sky130_fd_sc_hd__ha_4 _27694_ (.A(\hash.CA2.p5[21] ),
    .B(net1079),
    .COUT(_13494_),
    .SUM(_13495_));
 sky130_fd_sc_hd__ha_2 _27695_ (.A(\hash.CA2.p5[23] ),
    .B(_13393_),
    .COUT(_13496_),
    .SUM(_13497_));
 sky130_fd_sc_hd__ha_2 _27696_ (.A(\hash.CA2.p5[22] ),
    .B(_13386_),
    .COUT(_13498_),
    .SUM(_13499_));
 sky130_fd_sc_hd__ha_1 _27697_ (.A(\hash.CA2.p5[24] ),
    .B(_13400_),
    .COUT(_13500_),
    .SUM(_13501_));
 sky130_fd_sc_hd__ha_2 _27698_ (.A(\hash.CA2.p5[23] ),
    .B(_13393_),
    .COUT(_13502_),
    .SUM(_13503_));
 sky130_fd_sc_hd__ha_1 _27699_ (.A(\hash.CA2.p5[25] ),
    .B(_13407_),
    .COUT(_13504_),
    .SUM(_13505_));
 sky130_fd_sc_hd__ha_4 _27700_ (.A(_13414_),
    .B(\hash.CA2.p5[26] ),
    .COUT(_13506_),
    .SUM(_13507_));
 sky130_fd_sc_hd__ha_1 _27701_ (.A(\hash.CA2.p5[25] ),
    .B(_13407_),
    .COUT(_13508_),
    .SUM(_13509_));
 sky130_fd_sc_hd__ha_4 _27702_ (.A(\hash.CA2.p5[27] ),
    .B(_13421_),
    .COUT(_13510_),
    .SUM(_13511_));
 sky130_fd_sc_hd__ha_1 _27703_ (.A(\hash.CA2.p5[26] ),
    .B(_13414_),
    .COUT(_13512_),
    .SUM(_13513_));
 sky130_fd_sc_hd__ha_4 _27704_ (.A(\hash.CA2.p5[28] ),
    .B(_13428_),
    .COUT(_13514_),
    .SUM(_13515_));
 sky130_fd_sc_hd__ha_4 _27705_ (.A(\hash.CA2.p5[29] ),
    .B(_13435_),
    .COUT(_13516_),
    .SUM(_13517_));
 sky130_fd_sc_hd__ha_1 _27706_ (.A(\hash.CA2.p5[30] ),
    .B(_13442_),
    .COUT(_13518_),
    .SUM(_13519_));
 sky130_fd_sc_hd__ha_1 _27707_ (.A(net417),
    .B(net412),
    .COUT(_13520_),
    .SUM(_00643_));
 sky130_fd_sc_hd__ha_1 _27708_ (.A(net537),
    .B(\count15_1[2] ),
    .COUT(_13521_),
    .SUM(_00644_));
 sky130_fd_sc_hd__ha_1 _27709_ (.A(net556),
    .B(\count16_1[2] ),
    .COUT(_13522_),
    .SUM(_00645_));
 sky130_fd_sc_hd__ha_1 _27710_ (.A(net435),
    .B(\count2_2[2] ),
    .COUT(_13523_),
    .SUM(_00646_));
 sky130_fd_sc_hd__ha_1 _27711_ (.A(net544),
    .B(\count7_2[2] ),
    .COUT(_13524_),
    .SUM(_00647_));
 sky130_fd_sc_hd__ha_1 _27712_ (.A(net517),
    .B(net557),
    .COUT(_13525_),
    .SUM(_00648_));
 sky130_fd_sc_hd__ha_1 _27713_ (.A(net477),
    .B(\count16_2[2] ),
    .COUT(_13526_),
    .SUM(_00649_));
 sky130_fd_sc_hd__ha_4 _27714_ (.A(_00650_),
    .B(_13527_),
    .COUT(_13528_),
    .SUM(_00651_));
 sky130_fd_sc_hd__ha_4 _27715_ (.A(_00650_),
    .B(\count_1[2] ),
    .COUT(_13529_),
    .SUM(_13530_));
 sky130_fd_sc_hd__ha_4 _27716_ (.A(\count_1[1] ),
    .B(_13527_),
    .COUT(_13531_),
    .SUM(_13532_));
 sky130_fd_sc_hd__ha_4 _27717_ (.A(\count_1[1] ),
    .B(\count_1[2] ),
    .COUT(_13533_),
    .SUM(_13534_));
 sky130_fd_sc_hd__ha_4 _27718_ (.A(_00652_),
    .B(_13535_),
    .COUT(_13536_),
    .SUM(_00653_));
 sky130_fd_sc_hd__ha_4 _27719_ (.A(_00652_),
    .B(\count_2[2] ),
    .COUT(_13537_),
    .SUM(_13538_));
 sky130_fd_sc_hd__ha_4 _27720_ (.A(\count_2[1] ),
    .B(_13535_),
    .COUT(_13539_),
    .SUM(_13540_));
 sky130_fd_sc_hd__ha_4 _27721_ (.A(\count_2[1] ),
    .B(\count_2[2] ),
    .COUT(_13541_),
    .SUM(_13542_));
 sky130_fd_sc_hd__ha_1 _27722_ (.A(_00658_),
    .B(_13543_),
    .COUT(_13544_),
    .SUM(_13545_));
 sky130_fd_sc_hd__ha_1 _27723_ (.A(net456),
    .B(net551),
    .COUT(_13546_),
    .SUM(_00642_));
 sky130_fd_sc_hd__ha_1 _27724_ (.A(_13547_),
    .B(_13548_),
    .COUT(_13549_),
    .SUM(_13550_));
 sky130_fd_sc_hd__ha_1 _27725_ (.A(_13551_),
    .B(_13552_),
    .COUT(_13553_),
    .SUM(_13554_));
 sky130_fd_sc_hd__ha_4 _27726_ (.A(_13555_),
    .B(_13556_),
    .COUT(_13557_),
    .SUM(_13558_));
 sky130_fd_sc_hd__ha_1 _27727_ (.A(_13559_),
    .B(_13560_),
    .COUT(_13561_),
    .SUM(_13562_));
 sky130_fd_sc_hd__ha_1 _27728_ (.A(_13563_),
    .B(_13564_),
    .COUT(_13565_),
    .SUM(_13566_));
 sky130_fd_sc_hd__ha_1 _27729_ (.A(_13567_),
    .B(_13568_),
    .COUT(_13569_),
    .SUM(_13570_));
 sky130_fd_sc_hd__ha_1 _27730_ (.A(_13571_),
    .B(_13572_),
    .COUT(_13573_),
    .SUM(_13574_));
 sky130_fd_sc_hd__ha_4 _27731_ (.A(_13575_),
    .B(_13576_),
    .COUT(_13577_),
    .SUM(_13578_));
 sky130_fd_sc_hd__ha_2 _27732_ (.A(_13579_),
    .B(_13580_),
    .COUT(_13581_),
    .SUM(_13582_));
 sky130_fd_sc_hd__ha_4 _27733_ (.A(_13583_),
    .B(_13584_),
    .COUT(_13585_),
    .SUM(_13586_));
 sky130_fd_sc_hd__ha_1 _27734_ (.A(_13587_),
    .B(_13588_),
    .COUT(_13589_),
    .SUM(_13590_));
 sky130_fd_sc_hd__ha_1 _27735_ (.A(_13591_),
    .B(_13592_),
    .COUT(_13593_),
    .SUM(_13594_));
 sky130_fd_sc_hd__ha_4 _27736_ (.A(_13595_),
    .B(_13596_),
    .COUT(_13597_),
    .SUM(_13598_));
 sky130_fd_sc_hd__ha_2 _27737_ (.A(_13599_),
    .B(_13600_),
    .COUT(_13601_),
    .SUM(_13602_));
 sky130_fd_sc_hd__ha_2 _27738_ (.A(_13603_),
    .B(_13604_),
    .COUT(_13605_),
    .SUM(_13606_));
 sky130_fd_sc_hd__ha_2 _27739_ (.A(_13607_),
    .B(_13608_),
    .COUT(_13609_),
    .SUM(_13610_));
 sky130_fd_sc_hd__ha_1 _27740_ (.A(_13611_),
    .B(_13612_),
    .COUT(_13613_),
    .SUM(_13614_));
 sky130_fd_sc_hd__ha_4 _27741_ (.A(_13615_),
    .B(_13616_),
    .COUT(_13617_),
    .SUM(_13618_));
 sky130_fd_sc_hd__ha_4 _27742_ (.A(_13619_),
    .B(_13620_),
    .COUT(_13621_),
    .SUM(_13622_));
 sky130_fd_sc_hd__ha_4 _27743_ (.A(_13623_),
    .B(_13624_),
    .COUT(_13625_),
    .SUM(_13626_));
 sky130_fd_sc_hd__ha_4 _27744_ (.A(_13627_),
    .B(_13628_),
    .COUT(_13629_),
    .SUM(_13630_));
 sky130_fd_sc_hd__ha_1 _27745_ (.A(_13631_),
    .B(_13632_),
    .COUT(_13633_),
    .SUM(_13634_));
 sky130_fd_sc_hd__ha_1 _27746_ (.A(_13635_),
    .B(_13636_),
    .COUT(_13637_),
    .SUM(_13638_));
 sky130_fd_sc_hd__ha_2 _27747_ (.A(_13639_),
    .B(_13640_),
    .COUT(_13641_),
    .SUM(_13642_));
 sky130_fd_sc_hd__ha_1 _27748_ (.A(_13643_),
    .B(_13644_),
    .COUT(_13645_),
    .SUM(_13646_));
 sky130_fd_sc_hd__ha_1 _27749_ (.A(_13647_),
    .B(_13648_),
    .COUT(_13649_),
    .SUM(_13650_));
 sky130_fd_sc_hd__ha_1 _27750_ (.A(_13651_),
    .B(_13652_),
    .COUT(_13653_),
    .SUM(_13654_));
 sky130_fd_sc_hd__ha_1 _27751_ (.A(_13655_),
    .B(_13656_),
    .COUT(_13657_),
    .SUM(_13658_));
 sky130_fd_sc_hd__ha_1 _27752_ (.A(_13659_),
    .B(_13660_),
    .COUT(_13661_),
    .SUM(_13662_));
 sky130_fd_sc_hd__ha_1 _27753_ (.A(_13663_),
    .B(_13664_),
    .COUT(_13665_),
    .SUM(_13666_));
 sky130_fd_sc_hd__ha_1 _27754_ (.A(_13667_),
    .B(_13668_),
    .COUT(_12378_),
    .SUM(\hash.CA1.p4[1] ));
 sky130_fd_sc_hd__ha_1 _27755_ (.A(_12899_),
    .B(\hash.CA1.p4[1] ),
    .COUT(_13669_),
    .SUM(_13670_));
 sky130_fd_sc_hd__ha_1 _27756_ (.A(_12379_),
    .B(_12377_),
    .COUT(_13671_),
    .SUM(_13672_));
 sky130_fd_sc_hd__ha_1 _27757_ (.A(\hash.CA1.p4[2] ),
    .B(_13673_),
    .COUT(_13674_),
    .SUM(_13675_));
 sky130_fd_sc_hd__ha_1 _27758_ (.A(_12376_),
    .B(_13676_),
    .COUT(_13677_),
    .SUM(_13678_));
 sky130_fd_sc_hd__ha_1 _27759_ (.A(\hash.CA1.p4[3] ),
    .B(_13679_),
    .COUT(_13680_),
    .SUM(_13681_));
 sky130_fd_sc_hd__ha_1 _27760_ (.A(_13682_),
    .B(_12388_),
    .COUT(_13683_),
    .SUM(_13684_));
 sky130_fd_sc_hd__ha_4 _27761_ (.A(\hash.CA1.p4[4] ),
    .B(_13685_),
    .COUT(_13686_),
    .SUM(_13687_));
 sky130_fd_sc_hd__ha_1 _27762_ (.A(_12387_),
    .B(_13688_),
    .COUT(_13689_),
    .SUM(_13690_));
 sky130_fd_sc_hd__ha_4 _27763_ (.A(\hash.CA1.p4[5] ),
    .B(_13691_),
    .COUT(_13692_),
    .SUM(_13693_));
 sky130_fd_sc_hd__ha_2 _27764_ (.A(_13694_),
    .B(_12396_),
    .COUT(_13695_),
    .SUM(_13696_));
 sky130_fd_sc_hd__ha_4 _27765_ (.A(\hash.CA1.p4[6] ),
    .B(_13697_),
    .COUT(_13698_),
    .SUM(_13699_));
 sky130_fd_sc_hd__ha_1 _27766_ (.A(_12395_),
    .B(_13700_),
    .COUT(_13701_),
    .SUM(_13702_));
 sky130_fd_sc_hd__ha_2 _27767_ (.A(\hash.CA1.p4[7] ),
    .B(_13703_),
    .COUT(_13704_),
    .SUM(_13705_));
 sky130_fd_sc_hd__ha_1 _27768_ (.A(_13706_),
    .B(_13707_),
    .COUT(_13708_),
    .SUM(_13709_));
 sky130_fd_sc_hd__ha_1 _27769_ (.A(\hash.CA1.p4[8] ),
    .B(_13710_),
    .COUT(_13711_),
    .SUM(_13712_));
 sky130_fd_sc_hd__ha_4 _27770_ (.A(_13713_),
    .B(_12409_),
    .COUT(_13714_),
    .SUM(_13715_));
 sky130_fd_sc_hd__ha_1 _27771_ (.A(\hash.CA1.p4[9] ),
    .B(_13716_),
    .COUT(_13717_),
    .SUM(_13718_));
 sky130_fd_sc_hd__ha_4 _27772_ (.A(_12408_),
    .B(_12412_),
    .COUT(_13719_),
    .SUM(_13720_));
 sky130_fd_sc_hd__ha_1 _27773_ (.A(\hash.CA1.p4[10] ),
    .B(_13721_),
    .COUT(_13722_),
    .SUM(_13723_));
 sky130_fd_sc_hd__ha_4 _27774_ (.A(_12411_),
    .B(_13724_),
    .COUT(_13725_),
    .SUM(_13726_));
 sky130_fd_sc_hd__ha_2 _27775_ (.A(\hash.CA1.p4[11] ),
    .B(_13727_),
    .COUT(_13728_),
    .SUM(_13729_));
 sky130_fd_sc_hd__ha_4 _27776_ (.A(_13730_),
    .B(_13731_),
    .COUT(_13732_),
    .SUM(_13733_));
 sky130_fd_sc_hd__ha_2 _27777_ (.A(\hash.CA1.p4[12] ),
    .B(_13734_),
    .COUT(_13735_),
    .SUM(_13736_));
 sky130_fd_sc_hd__ha_1 _27778_ (.A(_13737_),
    .B(_12425_),
    .COUT(_13738_),
    .SUM(_13739_));
 sky130_fd_sc_hd__ha_4 _27779_ (.A(\hash.CA1.p4[13] ),
    .B(_13740_),
    .COUT(_13741_),
    .SUM(_13742_));
 sky130_fd_sc_hd__ha_1 _27780_ (.A(_12424_),
    .B(_13743_),
    .COUT(_13744_),
    .SUM(_13745_));
 sky130_fd_sc_hd__ha_2 _27781_ (.A(\hash.CA1.p4[14] ),
    .B(_13746_),
    .COUT(_13747_),
    .SUM(_13748_));
 sky130_fd_sc_hd__ha_2 _27782_ (.A(_13749_),
    .B(_13750_),
    .COUT(_13751_),
    .SUM(_13752_));
 sky130_fd_sc_hd__ha_1 _27783_ (.A(\hash.CA1.p4[15] ),
    .B(_13753_),
    .COUT(_13754_),
    .SUM(_13755_));
 sky130_fd_sc_hd__ha_1 _27784_ (.A(_13756_),
    .B(_13757_),
    .COUT(_13758_),
    .SUM(_13759_));
 sky130_fd_sc_hd__ha_1 _27785_ (.A(\hash.CA1.p4[16] ),
    .B(_13760_),
    .COUT(_13761_),
    .SUM(_13762_));
 sky130_fd_sc_hd__ha_2 _27786_ (.A(_13763_),
    .B(_13764_),
    .COUT(_13765_),
    .SUM(_13766_));
 sky130_fd_sc_hd__ha_1 _27787_ (.A(\hash.CA1.p4[17] ),
    .B(_13767_),
    .COUT(_13768_),
    .SUM(_13769_));
 sky130_fd_sc_hd__ha_2 _27788_ (.A(_13770_),
    .B(_12448_),
    .COUT(_13771_),
    .SUM(_13772_));
 sky130_fd_sc_hd__ha_1 _27789_ (.A(\hash.CA1.p4[18] ),
    .B(_13773_),
    .COUT(_13774_),
    .SUM(_13775_));
 sky130_fd_sc_hd__ha_4 _27790_ (.A(_12447_),
    .B(_12451_),
    .COUT(_13776_),
    .SUM(_13777_));
 sky130_fd_sc_hd__ha_1 _27791_ (.A(\hash.CA1.p4[19] ),
    .B(_13778_),
    .COUT(_13779_),
    .SUM(_13780_));
 sky130_fd_sc_hd__ha_4 _27792_ (.A(_12450_),
    .B(_12454_),
    .COUT(_13781_),
    .SUM(_13782_));
 sky130_fd_sc_hd__ha_1 _27793_ (.A(\hash.CA1.p4[20] ),
    .B(_13783_),
    .COUT(_13784_),
    .SUM(_13785_));
 sky130_fd_sc_hd__ha_4 _27794_ (.A(_12453_),
    .B(_12457_),
    .COUT(_13786_),
    .SUM(_13787_));
 sky130_fd_sc_hd__ha_1 _27795_ (.A(\hash.CA1.p4[21] ),
    .B(_13788_),
    .COUT(_13789_),
    .SUM(_13790_));
 sky130_fd_sc_hd__ha_1 _27796_ (.A(_12456_),
    .B(_12460_),
    .COUT(_13791_),
    .SUM(_13792_));
 sky130_fd_sc_hd__ha_1 _27797_ (.A(\hash.CA1.p4[22] ),
    .B(_13793_),
    .COUT(_13794_),
    .SUM(_13795_));
 sky130_fd_sc_hd__ha_1 _27798_ (.A(_12459_),
    .B(_13796_),
    .COUT(_13797_),
    .SUM(_13798_));
 sky130_fd_sc_hd__ha_1 _27799_ (.A(\hash.CA1.p4[23] ),
    .B(_13799_),
    .COUT(_13800_),
    .SUM(_13801_));
 sky130_fd_sc_hd__ha_1 _27800_ (.A(_13802_),
    .B(_13803_),
    .COUT(_13804_),
    .SUM(_13805_));
 sky130_fd_sc_hd__ha_1 _27801_ (.A(\hash.CA1.p4[24] ),
    .B(_13806_),
    .COUT(_13807_),
    .SUM(_13808_));
 sky130_fd_sc_hd__ha_1 _27802_ (.A(_13809_),
    .B(_13810_),
    .COUT(_13811_),
    .SUM(_13812_));
 sky130_fd_sc_hd__ha_1 _27803_ (.A(\hash.CA1.p4[25] ),
    .B(_13813_),
    .COUT(_13814_),
    .SUM(_13815_));
 sky130_fd_sc_hd__ha_1 _27804_ (.A(_13816_),
    .B(_13817_),
    .COUT(_13818_),
    .SUM(_13819_));
 sky130_fd_sc_hd__ha_2 _27805_ (.A(\hash.CA1.p4[26] ),
    .B(_06287_),
    .COUT(_13821_),
    .SUM(_13822_));
 sky130_fd_sc_hd__ha_4 _27806_ (.A(_13823_),
    .B(_13824_),
    .COUT(_13825_),
    .SUM(_13826_));
 sky130_fd_sc_hd__ha_2 _27807_ (.A(\hash.CA1.p4[27] ),
    .B(_13827_),
    .COUT(_13828_),
    .SUM(_13829_));
 sky130_fd_sc_hd__ha_4 _27808_ (.A(_13830_),
    .B(_13831_),
    .COUT(_13832_),
    .SUM(_13833_));
 sky130_fd_sc_hd__ha_1 _27809_ (.A(\hash.CA1.p4[28] ),
    .B(_13834_),
    .COUT(_13835_),
    .SUM(_13836_));
 sky130_fd_sc_hd__ha_2 _27810_ (.A(_13837_),
    .B(_12493_),
    .COUT(_13838_),
    .SUM(_13839_));
 sky130_fd_sc_hd__ha_1 _27811_ (.A(\hash.CA1.p4[29] ),
    .B(_13840_),
    .COUT(_13841_),
    .SUM(_13842_));
 sky130_fd_sc_hd__ha_1 _27812_ (.A(_12492_),
    .B(_12496_),
    .COUT(_13843_),
    .SUM(_13844_));
 sky130_fd_sc_hd__ha_1 _27813_ (.A(\hash.CA1.p4[30] ),
    .B(_13845_),
    .COUT(_13846_),
    .SUM(_13847_));
 sky130_fd_sc_hd__ha_4 _27814_ (.A(_12653_),
    .B(_12505_),
    .COUT(_13848_),
    .SUM(_11578_));
 sky130_fd_sc_hd__ha_1 _27815_ (.A(_00843_),
    .B(_12368_),
    .COUT(_13849_),
    .SUM(_13850_));
 sky130_fd_sc_hd__ha_4 _27816_ (.A(_00813_),
    .B(_13851_),
    .COUT(_13852_),
    .SUM(_13853_));
 sky130_fd_sc_hd__ha_4 _27817_ (.A(_13854_),
    .B(_00781_),
    .COUT(_13855_),
    .SUM(_13856_));
 sky130_fd_sc_hd__ha_4 _27818_ (.A(_12657_),
    .B(_13857_),
    .COUT(_13858_),
    .SUM(_11577_));
 sky130_fd_sc_hd__ha_4 _27819_ (.A(_12899_),
    .B(_13673_),
    .COUT(_13859_),
    .SUM(_11576_));
 sky130_fd_sc_hd__ha_4 _27820_ (.A(\hash.CA1.b[1] ),
    .B(\hash.CA1.b[0] ),
    .COUT(_13860_),
    .SUM(_11575_));
 sky130_fd_sc_hd__ha_4 _27821_ (.A(\hash.CA1.k_i1[0] ),
    .B(\hash.CA1.w_i1[0] ),
    .COUT(_12497_),
    .SUM(_12654_));
 sky130_fd_sc_hd__ha_2 _27822_ (.A(_13861_),
    .B(_13862_),
    .COUT(_12500_),
    .SUM(_12887_));
 sky130_fd_sc_hd__ha_1 _27823_ (.A(\hash.CA1.k_i1[1] ),
    .B(\hash.CA1.w_i1[1] ),
    .COUT(_13863_),
    .SUM(_13864_));
 sky130_fd_sc_hd__ha_1 _27824_ (.A(_12501_),
    .B(_12502_),
    .COUT(_13865_),
    .SUM(_13866_));
 sky130_fd_sc_hd__ha_1 _27825_ (.A(\hash.CA1.k_i1[2] ),
    .B(\hash.CA1.w_i1[2] ),
    .COUT(_13867_),
    .SUM(_13868_));
 sky130_fd_sc_hd__ha_1 _27826_ (.A(_13869_),
    .B(_13870_),
    .COUT(_13871_),
    .SUM(_13872_));
 sky130_fd_sc_hd__ha_1 _27827_ (.A(_12506_),
    .B(_12512_),
    .COUT(_13873_),
    .SUM(_13874_));
 sky130_fd_sc_hd__ha_1 _27828_ (.A(\hash.CA1.k_i1[3] ),
    .B(\hash.CA1.w_i1[3] ),
    .COUT(_13875_),
    .SUM(_13876_));
 sky130_fd_sc_hd__ha_2 _27829_ (.A(_13877_),
    .B(_13878_),
    .COUT(_13879_),
    .SUM(_13880_));
 sky130_fd_sc_hd__ha_4 _27830_ (.A(_12511_),
    .B(_13881_),
    .COUT(_13882_),
    .SUM(_13883_));
 sky130_fd_sc_hd__ha_1 _27831_ (.A(\hash.CA1.k_i1[4] ),
    .B(\hash.CA1.w_i1[4] ),
    .COUT(_13884_),
    .SUM(_13885_));
 sky130_fd_sc_hd__ha_1 _27832_ (.A(_13887_),
    .B(_13886_),
    .COUT(_13888_),
    .SUM(_13889_));
 sky130_fd_sc_hd__ha_1 _27833_ (.A(_13890_),
    .B(_13891_),
    .COUT(_13892_),
    .SUM(_13893_));
 sky130_fd_sc_hd__ha_4 _27834_ (.A(\hash.CA1.k_i1[5] ),
    .B(\hash.CA1.w_i1[5] ),
    .COUT(_13894_),
    .SUM(_13895_));
 sky130_fd_sc_hd__ha_2 _27835_ (.A(_13897_),
    .B(_13896_),
    .COUT(_13898_),
    .SUM(_13899_));
 sky130_fd_sc_hd__ha_1 _27836_ (.A(_13900_),
    .B(_12527_),
    .COUT(_13901_),
    .SUM(_13902_));
 sky130_fd_sc_hd__ha_1 _27837_ (.A(\hash.CA1.k_i1[6] ),
    .B(\hash.CA1.w_i1[6] ),
    .COUT(_13903_),
    .SUM(_13904_));
 sky130_fd_sc_hd__ha_2 _27838_ (.A(_13905_),
    .B(_13906_),
    .COUT(_13907_),
    .SUM(_13908_));
 sky130_fd_sc_hd__ha_1 _27839_ (.A(_12526_),
    .B(_12532_),
    .COUT(_13909_),
    .SUM(_13910_));
 sky130_fd_sc_hd__ha_1 _27840_ (.A(\hash.CA1.k_i1[7] ),
    .B(\hash.CA1.w_i1[7] ),
    .COUT(_13911_),
    .SUM(_13912_));
 sky130_fd_sc_hd__ha_4 _27841_ (.A(_13913_),
    .B(_13914_),
    .COUT(_13915_),
    .SUM(_13916_));
 sky130_fd_sc_hd__ha_4 _27842_ (.A(_12531_),
    .B(_12537_),
    .COUT(_13917_),
    .SUM(_13918_));
 sky130_fd_sc_hd__ha_1 _27843_ (.A(\hash.CA1.k_i1[8] ),
    .B(\hash.CA1.w_i1[8] ),
    .COUT(_13919_),
    .SUM(_13920_));
 sky130_fd_sc_hd__ha_4 _27844_ (.A(_13921_),
    .B(_13922_),
    .COUT(_13923_),
    .SUM(_13924_));
 sky130_fd_sc_hd__ha_4 _27845_ (.A(_12536_),
    .B(_13925_),
    .COUT(_13926_),
    .SUM(_13927_));
 sky130_fd_sc_hd__ha_1 _27846_ (.A(\hash.CA1.k_i1[9] ),
    .B(\hash.CA1.w_i1[9] ),
    .COUT(_13928_),
    .SUM(_13929_));
 sky130_fd_sc_hd__ha_1 _27847_ (.A(_13930_),
    .B(_13931_),
    .COUT(_13932_),
    .SUM(_13933_));
 sky130_fd_sc_hd__ha_4 _27848_ (.A(_13934_),
    .B(_12547_),
    .COUT(_13935_),
    .SUM(_13936_));
 sky130_fd_sc_hd__ha_1 _27849_ (.A(\hash.CA1.k_i1[10] ),
    .B(\hash.CA1.w_i1[10] ),
    .COUT(_13937_),
    .SUM(_13938_));
 sky130_fd_sc_hd__ha_1 _27850_ (.A(_13939_),
    .B(_13940_),
    .COUT(_13941_),
    .SUM(_13942_));
 sky130_fd_sc_hd__ha_4 _27851_ (.A(_12546_),
    .B(_13943_),
    .COUT(_13944_),
    .SUM(_13945_));
 sky130_fd_sc_hd__ha_1 _27852_ (.A(\hash.CA1.k_i1[11] ),
    .B(\hash.CA1.w_i1[11] ),
    .COUT(_13946_),
    .SUM(_13947_));
 sky130_fd_sc_hd__ha_4 _27853_ (.A(_13948_),
    .B(_13949_),
    .COUT(_13950_),
    .SUM(_13951_));
 sky130_fd_sc_hd__ha_4 _27854_ (.A(_13952_),
    .B(_13953_),
    .COUT(_13954_),
    .SUM(_13955_));
 sky130_fd_sc_hd__ha_1 _27855_ (.A(\hash.CA1.k_i1[12] ),
    .B(\hash.CA1.w_i1[12] ),
    .COUT(_13956_),
    .SUM(_13957_));
 sky130_fd_sc_hd__ha_1 _27856_ (.A(_13958_),
    .B(_13959_),
    .COUT(_13960_),
    .SUM(_13961_));
 sky130_fd_sc_hd__ha_4 _27857_ (.A(_13962_),
    .B(_12562_),
    .COUT(_13963_),
    .SUM(_13964_));
 sky130_fd_sc_hd__ha_1 _27858_ (.A(\hash.CA1.k_i1[13] ),
    .B(\hash.CA1.w_i1[13] ),
    .COUT(_13965_),
    .SUM(_13966_));
 sky130_fd_sc_hd__ha_4 _27859_ (.A(_13967_),
    .B(_13968_),
    .COUT(_13969_),
    .SUM(_13970_));
 sky130_fd_sc_hd__ha_1 _27860_ (.A(_12561_),
    .B(_12567_),
    .COUT(_13971_),
    .SUM(_13972_));
 sky130_fd_sc_hd__ha_4 _27861_ (.A(\hash.CA1.k_i1[14] ),
    .B(\hash.CA1.w_i1[14] ),
    .COUT(_13973_),
    .SUM(_13974_));
 sky130_fd_sc_hd__ha_4 _27862_ (.A(_13975_),
    .B(_13976_),
    .COUT(_13977_),
    .SUM(_13978_));
 sky130_fd_sc_hd__ha_4 _27863_ (.A(_12566_),
    .B(_13979_),
    .COUT(_13980_),
    .SUM(_13981_));
 sky130_fd_sc_hd__ha_1 _27864_ (.A(\hash.CA1.k_i1[15] ),
    .B(\hash.CA1.w_i1[15] ),
    .COUT(_13982_),
    .SUM(_13983_));
 sky130_fd_sc_hd__ha_4 _27865_ (.A(_13984_),
    .B(_13985_),
    .COUT(_13986_),
    .SUM(_13987_));
 sky130_fd_sc_hd__ha_4 _27866_ (.A(_13988_),
    .B(_13989_),
    .COUT(_13990_),
    .SUM(_13991_));
 sky130_fd_sc_hd__ha_1 _27867_ (.A(\hash.CA1.k_i1[16] ),
    .B(\hash.CA1.w_i1[16] ),
    .COUT(_13992_),
    .SUM(_13993_));
 sky130_fd_sc_hd__ha_2 _27868_ (.A(_13994_),
    .B(_13995_),
    .COUT(_13996_),
    .SUM(_13997_));
 sky130_fd_sc_hd__ha_4 _27869_ (.A(_13998_),
    .B(_12582_),
    .COUT(_13999_),
    .SUM(_14000_));
 sky130_fd_sc_hd__ha_1 _27870_ (.A(\hash.CA1.k_i1[17] ),
    .B(\hash.CA1.w_i1[17] ),
    .COUT(_14001_),
    .SUM(_14002_));
 sky130_fd_sc_hd__ha_4 _27871_ (.A(_14003_),
    .B(_14004_),
    .COUT(_14005_),
    .SUM(_14006_));
 sky130_fd_sc_hd__ha_4 _27872_ (.A(_12581_),
    .B(_12587_),
    .COUT(_14007_),
    .SUM(_14008_));
 sky130_fd_sc_hd__ha_1 _27873_ (.A(\hash.CA1.k_i1[18] ),
    .B(\hash.CA1.w_i1[18] ),
    .COUT(_14009_),
    .SUM(_14010_));
 sky130_fd_sc_hd__ha_2 _27874_ (.A(_14011_),
    .B(_14012_),
    .COUT(_14013_),
    .SUM(_14014_));
 sky130_fd_sc_hd__ha_4 _27875_ (.A(_12586_),
    .B(_12592_),
    .COUT(_14015_),
    .SUM(_14016_));
 sky130_fd_sc_hd__ha_1 _27876_ (.A(\hash.CA1.k_i1[19] ),
    .B(\hash.CA1.w_i1[19] ),
    .COUT(_14017_),
    .SUM(_14018_));
 sky130_fd_sc_hd__ha_1 _27877_ (.A(_14019_),
    .B(_14020_),
    .COUT(_14021_),
    .SUM(_14022_));
 sky130_fd_sc_hd__ha_4 _27878_ (.A(_12591_),
    .B(_12597_),
    .COUT(_14023_),
    .SUM(_14024_));
 sky130_fd_sc_hd__ha_1 _27879_ (.A(\hash.CA1.k_i1[20] ),
    .B(\hash.CA1.w_i1[20] ),
    .COUT(_14025_),
    .SUM(_14026_));
 sky130_fd_sc_hd__ha_1 _27880_ (.A(_14027_),
    .B(_14028_),
    .COUT(_14029_),
    .SUM(_14030_));
 sky130_fd_sc_hd__ha_2 _27881_ (.A(_12596_),
    .B(_12602_),
    .COUT(_14031_),
    .SUM(_14032_));
 sky130_fd_sc_hd__ha_2 _27882_ (.A(\hash.CA1.k_i1[21] ),
    .B(\hash.CA1.w_i1[21] ),
    .COUT(_14033_),
    .SUM(_14034_));
 sky130_fd_sc_hd__ha_1 _27883_ (.A(_14035_),
    .B(_14036_),
    .COUT(_14037_),
    .SUM(_14038_));
 sky130_fd_sc_hd__ha_1 _27884_ (.A(_12601_),
    .B(_14039_),
    .COUT(_14040_),
    .SUM(_14041_));
 sky130_fd_sc_hd__ha_1 _27885_ (.A(\hash.CA1.k_i1[22] ),
    .B(\hash.CA1.w_i1[22] ),
    .COUT(_14042_),
    .SUM(_14043_));
 sky130_fd_sc_hd__ha_1 _27886_ (.A(_14044_),
    .B(_14045_),
    .COUT(_14046_),
    .SUM(_14047_));
 sky130_fd_sc_hd__ha_1 _27887_ (.A(_14048_),
    .B(_14049_),
    .COUT(_14050_),
    .SUM(_14051_));
 sky130_fd_sc_hd__ha_1 _27888_ (.A(\hash.CA1.k_i1[23] ),
    .B(\hash.CA1.w_i1[23] ),
    .COUT(_14052_),
    .SUM(_14053_));
 sky130_fd_sc_hd__ha_1 _27889_ (.A(_14054_),
    .B(_14055_),
    .COUT(_14056_),
    .SUM(_14057_));
 sky130_fd_sc_hd__ha_1 _27890_ (.A(_14058_),
    .B(_14059_),
    .COUT(_14060_),
    .SUM(_14061_));
 sky130_fd_sc_hd__ha_1 _27891_ (.A(\hash.CA1.k_i1[24] ),
    .B(\hash.CA1.w_i1[24] ),
    .COUT(_14062_),
    .SUM(_14063_));
 sky130_fd_sc_hd__ha_2 _27892_ (.A(_14064_),
    .B(_14065_),
    .COUT(_14066_),
    .SUM(_14067_));
 sky130_fd_sc_hd__ha_2 _27893_ (.A(_14068_),
    .B(_14069_),
    .COUT(_14070_),
    .SUM(_14071_));
 sky130_fd_sc_hd__ha_4 _27894_ (.A(\hash.CA1.k_i1[25] ),
    .B(\hash.CA1.w_i1[25] ),
    .COUT(_14072_),
    .SUM(_14073_));
 sky130_fd_sc_hd__ha_4 _27895_ (.A(_14074_),
    .B(_14075_),
    .COUT(_14076_),
    .SUM(_14077_));
 sky130_fd_sc_hd__ha_1 _27896_ (.A(_14078_),
    .B(_14079_),
    .COUT(_14080_),
    .SUM(_14081_));
 sky130_fd_sc_hd__ha_4 _27897_ (.A(\hash.CA1.k_i1[26] ),
    .B(\hash.CA1.w_i1[26] ),
    .COUT(_14082_),
    .SUM(_14083_));
 sky130_fd_sc_hd__ha_2 _27898_ (.A(_14084_),
    .B(_14085_),
    .COUT(_14086_),
    .SUM(_14087_));
 sky130_fd_sc_hd__ha_1 _27899_ (.A(_14088_),
    .B(_12632_),
    .COUT(_14089_),
    .SUM(_14090_));
 sky130_fd_sc_hd__ha_4 _27900_ (.A(\hash.CA1.k_i1[27] ),
    .B(\hash.CA1.w_i1[27] ),
    .COUT(_14091_),
    .SUM(_14092_));
 sky130_fd_sc_hd__ha_4 _27901_ (.A(_14093_),
    .B(_14094_),
    .COUT(_14095_),
    .SUM(_14096_));
 sky130_fd_sc_hd__ha_2 _27902_ (.A(_12631_),
    .B(_14097_),
    .COUT(_14098_),
    .SUM(_14099_));
 sky130_fd_sc_hd__ha_4 _27903_ (.A(\hash.CA1.k_i1[28] ),
    .B(\hash.CA1.w_i1[28] ),
    .COUT(_14100_),
    .SUM(_14101_));
 sky130_fd_sc_hd__ha_1 _27904_ (.A(_14102_),
    .B(_14103_),
    .COUT(_14104_),
    .SUM(_14105_));
 sky130_fd_sc_hd__ha_1 _27905_ (.A(_14106_),
    .B(_14107_),
    .COUT(_14108_),
    .SUM(_14109_));
 sky130_fd_sc_hd__ha_1 _27906_ (.A(\hash.CA1.k_i1[29] ),
    .B(\hash.CA1.w_i1[29] ),
    .COUT(_14110_),
    .SUM(_14111_));
 sky130_fd_sc_hd__ha_1 _27907_ (.A(_14112_),
    .B(_14113_),
    .COUT(_14114_),
    .SUM(_14115_));
 sky130_fd_sc_hd__ha_1 _27908_ (.A(_14116_),
    .B(_12647_),
    .COUT(_14117_),
    .SUM(_14118_));
 sky130_fd_sc_hd__ha_1 _27909_ (.A(\hash.CA1.k_i1[30] ),
    .B(\hash.CA1.w_i1[30] ),
    .COUT(_14119_),
    .SUM(_14120_));
 sky130_fd_sc_hd__ha_1 _27910_ (.A(_14121_),
    .B(_14122_),
    .COUT(_14123_),
    .SUM(_14124_));
 sky130_fd_sc_hd__ha_1 _27911_ (.A(_12646_),
    .B(_14125_),
    .COUT(_14126_),
    .SUM(_14127_));
 sky130_fd_sc_hd__ha_1 _27912_ (.A(_14128_),
    .B(_14129_),
    .COUT(_14130_),
    .SUM(_14131_));
 sky130_fd_sc_hd__ha_1 _27913_ (.A(_14132_),
    .B(_14133_),
    .COUT(_14134_),
    .SUM(_14135_));
 sky130_fd_sc_hd__ha_4 _27914_ (.A(_14136_),
    .B(_14137_),
    .COUT(_14138_),
    .SUM(_14139_));
 sky130_fd_sc_hd__ha_4 _27915_ (.A(_14140_),
    .B(_14141_),
    .COUT(_14142_),
    .SUM(_14143_));
 sky130_fd_sc_hd__ha_4 _27916_ (.A(_14144_),
    .B(_14145_),
    .COUT(_14146_),
    .SUM(_14147_));
 sky130_fd_sc_hd__ha_4 _27917_ (.A(_14148_),
    .B(_14149_),
    .COUT(_14150_),
    .SUM(_14151_));
 sky130_fd_sc_hd__ha_2 _27918_ (.A(_14152_),
    .B(_14153_),
    .COUT(_14154_),
    .SUM(_14155_));
 sky130_fd_sc_hd__ha_4 _27919_ (.A(_14156_),
    .B(_12722_),
    .COUT(_14157_),
    .SUM(_14158_));
 sky130_fd_sc_hd__ha_4 _27920_ (.A(_12730_),
    .B(_12721_),
    .COUT(_14159_),
    .SUM(_14160_));
 sky130_fd_sc_hd__ha_1 _27921_ (.A(_12729_),
    .B(_12739_),
    .COUT(_14161_),
    .SUM(_14162_));
 sky130_fd_sc_hd__ha_4 _27922_ (.A(_12738_),
    .B(_12745_),
    .COUT(_14163_),
    .SUM(_14164_));
 sky130_fd_sc_hd__ha_1 _27923_ (.A(_12744_),
    .B(_12751_),
    .COUT(_14165_),
    .SUM(_14166_));
 sky130_fd_sc_hd__ha_1 _27924_ (.A(_12750_),
    .B(_12758_),
    .COUT(_14167_),
    .SUM(_14168_));
 sky130_fd_sc_hd__ha_2 _27925_ (.A(_12757_),
    .B(_12766_),
    .COUT(_14169_),
    .SUM(_14170_));
 sky130_fd_sc_hd__ha_1 _27926_ (.A(_12765_),
    .B(_12773_),
    .COUT(_14171_),
    .SUM(_14172_));
 sky130_fd_sc_hd__ha_1 _27927_ (.A(_12772_),
    .B(_12779_),
    .COUT(_14173_),
    .SUM(_14174_));
 sky130_fd_sc_hd__ha_1 _27928_ (.A(_12778_),
    .B(_12785_),
    .COUT(_14175_),
    .SUM(_14176_));
 sky130_fd_sc_hd__ha_4 _27929_ (.A(_12784_),
    .B(_12791_),
    .COUT(_14177_),
    .SUM(_14178_));
 sky130_fd_sc_hd__ha_4 _27930_ (.A(_12790_),
    .B(_12800_),
    .COUT(_14179_),
    .SUM(_14180_));
 sky130_fd_sc_hd__ha_2 _27931_ (.A(_12799_),
    .B(_12809_),
    .COUT(_14181_),
    .SUM(_14182_));
 sky130_fd_sc_hd__ha_1 _27932_ (.A(_12808_),
    .B(_12816_),
    .COUT(_14183_),
    .SUM(_14184_));
 sky130_fd_sc_hd__ha_2 _27933_ (.A(_12815_),
    .B(_12825_),
    .COUT(_14185_),
    .SUM(_14186_));
 sky130_fd_sc_hd__ha_4 _27934_ (.A(_12824_),
    .B(_12832_),
    .COUT(_14187_),
    .SUM(_14188_));
 sky130_fd_sc_hd__ha_4 _27935_ (.A(_12831_),
    .B(_12841_),
    .COUT(_14189_),
    .SUM(_14190_));
 sky130_fd_sc_hd__ha_4 _27936_ (.A(_12840_),
    .B(_12847_),
    .COUT(_14191_),
    .SUM(_14192_));
 sky130_fd_sc_hd__ha_4 _27937_ (.A(_12846_),
    .B(_12855_),
    .COUT(_14193_),
    .SUM(_14194_));
 sky130_fd_sc_hd__ha_1 _27938_ (.A(_12854_),
    .B(_12863_),
    .COUT(_14195_),
    .SUM(_14196_));
 sky130_fd_sc_hd__ha_2 _27939_ (.A(_12862_),
    .B(_12869_),
    .COUT(_14197_),
    .SUM(_14198_));
 sky130_fd_sc_hd__ha_1 _27940_ (.A(_12868_),
    .B(_14199_),
    .COUT(_14200_),
    .SUM(_14201_));
 sky130_fd_sc_hd__ha_2 _27941_ (.A(_14202_),
    .B(_14203_),
    .COUT(_14204_),
    .SUM(\hash.CA1.p1[0] ));
 sky130_fd_sc_hd__ha_1 _27942_ (.A(_12656_),
    .B(_12887_),
    .COUT(_14205_),
    .SUM(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__ha_1 _27943_ (.A(_14205_),
    .B(_14206_),
    .COUT(_14207_),
    .SUM(\hash.CA1.p2[1] ));
 sky130_fd_sc_hd__ha_1 _27944_ (.A(_12888_),
    .B(_12507_),
    .COUT(_14208_),
    .SUM(\hash.CA1.p3[1] ));
 sky130_fd_sc_hd__ha_1 _27945_ (.A(\hash.CA1.c[0] ),
    .B(\hash.CA1.p4[0] ),
    .COUT(_12898_),
    .SUM(\hash.CA1.p5[0] ));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[1]$_SDFF_PP0_  (.D(_00907_),
    .Q(\count15_1[1] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[2]$_SDFF_PP0_  (.D(_00908_),
    .Q(\count15_1[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[3]$_SDFF_PP0_  (.D(_00909_),
    .Q(\count15_1[3] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[4]$_SDFF_PP0_  (.D(_00910_),
    .Q(\count15_1[4] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[5]$_SDFF_PP0_  (.D(_00911_),
    .Q(\count15_1[5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_2[1]$_SDFF_PP1_  (.D(_00912_),
    .Q(\count15_2[1] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_2[2]$_SDFF_PP0_  (.D(_00913_),
    .Q(\count15_2[2] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_2[3]$_SDFF_PP0_  (.D(_00914_),
    .Q(\count15_2[3] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_2[4]$_SDFF_PP0_  (.D(_00915_),
    .Q(\count15_2[4] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 \count15_2[5]$_SDFF_PP0_  (.D(_00916_),
    .Q(\count15_2[5] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[1]$_SDFF_PP0_  (.D(_00917_),
    .Q(\count16_1[1] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[2]$_SDFF_PP0_  (.D(_00918_),
    .Q(\count16_1[2] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_1[3]$_SDFF_PP0_  (.D(_00919_),
    .Q(\count16_1[3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[4]$_SDFF_PP0_  (.D(_00920_),
    .Q(\count16_1[4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[5]$_SDFF_PP0_  (.D(_00921_),
    .Q(\count16_1[5] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_2[1]$_SDFF_PP0_  (.D(_00922_),
    .Q(\count16_2[1] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_2[2]$_SDFF_PP0_  (.D(_00923_),
    .Q(\count16_2[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_2[3]$_SDFF_PP0_  (.D(_00924_),
    .Q(\count16_2[3] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_2[4]$_SDFF_PP0_  (.D(_00925_),
    .Q(\count16_2[4] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_2[5]$_SDFF_PP0_  (.D(_00926_),
    .Q(\count16_2[5] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[1]$_SDFF_PP1_  (.D(_00927_),
    .Q(\count2_1[1] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[2]$_SDFF_PP1_  (.D(_00928_),
    .Q(\count2_1[2] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[3]$_SDFF_PP1_  (.D(_00929_),
    .Q(\count2_1[3] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[4]$_SDFF_PP0_  (.D(_00930_),
    .Q(\count2_1[4] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[5]$_SDFF_PP0_  (.D(_00931_),
    .Q(\count2_1[5] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 \count2_2[1]$_SDFF_PP1_  (.D(_00932_),
    .Q(\count2_2[1] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[2]$_SDFF_PP1_  (.D(_00933_),
    .Q(\count2_2[2] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[3]$_SDFF_PP1_  (.D(_00934_),
    .Q(\count2_2[3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[4]$_SDFF_PP0_  (.D(_00935_),
    .Q(\count2_2[4] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 \count2_2[5]$_SDFF_PP0_  (.D(_00936_),
    .Q(\count2_2[5] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[1]$_SDFF_PP0_  (.D(_00937_),
    .Q(\count7_1[1] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[2]$_SDFF_PP0_  (.D(_00938_),
    .Q(\count7_1[2] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[3]$_SDFF_PP1_  (.D(_00939_),
    .Q(\count7_1[3] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[4]$_SDFF_PP0_  (.D(_00940_),
    .Q(\count7_1[4] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[5]$_SDFF_PP0_  (.D(_00941_),
    .Q(\count7_1[5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[1]$_SDFF_PP1_  (.D(_00942_),
    .Q(\count7_2[1] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[2]$_SDFF_PP0_  (.D(_00943_),
    .Q(\count7_2[2] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[3]$_SDFF_PP1_  (.D(_00944_),
    .Q(\count7_2[3] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[4]$_SDFF_PP0_  (.D(_00945_),
    .Q(\count7_2[4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[5]$_SDFF_PP0_  (.D(_00946_),
    .Q(\count7_2[5] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[1]$_SDFFE_PP0N_  (.D(_00947_),
    .Q(\count_1[1] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[2]$_SDFFE_PP0N_  (.D(_00948_),
    .Q(\count_1[2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[3]$_SDFFE_PP0N_  (.D(_00949_),
    .Q(\count_1[3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[4]$_SDFFE_PP1N_  (.D(_00950_),
    .Q(\count_1[4] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[5]$_SDFFE_PP0N_  (.D(_00951_),
    .Q(\count_1[5] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[1]$_SDFFE_PP0N_  (.D(_00952_),
    .Q(\count_2[1] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[2]$_SDFFE_PP0N_  (.D(_00953_),
    .Q(\count_2[2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[3]$_SDFFE_PP0N_  (.D(_00954_),
    .Q(\count_2[3] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[4]$_SDFFE_PP1N_  (.D(_00955_),
    .Q(\count_2[4] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[5]$_SDFFE_PP0N_  (.D(_00956_),
    .Q(\count_2[5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[6]$_SDFFE_PP0N_  (.D(_00957_),
    .Q(\count_2[6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[1]$_SDFFE_PP0N_  (.D(_00958_),
    .Q(\count_hash1[1] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[2]$_SDFFE_PP0N_  (.D(_00959_),
    .Q(\count_hash1[2] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[3]$_SDFFE_PP0N_  (.D(_00960_),
    .Q(\count_hash1[3] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[4]$_SDFFE_PP0N_  (.D(_00961_),
    .Q(\count_hash1[4] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[5]$_SDFFE_PP0N_  (.D(_00962_),
    .Q(\count_hash1[5] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[6]$_SDFFE_PP0N_  (.D(_00963_),
    .Q(\count_hash1[6] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[1]$_SDFFE_PP0N_  (.D(_00964_),
    .Q(\count_hash2[1] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[2]$_SDFFE_PP0N_  (.D(_00965_),
    .Q(\count_hash2[2] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[3]$_SDFFE_PP0N_  (.D(_00966_),
    .Q(\count_hash2[3] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[4]$_SDFFE_PP0N_  (.D(_00967_),
    .Q(\count_hash2[4] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[5]$_SDFFE_PP0N_  (.D(_00968_),
    .Q(\count_hash2[5] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \done$_DFFE_PN_  (.D(_00128_),
    .DE(_09731_),
    .Q(done),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[0]$_DFF_P_  (.D(\hash.CA1.S0.X[0] ),
    .Q(\hash.CA2.a_dash[0] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[10]$_DFF_P_  (.D(\hash.CA1.S0.X[10] ),
    .Q(\hash.CA2.a_dash[10] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[11]$_DFF_P_  (.D(\hash.CA1.S0.X[11] ),
    .Q(\hash.CA2.a_dash[11] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[12]$_DFF_P_  (.D(\hash.CA1.S0.X[12] ),
    .Q(\hash.CA2.a_dash[12] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[13]$_DFF_P_  (.D(\hash.CA1.S0.X[13] ),
    .Q(\hash.CA2.a_dash[13] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[14]$_DFF_P_  (.D(\hash.CA1.S0.X[14] ),
    .Q(\hash.CA2.a_dash[14] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[15]$_DFF_P_  (.D(\hash.CA1.S0.X[15] ),
    .Q(\hash.CA2.a_dash[15] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[16]$_DFF_P_  (.D(\hash.CA1.S0.X[16] ),
    .Q(\hash.CA2.a_dash[16] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[17]$_DFF_P_  (.D(\hash.CA1.S0.X[17] ),
    .Q(\hash.CA2.a_dash[17] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[18]$_DFF_P_  (.D(\hash.CA1.S0.X[18] ),
    .Q(\hash.CA2.a_dash[18] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[19]$_DFF_P_  (.D(\hash.CA1.S0.X[19] ),
    .Q(\hash.CA2.a_dash[19] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[1]$_DFF_P_  (.D(\hash.CA1.S0.X[1] ),
    .Q(\hash.CA2.a_dash[1] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[20]$_DFF_P_  (.D(_06148_),
    .Q(\hash.CA2.a_dash[20] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[21]$_DFF_P_  (.D(_06156_),
    .Q(\hash.CA2.a_dash[21] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[22]$_DFF_P_  (.D(\hash.CA1.S0.X[22] ),
    .Q(\hash.CA2.a_dash[22] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[23]$_DFF_P_  (.D(\hash.CA1.S0.X[23] ),
    .Q(\hash.CA2.a_dash[23] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[24]$_DFF_P_  (.D(_06179_),
    .Q(\hash.CA2.a_dash[24] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[25]$_DFF_P_  (.D(\hash.CA1.S0.X[25] ),
    .Q(\hash.CA2.a_dash[25] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[26]$_DFF_P_  (.D(_06201_),
    .Q(\hash.CA2.a_dash[26] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[27]$_DFF_P_  (.D(_06211_),
    .Q(\hash.CA2.a_dash[27] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[28]$_DFF_P_  (.D(\hash.CA1.S0.X[28] ),
    .Q(\hash.CA2.a_dash[28] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[29]$_DFF_P_  (.D(\hash.CA1.S0.X[29] ),
    .Q(\hash.CA2.a_dash[29] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[2]$_DFF_P_  (.D(\hash.CA1.S0.X[2] ),
    .Q(\hash.CA2.a_dash[2] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[30]$_DFF_P_  (.D(_06234_),
    .Q(\hash.CA2.a_dash[30] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[31]$_DFF_P_  (.D(\hash.CA1.S0.X[31] ),
    .Q(\hash.CA2.a_dash[31] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[3]$_DFF_P_  (.D(\hash.CA1.S0.X[3] ),
    .Q(\hash.CA2.a_dash[3] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[4]$_DFF_P_  (.D(_06010_),
    .Q(\hash.CA2.a_dash[4] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[5]$_DFF_P_  (.D(\hash.CA1.S0.X[5] ),
    .Q(\hash.CA2.a_dash[5] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[6]$_DFF_P_  (.D(\hash.CA1.S0.X[6] ),
    .Q(\hash.CA2.a_dash[6] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[7]$_DFF_P_  (.D(\hash.CA1.S0.X[7] ),
    .Q(\hash.CA2.a_dash[7] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[8]$_DFF_P_  (.D(_06043_),
    .Q(\hash.CA2.a_dash[8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[9]$_DFF_P_  (.D(\hash.CA1.S0.X[9] ),
    .Q(\hash.CA2.a_dash[9] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[0]$_DFF_P_  (.D(\hash.CA1.b[0] ),
    .Q(\hash.CA2.b_dash[0] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[10]$_DFF_P_  (.D(\hash.CA1.b[10] ),
    .Q(\hash.CA2.b_dash[10] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[11]$_DFF_P_  (.D(\hash.CA1.b[11] ),
    .Q(\hash.CA2.b_dash[11] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[12]$_DFF_P_  (.D(_06283_),
    .Q(\hash.CA2.b_dash[12] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[13]$_DFF_P_  (.D(\hash.CA1.b[13] ),
    .Q(\hash.CA2.b_dash[13] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[14]$_DFF_P_  (.D(\hash.CA1.b[14] ),
    .Q(\hash.CA2.b_dash[14] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[15]$_DFF_P_  (.D(\hash.CA1.b[15] ),
    .Q(\hash.CA2.b_dash[15] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[16]$_DFF_P_  (.D(\hash.CA1.b[16] ),
    .Q(\hash.CA2.b_dash[16] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[17]$_DFF_P_  (.D(\hash.CA1.b[17] ),
    .Q(\hash.CA2.b_dash[17] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[18]$_DFF_P_  (.D(\hash.CA1.b[18] ),
    .Q(\hash.CA2.b_dash[18] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[19]$_DFF_P_  (.D(_06284_),
    .Q(\hash.CA2.b_dash[19] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[1]$_DFF_P_  (.D(\hash.CA1.b[1] ),
    .Q(\hash.CA2.b_dash[1] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[20]$_DFF_P_  (.D(\hash.CA1.b[20] ),
    .Q(\hash.CA2.b_dash[20] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[21]$_DFF_P_  (.D(\hash.CA1.b[21] ),
    .Q(\hash.CA2.b_dash[21] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[22]$_DFF_P_  (.D(\hash.CA1.b[22] ),
    .Q(\hash.CA2.b_dash[22] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[23]$_DFF_P_  (.D(_06285_),
    .Q(\hash.CA2.b_dash[23] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[24]$_DFF_P_  (.D(\hash.CA1.b[24] ),
    .Q(\hash.CA2.b_dash[24] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[25]$_DFF_P_  (.D(\hash.CA1.b[25] ),
    .Q(\hash.CA2.b_dash[25] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[26]$_DFF_P_  (.D(\hash.CA1.b[26] ),
    .Q(\hash.CA2.b_dash[26] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[27]$_DFF_P_  (.D(\hash.CA1.b[27] ),
    .Q(\hash.CA2.b_dash[27] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[28]$_DFF_P_  (.D(\hash.CA1.b[28] ),
    .Q(\hash.CA2.b_dash[28] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[29]$_DFF_P_  (.D(\hash.CA1.b[29] ),
    .Q(\hash.CA2.b_dash[29] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[2]$_DFF_P_  (.D(\hash.CA1.b[2] ),
    .Q(\hash.CA2.b_dash[2] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[30]$_DFF_P_  (.D(\hash.CA1.b[30] ),
    .Q(\hash.CA2.b_dash[30] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[31]$_DFF_P_  (.D(\hash.CA1.b[31] ),
    .Q(\hash.CA2.b_dash[31] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[3]$_DFF_P_  (.D(\hash.CA1.b[3] ),
    .Q(\hash.CA2.b_dash[3] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[4]$_DFF_P_  (.D(\hash.CA1.b[4] ),
    .Q(\hash.CA2.b_dash[4] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[5]$_DFF_P_  (.D(\hash.CA1.b[5] ),
    .Q(\hash.CA2.b_dash[5] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[6]$_DFF_P_  (.D(\hash.CA1.b[6] ),
    .Q(\hash.CA2.b_dash[6] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[7]$_DFF_P_  (.D(\hash.CA1.b[7] ),
    .Q(\hash.CA2.b_dash[7] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[8]$_DFF_P_  (.D(_06279_),
    .Q(\hash.CA2.b_dash[8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[9]$_DFF_P_  (.D(_06280_),
    .Q(\hash.CA2.b_dash[9] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[0]$_DFF_P_  (.D(\hash.CA1.S1.X[0] ),
    .Q(\hash.CA2.e_dash[0] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[10]$_DFF_P_  (.D(\hash.CA1.S1.X[10] ),
    .Q(\hash.CA2.e_dash[10] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[11]$_DFF_P_  (.D(_06575_),
    .Q(\hash.CA2.e_dash[11] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[12]$_DFF_P_  (.D(\hash.CA1.S1.X[12] ),
    .Q(\hash.CA2.e_dash[12] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[13]$_DFF_P_  (.D(\hash.CA1.S1.X[13] ),
    .Q(\hash.CA2.e_dash[13] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[14]$_DFF_P_  (.D(\hash.CA1.S1.X[14] ),
    .Q(\hash.CA2.e_dash[14] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[15]$_DFF_P_  (.D(_06610_),
    .Q(\hash.CA2.e_dash[15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[16]$_DFF_P_  (.D(\hash.CA1.S1.X[16] ),
    .Q(\hash.CA2.e_dash[16] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[17]$_DFF_P_  (.D(\hash.CA1.S1.X[17] ),
    .Q(\hash.CA2.e_dash[17] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[18]$_DFF_P_  (.D(\hash.CA1.S1.X[18] ),
    .Q(\hash.CA2.e_dash[18] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[19]$_DFF_P_  (.D(\hash.CA1.S1.X[19] ),
    .Q(\hash.CA2.e_dash[19] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[1]$_DFF_P_  (.D(\hash.CA1.S1.X[1] ),
    .Q(\hash.CA2.e_dash[1] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[20]$_DFF_P_  (.D(\hash.CA1.S1.X[20] ),
    .Q(\hash.CA2.e_dash[20] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[21]$_DFF_P_  (.D(\hash.CA1.S1.X[21] ),
    .Q(\hash.CA2.e_dash[21] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[22]$_DFF_P_  (.D(\hash.CA1.S1.X[22] ),
    .Q(\hash.CA2.e_dash[22] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[23]$_DFF_P_  (.D(\hash.CA1.S1.X[23] ),
    .Q(\hash.CA2.e_dash[23] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[24]$_DFF_P_  (.D(\hash.CA1.S1.X[24] ),
    .Q(\hash.CA2.e_dash[24] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[25]$_DFF_P_  (.D(net1053),
    .Q(\hash.CA2.e_dash[25] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[26]$_DFF_P_  (.D(net1054),
    .Q(\hash.CA2.e_dash[26] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[27]$_DFF_P_  (.D(_06699_),
    .Q(\hash.CA2.e_dash[27] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[28]$_DFF_P_  (.D(_06707_),
    .Q(\hash.CA2.e_dash[28] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[29]$_DFF_P_  (.D(\hash.CA1.S1.X[29] ),
    .Q(\hash.CA2.e_dash[29] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[2]$_DFF_P_  (.D(\hash.CA1.S1.X[2] ),
    .Q(\hash.CA2.e_dash[2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[30]$_DFF_P_  (.D(net1046),
    .Q(\hash.CA2.e_dash[30] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[31]$_DFF_P_  (.D(\hash.CA1.S1.X[31] ),
    .Q(\hash.CA2.e_dash[31] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[3]$_DFF_P_  (.D(\hash.CA1.S1.X[3] ),
    .Q(\hash.CA2.e_dash[3] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[4]$_DFF_P_  (.D(\hash.CA1.S1.X[4] ),
    .Q(\hash.CA2.e_dash[4] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[5]$_DFF_P_  (.D(\hash.CA1.S1.X[5] ),
    .Q(\hash.CA2.e_dash[5] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[6]$_DFF_P_  (.D(\hash.CA1.S1.X[6] ),
    .Q(\hash.CA2.e_dash[6] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[7]$_DFF_P_  (.D(\hash.CA1.S1.X[7] ),
    .Q(\hash.CA2.e_dash[7] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[8]$_DFF_P_  (.D(_06552_),
    .Q(\hash.CA2.e_dash[8] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[9]$_DFF_P_  (.D(\hash.CA1.S1.X[9] ),
    .Q(\hash.CA2.e_dash[9] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[0]$_DFF_P_  (.D(\hash.CA1.f[0] ),
    .Q(\hash.CA2.f_dash[0] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[10]$_DFF_P_  (.D(\hash.CA1.f[10] ),
    .Q(\hash.CA2.f_dash[10] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[11]$_DFF_P_  (.D(\hash.CA1.f[11] ),
    .Q(\hash.CA2.f_dash[11] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[12]$_DFF_P_  (.D(\hash.CA1.f[12] ),
    .Q(\hash.CA2.f_dash[12] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[13]$_DFF_P_  (.D(\hash.CA1.f[13] ),
    .Q(\hash.CA2.f_dash[13] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[14]$_DFF_P_  (.D(\hash.CA1.f[14] ),
    .Q(\hash.CA2.f_dash[14] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[15]$_DFF_P_  (.D(\hash.CA1.f[15] ),
    .Q(\hash.CA2.f_dash[15] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[16]$_DFF_P_  (.D(\hash.CA1.f[16] ),
    .Q(\hash.CA2.f_dash[16] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[17]$_DFF_P_  (.D(\hash.CA1.f[17] ),
    .Q(\hash.CA2.f_dash[17] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[18]$_DFF_P_  (.D(_06467_),
    .Q(\hash.CA2.f_dash[18] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[19]$_DFF_P_  (.D(\hash.CA1.f[19] ),
    .Q(\hash.CA2.f_dash[19] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[1]$_DFF_P_  (.D(\hash.CA1.f[1] ),
    .Q(\hash.CA2.f_dash[1] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[20]$_DFF_P_  (.D(\hash.CA1.f[20] ),
    .Q(\hash.CA2.f_dash[20] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[21]$_DFF_P_  (.D(\hash.CA1.f[21] ),
    .Q(\hash.CA2.f_dash[21] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[22]$_DFF_P_  (.D(\hash.CA1.f[22] ),
    .Q(\hash.CA2.f_dash[22] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[23]$_DFF_P_  (.D(\hash.CA1.f[23] ),
    .Q(\hash.CA2.f_dash[23] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[24]$_DFF_P_  (.D(_06487_),
    .Q(\hash.CA2.f_dash[24] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[25]$_DFF_P_  (.D(\hash.CA1.f[25] ),
    .Q(\hash.CA2.f_dash[25] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[26]$_DFF_P_  (.D(\hash.CA1.f[26] ),
    .Q(\hash.CA2.f_dash[26] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[27]$_DFF_P_  (.D(\hash.CA1.f[27] ),
    .Q(\hash.CA2.f_dash[27] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[28]$_DFF_P_  (.D(\hash.CA1.f[28] ),
    .Q(\hash.CA2.f_dash[28] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[29]$_DFF_P_  (.D(\hash.CA1.f[29] ),
    .Q(\hash.CA2.f_dash[29] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[2]$_DFF_P_  (.D(\hash.CA1.f[2] ),
    .Q(\hash.CA2.f_dash[2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[30]$_DFF_P_  (.D(\hash.CA1.f[30] ),
    .Q(\hash.CA2.f_dash[30] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[31]$_DFF_P_  (.D(\hash.CA1.f[31] ),
    .Q(\hash.CA2.f_dash[31] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[3]$_DFF_P_  (.D(\hash.CA1.f[3] ),
    .Q(\hash.CA2.f_dash[3] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[4]$_DFF_P_  (.D(\hash.CA1.f[4] ),
    .Q(\hash.CA2.f_dash[4] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[5]$_DFF_P_  (.D(\hash.CA1.f[5] ),
    .Q(\hash.CA2.f_dash[5] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[6]$_DFF_P_  (.D(\hash.CA1.f[6] ),
    .Q(\hash.CA2.f_dash[6] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[7]$_DFF_P_  (.D(\hash.CA1.f[7] ),
    .Q(\hash.CA2.f_dash[7] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[8]$_DFF_P_  (.D(\hash.CA1.f[8] ),
    .Q(\hash.CA2.f_dash[8] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[9]$_DFF_P_  (.D(_06438_),
    .Q(\hash.CA2.f_dash[9] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[0]$_DFFE_PN_  (.D(_00658_),
    .DE(_00906_),
    .Q(net923),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[10]$_DFFE_PN_  (.D(_00659_),
    .DE(_00906_),
    .Q(net934),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[11]$_DFFE_PN_  (.D(_00660_),
    .DE(_00906_),
    .Q(net935),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[12]$_DFFE_PN_  (.D(_00661_),
    .DE(_00906_),
    .Q(net936),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[13]$_DFFE_PN_  (.D(_00662_),
    .DE(_00906_),
    .Q(net937),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[14]$_DFFE_PN_  (.D(_00663_),
    .DE(_00906_),
    .Q(net938),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[15]$_DFFE_PN_  (.D(_00664_),
    .DE(_00906_),
    .Q(net939),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[16]$_DFFE_PN_  (.D(_00665_),
    .DE(_00906_),
    .Q(net941),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[17]$_DFFE_PN_  (.D(_00666_),
    .DE(_00906_),
    .Q(net942),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[18]$_DFFE_PN_  (.D(_00667_),
    .DE(_00906_),
    .Q(net943),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[19]$_DFFE_PN_  (.D(_00668_),
    .DE(_00906_),
    .Q(net944),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[1]$_DFFE_PN_  (.D(_00669_),
    .DE(_00906_),
    .Q(net924),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[20]$_DFFE_PN_  (.D(_00670_),
    .DE(_00906_),
    .Q(net945),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[21]$_DFFE_PN_  (.D(_00671_),
    .DE(_00906_),
    .Q(net946),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[22]$_DFFE_PN_  (.D(_00672_),
    .DE(_00906_),
    .Q(net947),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[23]$_DFFE_PN_  (.D(_00673_),
    .DE(_00906_),
    .Q(net948),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[24]$_DFFE_PN_  (.D(_00674_),
    .DE(_00906_),
    .Q(net949),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[25]$_DFFE_PN_  (.D(_00675_),
    .DE(_00906_),
    .Q(net950),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[26]$_DFFE_PN_  (.D(_00676_),
    .DE(_00906_),
    .Q(net952),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[27]$_DFFE_PN_  (.D(_00677_),
    .DE(_00906_),
    .Q(net953),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[28]$_DFFE_PN_  (.D(_00678_),
    .DE(_00906_),
    .Q(net954),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[29]$_DFFE_PN_  (.D(_00679_),
    .DE(_00906_),
    .Q(net955),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[2]$_DFFE_PN_  (.D(_00680_),
    .DE(_00906_),
    .Q(net925),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[30]$_DFFE_PN_  (.D(_00681_),
    .DE(_00906_),
    .Q(net956),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[31]$_DFFE_PN_  (.D(_00682_),
    .DE(_00906_),
    .Q(net957),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[3]$_DFFE_PN_  (.D(_00683_),
    .DE(_00906_),
    .Q(net926),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[4]$_DFFE_PN_  (.D(_00684_),
    .DE(_00906_),
    .Q(net927),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[5]$_DFFE_PN_  (.D(_00685_),
    .DE(_00906_),
    .Q(net928),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[6]$_DFFE_PN_  (.D(_00686_),
    .DE(_00906_),
    .Q(net930),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[7]$_DFFE_PN_  (.D(_00687_),
    .DE(_00906_),
    .Q(net931),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[8]$_DFFE_PN_  (.D(_00688_),
    .DE(_00906_),
    .Q(net932),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[9]$_DFFE_PN_  (.D(_00689_),
    .DE(_00906_),
    .Q(net933),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[0]$_DFFE_PN_  (.D(_00690_),
    .DE(_00906_),
    .Q(net887),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[10]$_DFFE_PN_  (.D(_00691_),
    .DE(_00906_),
    .Q(net899),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[11]$_DFFE_PN_  (.D(_00692_),
    .DE(_00906_),
    .Q(net900),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[12]$_DFFE_PN_  (.D(_00693_),
    .DE(_00906_),
    .Q(net901),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[13]$_DFFE_PN_  (.D(_00694_),
    .DE(_00906_),
    .Q(net902),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[14]$_DFFE_PN_  (.D(_00695_),
    .DE(_00906_),
    .Q(net903),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[15]$_DFFE_PN_  (.D(_00696_),
    .DE(_00906_),
    .Q(net904),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[16]$_DFFE_PN_  (.D(_00697_),
    .DE(_00906_),
    .Q(net905),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[17]$_DFFE_PN_  (.D(_00698_),
    .DE(_00906_),
    .Q(net906),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[18]$_DFFE_PN_  (.D(_00699_),
    .DE(_00906_),
    .Q(net908),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[19]$_DFFE_PN_  (.D(_00700_),
    .DE(_00906_),
    .Q(net909),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[1]$_DFFE_PN_  (.D(_11575_),
    .DE(_00906_),
    .Q(net888),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[20]$_DFFE_PN_  (.D(_00701_),
    .DE(_00906_),
    .Q(net910),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[21]$_DFFE_PN_  (.D(_00702_),
    .DE(_00906_),
    .Q(net911),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[22]$_DFFE_PN_  (.D(_00703_),
    .DE(_00906_),
    .Q(net912),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[23]$_DFFE_PN_  (.D(_00704_),
    .DE(_00906_),
    .Q(net913),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[24]$_DFFE_PN_  (.D(_00705_),
    .DE(_00906_),
    .Q(net914),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[25]$_DFFE_PN_  (.D(_00706_),
    .DE(_00906_),
    .Q(net915),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[26]$_DFFE_PN_  (.D(_00707_),
    .DE(_00906_),
    .Q(net916),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[27]$_DFFE_PN_  (.D(_00708_),
    .DE(_00906_),
    .Q(net917),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[28]$_DFFE_PN_  (.D(_00709_),
    .DE(_00906_),
    .Q(net919),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[29]$_DFFE_PN_  (.D(_00710_),
    .DE(_00906_),
    .Q(net920),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[2]$_DFFE_PN_  (.D(_00711_),
    .DE(_00906_),
    .Q(net889),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[30]$_DFFE_PN_  (.D(_00712_),
    .DE(_00906_),
    .Q(net921),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[31]$_DFFE_PN_  (.D(_00713_),
    .DE(_00906_),
    .Q(net922),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[3]$_DFFE_PN_  (.D(_00714_),
    .DE(_00906_),
    .Q(net890),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[4]$_DFFE_PN_  (.D(_00715_),
    .DE(_00906_),
    .Q(net891),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[5]$_DFFE_PN_  (.D(_00716_),
    .DE(_00906_),
    .Q(net892),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[6]$_DFFE_PN_  (.D(_00717_),
    .DE(_00906_),
    .Q(net893),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[7]$_DFFE_PN_  (.D(_00718_),
    .DE(_00906_),
    .Q(net894),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[8]$_DFFE_PN_  (.D(_00719_),
    .DE(_00906_),
    .Q(net897),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[9]$_DFFE_PN_  (.D(_00720_),
    .DE(_00906_),
    .Q(net898),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[0]$_DFFE_PN_  (.D(\hash.CA1.c[0] ),
    .DE(_00906_),
    .Q(net852),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[10]$_DFFE_PN_  (.D(_00750_),
    .DE(_00906_),
    .Q(net863),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[11]$_DFFE_PN_  (.D(_00722_),
    .DE(_00906_),
    .Q(net864),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[12]$_DFFE_PN_  (.D(_00723_),
    .DE(_00906_),
    .Q(net865),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[13]$_DFFE_PN_  (.D(_00724_),
    .DE(_00906_),
    .Q(net866),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[14]$_DFFE_PN_  (.D(_00725_),
    .DE(_00906_),
    .Q(net867),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[15]$_DFFE_PN_  (.D(_00726_),
    .DE(_00906_),
    .Q(net868),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[16]$_DFFE_PN_  (.D(_00727_),
    .DE(_00906_),
    .Q(net869),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[17]$_DFFE_PN_  (.D(_00728_),
    .DE(_00906_),
    .Q(net870),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[18]$_DFFE_PN_  (.D(_00729_),
    .DE(_00906_),
    .Q(net871),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[19]$_DFFE_PN_  (.D(_00730_),
    .DE(_00906_),
    .Q(net872),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[1]$_DFFE_PN_  (.D(_00721_),
    .DE(_00906_),
    .Q(net853),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[20]$_DFFE_PN_  (.D(_00731_),
    .DE(_00906_),
    .Q(net874),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[21]$_DFFE_PN_  (.D(_00732_),
    .DE(_00906_),
    .Q(net875),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[22]$_DFFE_PN_  (.D(_00733_),
    .DE(_00906_),
    .Q(net876),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[23]$_DFFE_PN_  (.D(_00734_),
    .DE(_00906_),
    .Q(net877),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[24]$_DFFE_PN_  (.D(_00735_),
    .DE(_00906_),
    .Q(net878),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[25]$_DFFE_PN_  (.D(_00736_),
    .DE(_00906_),
    .Q(net879),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[26]$_DFFE_PN_  (.D(_00737_),
    .DE(_00906_),
    .Q(net880),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[27]$_DFFE_PN_  (.D(_00738_),
    .DE(_00906_),
    .Q(net881),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[28]$_DFFE_PN_  (.D(_00739_),
    .DE(_00906_),
    .Q(net882),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[29]$_DFFE_PN_  (.D(_00740_),
    .DE(_00906_),
    .Q(net883),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[2]$_DFFE_PN_  (.D(_11576_),
    .DE(_00906_),
    .Q(net854),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[30]$_DFFE_PN_  (.D(_00741_),
    .DE(_00906_),
    .Q(net885),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[31]$_DFFE_PN_  (.D(_00743_),
    .DE(_00906_),
    .Q(net886),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[3]$_DFFE_PN_  (.D(_00742_),
    .DE(_00906_),
    .Q(net855),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[4]$_DFFE_PN_  (.D(_00744_),
    .DE(_00906_),
    .Q(net856),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[5]$_DFFE_PN_  (.D(_00745_),
    .DE(_00906_),
    .Q(net857),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[6]$_DFFE_PN_  (.D(_00746_),
    .DE(_00906_),
    .Q(net858),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[7]$_DFFE_PN_  (.D(_00747_),
    .DE(_00906_),
    .Q(net859),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[8]$_DFFE_PN_  (.D(_00748_),
    .DE(_00906_),
    .Q(net860),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[9]$_DFFE_PN_  (.D(_00749_),
    .DE(_00906_),
    .Q(net861),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[0]$_DFFE_PN_  (.D(\hash.CA1.d[0] ),
    .DE(_00906_),
    .Q(net816),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[10]$_DFFE_PN_  (.D(_00780_),
    .DE(_00906_),
    .Q(net827),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[11]$_DFFE_PN_  (.D(_00752_),
    .DE(_00906_),
    .Q(net828),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[12]$_DFFE_PN_  (.D(_00753_),
    .DE(_00906_),
    .Q(net830),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[13]$_DFFE_PN_  (.D(_00754_),
    .DE(_00906_),
    .Q(net831),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[14]$_DFFE_PN_  (.D(_00755_),
    .DE(_00906_),
    .Q(net832),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[15]$_DFFE_PN_  (.D(_00756_),
    .DE(_00906_),
    .Q(net833),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[16]$_DFFE_PN_  (.D(_00757_),
    .DE(_00906_),
    .Q(net834),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[17]$_DFFE_PN_  (.D(_00758_),
    .DE(_00906_),
    .Q(net835),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[18]$_DFFE_PN_  (.D(_00759_),
    .DE(_00906_),
    .Q(net836),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[19]$_DFFE_PN_  (.D(_00760_),
    .DE(_00906_),
    .Q(net837),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[1]$_DFFE_PN_  (.D(_00751_),
    .DE(_00906_),
    .Q(net817),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[20]$_DFFE_PN_  (.D(_00761_),
    .DE(_00906_),
    .Q(net838),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[21]$_DFFE_PN_  (.D(_00762_),
    .DE(_00906_),
    .Q(net839),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[22]$_DFFE_PN_  (.D(_00763_),
    .DE(_00906_),
    .Q(net841),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[23]$_DFFE_PN_  (.D(_00764_),
    .DE(_00906_),
    .Q(net842),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[24]$_DFFE_PN_  (.D(_00765_),
    .DE(_00906_),
    .Q(net843),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[25]$_DFFE_PN_  (.D(_00766_),
    .DE(_00906_),
    .Q(net844),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[26]$_DFFE_PN_  (.D(_00767_),
    .DE(_00906_),
    .Q(net845),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[27]$_DFFE_PN_  (.D(_00768_),
    .DE(_00906_),
    .Q(net846),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[28]$_DFFE_PN_  (.D(_00769_),
    .DE(_00906_),
    .Q(net847),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[29]$_DFFE_PN_  (.D(_00770_),
    .DE(_00906_),
    .Q(net848),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[2]$_DFFE_PN_  (.D(_11577_),
    .DE(_00906_),
    .Q(net819),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[30]$_DFFE_PN_  (.D(_00771_),
    .DE(_00906_),
    .Q(net849),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[31]$_DFFE_PN_  (.D(_00773_),
    .DE(_00906_),
    .Q(net850),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[3]$_DFFE_PN_  (.D(_00772_),
    .DE(_00906_),
    .Q(net820),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[4]$_DFFE_PN_  (.D(_00774_),
    .DE(_00906_),
    .Q(net821),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[5]$_DFFE_PN_  (.D(_00775_),
    .DE(_00906_),
    .Q(net822),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[6]$_DFFE_PN_  (.D(_00776_),
    .DE(_00906_),
    .Q(net823),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[7]$_DFFE_PN_  (.D(_00777_),
    .DE(_00906_),
    .Q(net824),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[8]$_DFFE_PN_  (.D(_00778_),
    .DE(_00906_),
    .Q(net825),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[9]$_DFFE_PN_  (.D(_00779_),
    .DE(_00906_),
    .Q(net826),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[0]$_DFFE_PN_  (.D(_00781_),
    .DE(_00906_),
    .Q(net1036),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[10]$_DFFE_PN_  (.D(_00782_),
    .DE(_00906_),
    .Q(net792),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[11]$_DFFE_PN_  (.D(_00783_),
    .DE(_00906_),
    .Q(net793),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[12]$_DFFE_PN_  (.D(_00784_),
    .DE(_00906_),
    .Q(net794),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[13]$_DFFE_PN_  (.D(_00785_),
    .DE(_00906_),
    .Q(net795),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[14]$_DFFE_PN_  (.D(_00786_),
    .DE(_00906_),
    .Q(net797),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[15]$_DFFE_PN_  (.D(_00787_),
    .DE(_00906_),
    .Q(net798),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[16]$_DFFE_PN_  (.D(_00788_),
    .DE(_00906_),
    .Q(net799),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[17]$_DFFE_PN_  (.D(_00789_),
    .DE(_00906_),
    .Q(net800),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[18]$_DFFE_PN_  (.D(_00790_),
    .DE(_00906_),
    .Q(net801),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[19]$_DFFE_PN_  (.D(_00791_),
    .DE(_00906_),
    .Q(net802),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[1]$_DFFE_PN_  (.D(_00792_),
    .DE(_00906_),
    .Q(net1037),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[20]$_DFFE_PN_  (.D(_00793_),
    .DE(_00906_),
    .Q(net803),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[21]$_DFFE_PN_  (.D(_00794_),
    .DE(_00906_),
    .Q(net804),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[22]$_DFFE_PN_  (.D(_00795_),
    .DE(_00906_),
    .Q(net805),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[23]$_DFFE_PN_  (.D(_00796_),
    .DE(_00906_),
    .Q(net806),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[24]$_DFFE_PN_  (.D(_00797_),
    .DE(_00906_),
    .Q(net808),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[25]$_DFFE_PN_  (.D(_00798_),
    .DE(_00906_),
    .Q(net809),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[26]$_DFFE_PN_  (.D(_00799_),
    .DE(_00906_),
    .Q(net810),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[27]$_DFFE_PN_  (.D(_00800_),
    .DE(_00906_),
    .Q(net811),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[28]$_DFFE_PN_  (.D(_00801_),
    .DE(_00906_),
    .Q(net812),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[29]$_DFFE_PN_  (.D(_00802_),
    .DE(_00906_),
    .Q(net813),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[2]$_DFFE_PN_  (.D(_00803_),
    .DE(_00906_),
    .Q(net1038),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[30]$_DFFE_PN_  (.D(_00804_),
    .DE(_00906_),
    .Q(net814),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[31]$_DFFE_PN_  (.D(_00805_),
    .DE(_00906_),
    .Q(net815),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[3]$_DFFE_PN_  (.D(_00806_),
    .DE(_00906_),
    .Q(net1039),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[4]$_DFFE_PN_  (.D(_00807_),
    .DE(_00906_),
    .Q(net786),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[5]$_DFFE_PN_  (.D(_00808_),
    .DE(_00906_),
    .Q(net787),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[6]$_DFFE_PN_  (.D(_00809_),
    .DE(_00906_),
    .Q(net788),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[7]$_DFFE_PN_  (.D(_00810_),
    .DE(_00906_),
    .Q(net789),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[8]$_DFFE_PN_  (.D(_00811_),
    .DE(_00906_),
    .Q(net790),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[9]$_DFFE_PN_  (.D(_00812_),
    .DE(_00906_),
    .Q(net791),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[0]$_DFFE_PN_  (.D(\hash.CA1.f[0] ),
    .DE(_00906_),
    .Q(net1001),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[10]$_DFFE_PN_  (.D(_00841_),
    .DE(_00906_),
    .Q(net1012),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[11]$_DFFE_PN_  (.D(_00842_),
    .DE(_00906_),
    .Q(net1013),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[12]$_DFFE_PN_  (.D(_00814_),
    .DE(_00906_),
    .Q(net1014),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[13]$_DFFE_PN_  (.D(_00815_),
    .DE(_00906_),
    .Q(net1015),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[14]$_DFFE_PN_  (.D(_00816_),
    .DE(_00906_),
    .Q(net1016),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[15]$_DFFE_PN_  (.D(_00817_),
    .DE(_00906_),
    .Q(net1017),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[16]$_DFFE_PN_  (.D(_00818_),
    .DE(_00906_),
    .Q(net1019),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[17]$_DFFE_PN_  (.D(_00819_),
    .DE(_00906_),
    .Q(net1020),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[18]$_DFFE_PN_  (.D(_00820_),
    .DE(_00906_),
    .Q(net1021),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[19]$_DFFE_PN_  (.D(_00821_),
    .DE(_00906_),
    .Q(net1022),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[1]$_DFFE_PN_  (.D(\hash.CA1.f[1] ),
    .DE(_00906_),
    .Q(net1002),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[20]$_DFFE_PN_  (.D(_00822_),
    .DE(_00906_),
    .Q(net1023),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[21]$_DFFE_PN_  (.D(_00823_),
    .DE(_00906_),
    .Q(net1024),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[22]$_DFFE_PN_  (.D(_00825_),
    .DE(_00906_),
    .Q(net1025),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[23]$_DFFE_PN_  (.D(_00826_),
    .DE(_00906_),
    .Q(net1026),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[24]$_DFFE_PN_  (.D(_00827_),
    .DE(_00906_),
    .Q(net1027),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[25]$_DFFE_PN_  (.D(_00828_),
    .DE(_00906_),
    .Q(net1028),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[26]$_DFFE_PN_  (.D(_00829_),
    .DE(_00906_),
    .Q(net1030),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[27]$_DFFE_PN_  (.D(_00830_),
    .DE(_00906_),
    .Q(net1031),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[28]$_DFFE_PN_  (.D(_00831_),
    .DE(_00906_),
    .Q(net1032),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[29]$_DFFE_PN_  (.D(_00832_),
    .DE(_00906_),
    .Q(net1033),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[2]$_DFFE_PN_  (.D(_00813_),
    .DE(_00906_),
    .Q(net1003),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[30]$_DFFE_PN_  (.D(_00833_),
    .DE(_00906_),
    .Q(net1034),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[31]$_DFFE_PN_  (.D(_00834_),
    .DE(_00906_),
    .Q(net1035),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[3]$_DFFE_PN_  (.D(_00824_),
    .DE(_00906_),
    .Q(net1004),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[4]$_DFFE_PN_  (.D(_00835_),
    .DE(_00906_),
    .Q(net1005),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[5]$_DFFE_PN_  (.D(_00836_),
    .DE(_00906_),
    .Q(net1006),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[6]$_DFFE_PN_  (.D(_00837_),
    .DE(_00906_),
    .Q(net1008),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[7]$_DFFE_PN_  (.D(_00838_),
    .DE(_00906_),
    .Q(net1009),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[8]$_DFFE_PN_  (.D(_00839_),
    .DE(_00906_),
    .Q(net1010),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[9]$_DFFE_PN_  (.D(_00840_),
    .DE(_00906_),
    .Q(net1011),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[0]$_DFFE_PN_  (.D(_00843_),
    .DE(_00906_),
    .Q(net966),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[10]$_DFFE_PN_  (.D(_00844_),
    .DE(_00906_),
    .Q(net977),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[11]$_DFFE_PN_  (.D(_00845_),
    .DE(_00906_),
    .Q(net978),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[12]$_DFFE_PN_  (.D(_00846_),
    .DE(_00906_),
    .Q(net979),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[13]$_DFFE_PN_  (.D(_00847_),
    .DE(_00906_),
    .Q(net980),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[14]$_DFFE_PN_  (.D(_00848_),
    .DE(_00906_),
    .Q(net981),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[15]$_DFFE_PN_  (.D(_00849_),
    .DE(_00906_),
    .Q(net982),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[16]$_DFFE_PN_  (.D(_00850_),
    .DE(_00906_),
    .Q(net983),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[17]$_DFFE_PN_  (.D(_00851_),
    .DE(_00906_),
    .Q(net984),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[18]$_DFFE_PN_  (.D(_00852_),
    .DE(_00906_),
    .Q(net986),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[19]$_DFFE_PN_  (.D(_00853_),
    .DE(_00906_),
    .Q(net987),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[1]$_DFFE_PN_  (.D(_00854_),
    .DE(_00906_),
    .Q(net967),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[20]$_DFFE_PN_  (.D(_00855_),
    .DE(_00906_),
    .Q(net988),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[21]$_DFFE_PN_  (.D(_00856_),
    .DE(_00906_),
    .Q(net989),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[22]$_DFFE_PN_  (.D(_00857_),
    .DE(_00906_),
    .Q(net990),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[23]$_DFFE_PN_  (.D(_00858_),
    .DE(_00906_),
    .Q(net991),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[24]$_DFFE_PN_  (.D(_00859_),
    .DE(_00906_),
    .Q(net992),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[25]$_DFFE_PN_  (.D(_00860_),
    .DE(_00906_),
    .Q(net993),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[26]$_DFFE_PN_  (.D(_00861_),
    .DE(_00906_),
    .Q(net994),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[27]$_DFFE_PN_  (.D(_00862_),
    .DE(_00906_),
    .Q(net995),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[28]$_DFFE_PN_  (.D(_00863_),
    .DE(_00906_),
    .Q(net997),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[29]$_DFFE_PN_  (.D(_00864_),
    .DE(_00906_),
    .Q(net998),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[2]$_DFFE_PN_  (.D(_00865_),
    .DE(_00906_),
    .Q(net968),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[30]$_DFFE_PN_  (.D(_00866_),
    .DE(_00906_),
    .Q(net999),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[31]$_DFFE_PN_  (.D(_00867_),
    .DE(_00906_),
    .Q(net1000),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[3]$_DFFE_PN_  (.D(_00868_),
    .DE(_00906_),
    .Q(net969),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[4]$_DFFE_PN_  (.D(_00869_),
    .DE(_00906_),
    .Q(net970),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[5]$_DFFE_PN_  (.D(_00870_),
    .DE(_00906_),
    .Q(net971),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[6]$_DFFE_PN_  (.D(_00871_),
    .DE(_00906_),
    .Q(net972),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[7]$_DFFE_PN_  (.D(_00872_),
    .DE(_00906_),
    .Q(net973),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[8]$_DFFE_PN_  (.D(_00873_),
    .DE(_00906_),
    .Q(net975),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[9]$_DFFE_PN_  (.D(_00874_),
    .DE(_00906_),
    .Q(net976),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[0]$_DFFE_PN_  (.D(_00875_),
    .DE(_00906_),
    .Q(net785),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[10]$_DFFE_PN_  (.D(_00876_),
    .DE(_00906_),
    .Q(net796),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[11]$_DFFE_PN_  (.D(_00877_),
    .DE(_00906_),
    .Q(net807),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[12]$_DFFE_PN_  (.D(_00878_),
    .DE(_00906_),
    .Q(net818),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[13]$_DFFE_PN_  (.D(_00879_),
    .DE(_00906_),
    .Q(net829),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[14]$_DFFE_PN_  (.D(_00880_),
    .DE(_00906_),
    .Q(net840),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[15]$_DFFE_PN_  (.D(_00881_),
    .DE(_00906_),
    .Q(net851),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[16]$_DFFE_PN_  (.D(_00882_),
    .DE(_00906_),
    .Q(net862),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[17]$_DFFE_PN_  (.D(_00883_),
    .DE(_00906_),
    .Q(net873),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[18]$_DFFE_PN_  (.D(_00884_),
    .DE(_00906_),
    .Q(net884),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[19]$_DFFE_PN_  (.D(_00885_),
    .DE(_00906_),
    .Q(net895),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[1]$_DFFE_PN_  (.D(_11578_),
    .DE(_00906_),
    .Q(net896),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[20]$_DFFE_PN_  (.D(_00886_),
    .DE(_00906_),
    .Q(net907),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[21]$_DFFE_PN_  (.D(_00887_),
    .DE(_00906_),
    .Q(net918),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[22]$_DFFE_PN_  (.D(_00888_),
    .DE(_00906_),
    .Q(net929),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[23]$_DFFE_PN_  (.D(_00889_),
    .DE(_00906_),
    .Q(net940),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[24]$_DFFE_PN_  (.D(_00890_),
    .DE(_00906_),
    .Q(net951),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[25]$_DFFE_PN_  (.D(_00891_),
    .DE(_00906_),
    .Q(net958),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[26]$_DFFE_PN_  (.D(_00892_),
    .DE(_00906_),
    .Q(net959),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[27]$_DFFE_PN_  (.D(_00893_),
    .DE(_00906_),
    .Q(net960),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[28]$_DFFE_PN_  (.D(_00894_),
    .DE(_00906_),
    .Q(net961),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[29]$_DFFE_PN_  (.D(_00895_),
    .DE(_00906_),
    .Q(net962),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[2]$_DFFE_PN_  (.D(_00896_),
    .DE(_00906_),
    .Q(net963),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[30]$_DFFE_PN_  (.D(_00897_),
    .DE(_00906_),
    .Q(net964),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[31]$_DFFE_PN_  (.D(_00898_),
    .DE(_00906_),
    .Q(net965),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[3]$_DFFE_PN_  (.D(_00899_),
    .DE(_00906_),
    .Q(net974),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[4]$_DFFE_PN_  (.D(_00900_),
    .DE(_00906_),
    .Q(net985),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[5]$_DFFE_PN_  (.D(_00901_),
    .DE(_00906_),
    .Q(net996),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[6]$_DFFE_PN_  (.D(_00902_),
    .DE(_00906_),
    .Q(net1007),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[7]$_DFFE_PN_  (.D(_00903_),
    .DE(_00906_),
    .Q(net1018),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[8]$_DFFE_PN_  (.D(_00904_),
    .DE(_00906_),
    .Q(net1029),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[9]$_DFFE_PN_  (.D(_00905_),
    .DE(_00906_),
    .Q(net1040),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p1_cap[0]$_DFF_P_  (.D(\hash.CA1.p1[0] ),
    .Q(\hash.CA2.p1[0] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[10]$_DFF_P_  (.D(\hash.CA1.p1[10] ),
    .Q(\hash.CA2.p1[10] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[11]$_DFF_P_  (.D(\hash.CA1.p1[11] ),
    .Q(\hash.CA2.p1[11] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[12]$_DFF_P_  (.D(\hash.CA1.p1[12] ),
    .Q(\hash.CA2.p1[12] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[13]$_DFF_P_  (.D(\hash.CA1.p1[13] ),
    .Q(\hash.CA2.p1[13] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[14]$_DFF_P_  (.D(\hash.CA1.p1[14] ),
    .Q(\hash.CA2.p1[14] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[15]$_DFF_P_  (.D(\hash.CA1.p1[15] ),
    .Q(\hash.CA2.p1[15] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[16]$_DFF_P_  (.D(\hash.CA1.p1[16] ),
    .Q(\hash.CA2.p1[16] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[17]$_DFF_P_  (.D(\hash.CA1.p1[17] ),
    .Q(\hash.CA2.p1[17] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[18]$_DFF_P_  (.D(\hash.CA1.p1[18] ),
    .Q(\hash.CA2.p1[18] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[19]$_DFF_P_  (.D(\hash.CA1.p1[19] ),
    .Q(\hash.CA2.p1[19] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[1]$_DFF_P_  (.D(\hash.CA1.p1[1] ),
    .Q(\hash.CA2.p1[1] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[20]$_DFF_P_  (.D(\hash.CA1.p1[20] ),
    .Q(\hash.CA2.p1[20] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[21]$_DFF_P_  (.D(\hash.CA1.p1[21] ),
    .Q(\hash.CA2.p1[21] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[22]$_DFF_P_  (.D(\hash.CA1.p1[22] ),
    .Q(\hash.CA2.p1[22] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[23]$_DFF_P_  (.D(\hash.CA1.p1[23] ),
    .Q(\hash.CA2.p1[23] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[24]$_DFF_P_  (.D(\hash.CA1.p1[24] ),
    .Q(\hash.CA2.p1[24] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[25]$_DFF_P_  (.D(\hash.CA1.p1[25] ),
    .Q(\hash.CA2.p1[25] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[26]$_DFF_P_  (.D(\hash.CA1.p1[26] ),
    .Q(\hash.CA2.p1[26] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[27]$_DFF_P_  (.D(\hash.CA1.p1[27] ),
    .Q(\hash.CA2.p1[27] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[28]$_DFF_P_  (.D(\hash.CA1.p1[28] ),
    .Q(\hash.CA2.p1[28] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[29]$_DFF_P_  (.D(\hash.CA1.p1[29] ),
    .Q(\hash.CA2.p1[29] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[2]$_DFF_P_  (.D(\hash.CA1.p1[2] ),
    .Q(\hash.CA2.p1[2] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[30]$_DFF_P_  (.D(\hash.CA1.p1[30] ),
    .Q(\hash.CA2.p1[30] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[31]$_DFF_P_  (.D(\hash.CA1.p1[31] ),
    .Q(\hash.CA2.p1[31] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[3]$_DFF_P_  (.D(\hash.CA1.p1[3] ),
    .Q(\hash.CA2.p1[3] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[4]$_DFF_P_  (.D(\hash.CA1.p1[4] ),
    .Q(\hash.CA2.p1[4] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[5]$_DFF_P_  (.D(\hash.CA1.p1[5] ),
    .Q(\hash.CA2.p1[5] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[6]$_DFF_P_  (.D(\hash.CA1.p1[6] ),
    .Q(\hash.CA2.p1[6] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[7]$_DFF_P_  (.D(\hash.CA1.p1[7] ),
    .Q(\hash.CA2.p1[7] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[8]$_DFF_P_  (.D(\hash.CA1.p1[8] ),
    .Q(\hash.CA2.p1[8] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[9]$_DFF_P_  (.D(\hash.CA1.p1[9] ),
    .Q(\hash.CA2.p1[9] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[0]$_DFF_P_  (.D(\hash.CA1.p2[0] ),
    .Q(\hash.CA2.S1.X[0] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[10]$_DFF_P_  (.D(\hash.CA1.p2[10] ),
    .Q(\hash.CA2.S1.X[10] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[11]$_DFF_P_  (.D(\hash.CA1.p2[11] ),
    .Q(\hash.CA2.S1.X[11] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[12]$_DFF_P_  (.D(\hash.CA1.p2[12] ),
    .Q(\hash.CA2.S1.X[12] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[13]$_DFF_P_  (.D(\hash.CA1.p2[13] ),
    .Q(\hash.CA2.S1.X[13] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[14]$_DFF_P_  (.D(\hash.CA1.p2[14] ),
    .Q(\hash.CA2.S1.X[14] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[15]$_DFF_P_  (.D(\hash.CA1.p2[15] ),
    .Q(\hash.CA2.S1.X[15] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[16]$_DFF_P_  (.D(\hash.CA1.p2[16] ),
    .Q(\hash.CA2.S1.X[16] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[17]$_DFF_P_  (.D(\hash.CA1.p2[17] ),
    .Q(\hash.CA2.S1.X[17] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[18]$_DFF_P_  (.D(\hash.CA1.p2[18] ),
    .Q(\hash.CA2.S1.X[18] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[19]$_DFF_P_  (.D(\hash.CA1.p2[19] ),
    .Q(\hash.CA2.S1.X[19] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[1]$_DFF_P_  (.D(\hash.CA1.p2[1] ),
    .Q(\hash.CA2.S1.X[1] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[20]$_DFF_P_  (.D(\hash.CA1.p2[20] ),
    .Q(\hash.CA2.S1.X[20] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[21]$_DFF_P_  (.D(\hash.CA1.p2[21] ),
    .Q(\hash.CA2.S1.X[21] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[22]$_DFF_P_  (.D(\hash.CA1.p2[22] ),
    .Q(\hash.CA2.S1.X[22] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[23]$_DFF_P_  (.D(\hash.CA1.p2[23] ),
    .Q(\hash.CA2.S1.X[23] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[24]$_DFF_P_  (.D(\hash.CA1.p2[24] ),
    .Q(\hash.CA2.S1.X[24] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[25]$_DFF_P_  (.D(\hash.CA1.p2[25] ),
    .Q(\hash.CA2.S1.X[25] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[26]$_DFF_P_  (.D(\hash.CA1.p2[26] ),
    .Q(\hash.CA2.S1.X[26] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[27]$_DFF_P_  (.D(\hash.CA1.p2[27] ),
    .Q(\hash.CA2.S1.X[27] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[28]$_DFF_P_  (.D(\hash.CA1.p2[28] ),
    .Q(\hash.CA2.S1.X[28] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[29]$_DFF_P_  (.D(\hash.CA1.p2[29] ),
    .Q(\hash.CA2.S1.X[29] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[2]$_DFF_P_  (.D(\hash.CA1.p2[2] ),
    .Q(\hash.CA2.S1.X[2] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[30]$_DFF_P_  (.D(\hash.CA1.p2[30] ),
    .Q(\hash.CA2.S1.X[30] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[31]$_DFF_P_  (.D(\hash.CA1.p2[31] ),
    .Q(\hash.CA2.S1.X[31] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[3]$_DFF_P_  (.D(\hash.CA1.p2[3] ),
    .Q(\hash.CA2.S1.X[3] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[4]$_DFF_P_  (.D(\hash.CA1.p2[4] ),
    .Q(\hash.CA2.S1.X[4] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[5]$_DFF_P_  (.D(\hash.CA1.p2[5] ),
    .Q(\hash.CA2.S1.X[5] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[6]$_DFF_P_  (.D(\hash.CA1.p2[6] ),
    .Q(\hash.CA2.S1.X[6] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[7]$_DFF_P_  (.D(\hash.CA1.p2[7] ),
    .Q(\hash.CA2.S1.X[7] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[8]$_DFF_P_  (.D(\hash.CA1.p2[8] ),
    .Q(\hash.CA2.S1.X[8] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[9]$_DFF_P_  (.D(\hash.CA1.p2[9] ),
    .Q(\hash.CA2.S1.X[9] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p3_cap[0]$_DFF_P_  (.D(\hash.CA1.p3[0] ),
    .Q(\hash.CA2.p3[0] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[10]$_DFF_P_  (.D(\hash.CA1.p3[10] ),
    .Q(\hash.CA2.p3[10] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[11]$_DFF_P_  (.D(\hash.CA1.p3[11] ),
    .Q(\hash.CA2.p3[11] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[12]$_DFF_P_  (.D(\hash.CA1.p3[12] ),
    .Q(\hash.CA2.p3[12] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[13]$_DFF_P_  (.D(\hash.CA1.p3[13] ),
    .Q(\hash.CA2.p3[13] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[14]$_DFF_P_  (.D(\hash.CA1.p3[14] ),
    .Q(\hash.CA2.p3[14] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[15]$_DFF_P_  (.D(\hash.CA1.p3[15] ),
    .Q(\hash.CA2.p3[15] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p3_cap[16]$_DFF_P_  (.D(\hash.CA1.p3[16] ),
    .Q(\hash.CA2.p3[16] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p3_cap[17]$_DFF_P_  (.D(\hash.CA1.p3[17] ),
    .Q(\hash.CA2.p3[17] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[18]$_DFF_P_  (.D(\hash.CA1.p3[18] ),
    .Q(\hash.CA2.p3[18] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[19]$_DFF_P_  (.D(\hash.CA1.p3[19] ),
    .Q(\hash.CA2.p3[19] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[1]$_DFF_P_  (.D(\hash.CA1.p3[1] ),
    .Q(\hash.CA2.p3[1] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[20]$_DFF_P_  (.D(\hash.CA1.p3[20] ),
    .Q(\hash.CA2.p3[20] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[21]$_DFF_P_  (.D(\hash.CA1.p3[21] ),
    .Q(\hash.CA2.p3[21] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[22]$_DFF_P_  (.D(\hash.CA1.p3[22] ),
    .Q(\hash.CA2.p3[22] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[23]$_DFF_P_  (.D(\hash.CA1.p3[23] ),
    .Q(\hash.CA2.p3[23] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[24]$_DFF_P_  (.D(\hash.CA1.p3[24] ),
    .Q(\hash.CA2.p3[24] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[25]$_DFF_P_  (.D(\hash.CA1.p3[25] ),
    .Q(\hash.CA2.p3[25] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[26]$_DFF_P_  (.D(\hash.CA1.p3[26] ),
    .Q(\hash.CA2.p3[26] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[27]$_DFF_P_  (.D(\hash.CA1.p3[27] ),
    .Q(\hash.CA2.p3[27] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[28]$_DFF_P_  (.D(\hash.CA1.p3[28] ),
    .Q(\hash.CA2.p3[28] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[29]$_DFF_P_  (.D(\hash.CA1.p3[29] ),
    .Q(\hash.CA2.p3[29] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[2]$_DFF_P_  (.D(\hash.CA1.p3[2] ),
    .Q(\hash.CA2.p3[2] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[30]$_DFF_P_  (.D(\hash.CA1.p3[30] ),
    .Q(\hash.CA2.p3[30] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[31]$_DFF_P_  (.D(\hash.CA1.p3[31] ),
    .Q(\hash.CA2.p3[31] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[3]$_DFF_P_  (.D(\hash.CA1.p3[3] ),
    .Q(\hash.CA2.p3[3] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[4]$_DFF_P_  (.D(\hash.CA1.p3[4] ),
    .Q(\hash.CA2.p3[4] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[5]$_DFF_P_  (.D(\hash.CA1.p3[5] ),
    .Q(\hash.CA2.p3[5] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[6]$_DFF_P_  (.D(\hash.CA1.p3[6] ),
    .Q(\hash.CA2.p3[6] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[7]$_DFF_P_  (.D(\hash.CA1.p3[7] ),
    .Q(\hash.CA2.p3[7] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[8]$_DFF_P_  (.D(\hash.CA1.p3[8] ),
    .Q(\hash.CA2.p3[8] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[9]$_DFF_P_  (.D(\hash.CA1.p3[9] ),
    .Q(\hash.CA2.p3[9] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[0]$_DFF_P_  (.D(\hash.CA1.p4[0] ),
    .Q(\hash.CA2.p4[0] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[10]$_DFF_P_  (.D(\hash.CA1.p4[10] ),
    .Q(\hash.CA2.p4[10] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[11]$_DFF_P_  (.D(\hash.CA1.p4[11] ),
    .Q(\hash.CA2.p4[11] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[12]$_DFF_P_  (.D(\hash.CA1.p4[12] ),
    .Q(\hash.CA2.p4[12] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[13]$_DFF_P_  (.D(\hash.CA1.p4[13] ),
    .Q(\hash.CA2.p4[13] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[14]$_DFF_P_  (.D(\hash.CA1.p4[14] ),
    .Q(\hash.CA2.p4[14] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[15]$_DFF_P_  (.D(\hash.CA1.p4[15] ),
    .Q(\hash.CA2.p4[15] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[16]$_DFF_P_  (.D(\hash.CA1.p4[16] ),
    .Q(\hash.CA2.p4[16] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[17]$_DFF_P_  (.D(\hash.CA1.p4[17] ),
    .Q(\hash.CA2.p4[17] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[18]$_DFF_P_  (.D(\hash.CA1.p4[18] ),
    .Q(\hash.CA2.p4[18] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[19]$_DFF_P_  (.D(\hash.CA1.p4[19] ),
    .Q(\hash.CA2.p4[19] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[1]$_DFF_P_  (.D(\hash.CA1.p4[1] ),
    .Q(\hash.CA2.p4[1] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[20]$_DFF_P_  (.D(\hash.CA1.p4[20] ),
    .Q(\hash.CA2.p4[20] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[21]$_DFF_P_  (.D(\hash.CA1.p4[21] ),
    .Q(\hash.CA2.p4[21] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[22]$_DFF_P_  (.D(\hash.CA1.p4[22] ),
    .Q(\hash.CA2.p4[22] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[23]$_DFF_P_  (.D(\hash.CA1.p4[23] ),
    .Q(\hash.CA2.p4[23] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[24]$_DFF_P_  (.D(\hash.CA1.p4[24] ),
    .Q(\hash.CA2.p4[24] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[25]$_DFF_P_  (.D(\hash.CA1.p4[25] ),
    .Q(\hash.CA2.p4[25] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[26]$_DFF_P_  (.D(\hash.CA1.p4[26] ),
    .Q(\hash.CA2.p4[26] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[27]$_DFF_P_  (.D(\hash.CA1.p4[27] ),
    .Q(\hash.CA2.p4[27] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[28]$_DFF_P_  (.D(\hash.CA1.p4[28] ),
    .Q(\hash.CA2.p4[28] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[29]$_DFF_P_  (.D(\hash.CA1.p4[29] ),
    .Q(\hash.CA2.p4[29] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[2]$_DFF_P_  (.D(\hash.CA1.p4[2] ),
    .Q(\hash.CA2.p4[2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[30]$_DFF_P_  (.D(\hash.CA1.p4[30] ),
    .Q(\hash.CA2.p4[30] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[31]$_DFF_P_  (.D(\hash.CA1.p4[31] ),
    .Q(\hash.CA2.p4[31] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[3]$_DFF_P_  (.D(\hash.CA1.p4[3] ),
    .Q(\hash.CA2.p4[3] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[4]$_DFF_P_  (.D(\hash.CA1.p4[4] ),
    .Q(\hash.CA2.p4[4] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[5]$_DFF_P_  (.D(\hash.CA1.p4[5] ),
    .Q(\hash.CA2.p4[5] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[6]$_DFF_P_  (.D(\hash.CA1.p4[6] ),
    .Q(\hash.CA2.p4[6] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[7]$_DFF_P_  (.D(\hash.CA1.p4[7] ),
    .Q(\hash.CA2.p4[7] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[8]$_DFF_P_  (.D(\hash.CA1.p4[8] ),
    .Q(\hash.CA2.p4[8] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[9]$_DFF_P_  (.D(\hash.CA1.p4[9] ),
    .Q(\hash.CA2.p4[9] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[0]$_DFF_P_  (.D(\hash.CA1.p5[0] ),
    .Q(\hash.CA2.p5[0] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[10]$_DFF_P_  (.D(\hash.CA1.p5[10] ),
    .Q(\hash.CA2.p5[10] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[11]$_DFF_P_  (.D(\hash.CA1.p5[11] ),
    .Q(\hash.CA2.p5[11] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[12]$_DFF_P_  (.D(\hash.CA1.p5[12] ),
    .Q(\hash.CA2.p5[12] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[13]$_DFF_P_  (.D(\hash.CA1.p5[13] ),
    .Q(\hash.CA2.p5[13] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[14]$_DFF_P_  (.D(\hash.CA1.p5[14] ),
    .Q(\hash.CA2.p5[14] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[15]$_DFF_P_  (.D(\hash.CA1.p5[15] ),
    .Q(\hash.CA2.p5[15] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[16]$_DFF_P_  (.D(\hash.CA1.p5[16] ),
    .Q(\hash.CA2.p5[16] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[17]$_DFF_P_  (.D(\hash.CA1.p5[17] ),
    .Q(\hash.CA2.p5[17] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[18]$_DFF_P_  (.D(\hash.CA1.p5[18] ),
    .Q(\hash.CA2.p5[18] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[19]$_DFF_P_  (.D(\hash.CA1.p5[19] ),
    .Q(\hash.CA2.p5[19] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[1]$_DFF_P_  (.D(\hash.CA1.p5[1] ),
    .Q(\hash.CA2.p5[1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[20]$_DFF_P_  (.D(\hash.CA1.p5[20] ),
    .Q(\hash.CA2.p5[20] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[21]$_DFF_P_  (.D(\hash.CA1.p5[21] ),
    .Q(\hash.CA2.p5[21] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[22]$_DFF_P_  (.D(\hash.CA1.p5[22] ),
    .Q(\hash.CA2.p5[22] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[23]$_DFF_P_  (.D(\hash.CA1.p5[23] ),
    .Q(\hash.CA2.p5[23] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[24]$_DFF_P_  (.D(\hash.CA1.p5[24] ),
    .Q(\hash.CA2.p5[24] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[25]$_DFF_P_  (.D(\hash.CA1.p5[25] ),
    .Q(\hash.CA2.p5[25] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[26]$_DFF_P_  (.D(\hash.CA1.p5[26] ),
    .Q(\hash.CA2.p5[26] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[27]$_DFF_P_  (.D(\hash.CA1.p5[27] ),
    .Q(\hash.CA2.p5[27] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[28]$_DFF_P_  (.D(\hash.CA1.p5[28] ),
    .Q(\hash.CA2.p5[28] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[29]$_DFF_P_  (.D(\hash.CA1.p5[29] ),
    .Q(\hash.CA2.p5[29] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[2]$_DFF_P_  (.D(\hash.CA1.p5[2] ),
    .Q(\hash.CA2.p5[2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[30]$_DFF_P_  (.D(\hash.CA1.p5[30] ),
    .Q(\hash.CA2.p5[30] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[31]$_DFF_P_  (.D(\hash.CA1.p5[31] ),
    .Q(\hash.CA2.p5[31] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[3]$_DFF_P_  (.D(\hash.CA1.p5[3] ),
    .Q(\hash.CA2.p5[3] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[4]$_DFF_P_  (.D(\hash.CA1.p5[4] ),
    .Q(\hash.CA2.p5[4] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[5]$_DFF_P_  (.D(\hash.CA1.p5[5] ),
    .Q(\hash.CA2.p5[5] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[6]$_DFF_P_  (.D(\hash.CA1.p5[6] ),
    .Q(\hash.CA2.p5[6] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[7]$_DFF_P_  (.D(\hash.CA1.p5[7] ),
    .Q(\hash.CA2.p5[7] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[8]$_DFF_P_  (.D(\hash.CA1.p5[8] ),
    .Q(\hash.CA2.p5[8] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[9]$_DFF_P_  (.D(\hash.CA1.p5[9] ),
    .Q(\hash.CA2.p5[9] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[0]$_SDFF_PP0_  (.D(_00969_),
    .Q(\hash.CA1.k_i1[0] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[10]$_SDFF_PP1_  (.D(_00970_),
    .Q(\hash.CA1.k_i1[10] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[11]$_SDFF_PP1_  (.D(_00971_),
    .Q(\hash.CA1.k_i1[11] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[12]$_SDFF_PP0_  (.D(_00972_),
    .Q(\hash.CA1.k_i1[12] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[13]$_SDFF_PP1_  (.D(_00973_),
    .Q(\hash.CA1.k_i1[13] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[14]$_SDFF_PP0_  (.D(_00974_),
    .Q(\hash.CA1.k_i1[14] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[15]$_SDFF_PP0_  (.D(_00975_),
    .Q(\hash.CA1.k_i1[15] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[16]$_SDFF_PP0_  (.D(_00976_),
    .Q(\hash.CA1.k_i1[16] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[17]$_SDFF_PP1_  (.D(_00977_),
    .Q(\hash.CA1.k_i1[17] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[18]$_SDFF_PP0_  (.D(_00978_),
    .Q(\hash.CA1.k_i1[18] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[19]$_SDFF_PP1_  (.D(_00979_),
    .Q(\hash.CA1.k_i1[19] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[1]$_SDFF_PP0_  (.D(_00980_),
    .Q(\hash.CA1.k_i1[1] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[20]$_SDFF_PP0_  (.D(_00981_),
    .Q(\hash.CA1.k_i1[20] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[21]$_SDFF_PP0_  (.D(_00982_),
    .Q(\hash.CA1.k_i1[21] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[22]$_SDFF_PP0_  (.D(_00983_),
    .Q(\hash.CA1.k_i1[22] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[23]$_SDFF_PP1_  (.D(_00984_),
    .Q(\hash.CA1.k_i1[23] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[24]$_SDFF_PP0_  (.D(_00985_),
    .Q(\hash.CA1.k_i1[24] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[25]$_SDFF_PP1_  (.D(_00986_),
    .Q(\hash.CA1.k_i1[25] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[26]$_SDFF_PP0_  (.D(_00987_),
    .Q(\hash.CA1.k_i1[26] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[27]$_SDFF_PP0_  (.D(_00988_),
    .Q(\hash.CA1.k_i1[27] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[28]$_SDFF_PP0_  (.D(_00989_),
    .Q(\hash.CA1.k_i1[28] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[29]$_SDFF_PP0_  (.D(_00990_),
    .Q(\hash.CA1.k_i1[29] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[2]$_SDFF_PP0_  (.D(_00991_),
    .Q(\hash.CA1.k_i1[2] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[30]$_SDFF_PP1_  (.D(_00992_),
    .Q(\hash.CA1.k_i1[30] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[31]$_SDFF_PP0_  (.D(_00993_),
    .Q(\hash.CA1.k_i1[31] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[3]$_SDFF_PP1_  (.D(_00994_),
    .Q(\hash.CA1.k_i1[3] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[4]$_SDFF_PP1_  (.D(_00995_),
    .Q(\hash.CA1.k_i1[4] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[5]$_SDFF_PP0_  (.D(_00996_),
    .Q(\hash.CA1.k_i1[5] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[6]$_SDFF_PP0_  (.D(_00997_),
    .Q(\hash.CA1.k_i1[6] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[7]$_SDFF_PP1_  (.D(_00998_),
    .Q(\hash.CA1.k_i1[7] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[8]$_SDFF_PP1_  (.D(_00999_),
    .Q(\hash.CA1.k_i1[8] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[9]$_SDFF_PP1_  (.D(_01000_),
    .Q(\hash.CA1.k_i1[9] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[0]$_SDFF_PP1_  (.D(_01001_),
    .Q(\hash.CA1.k_i2[0] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[10]$_SDFF_PP1_  (.D(_01002_),
    .Q(\hash.CA1.k_i2[10] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[11]$_SDFF_PP0_  (.D(_01003_),
    .Q(\hash.CA1.k_i2[11] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[12]$_SDFF_PP0_  (.D(_01004_),
    .Q(\hash.CA1.k_i2[12] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[13]$_SDFF_PP0_  (.D(_01005_),
    .Q(\hash.CA1.k_i2[13] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[14]$_SDFF_PP1_  (.D(_01006_),
    .Q(\hash.CA1.k_i2[14] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[15]$_SDFF_PP0_  (.D(_01007_),
    .Q(\hash.CA1.k_i2[15] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[16]$_SDFF_PP1_  (.D(_01008_),
    .Q(\hash.CA1.k_i2[16] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[17]$_SDFF_PP1_  (.D(_01009_),
    .Q(\hash.CA1.k_i2[17] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[18]$_SDFF_PP1_  (.D(_01010_),
    .Q(\hash.CA1.k_i2[18] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[19]$_SDFF_PP0_  (.D(_01011_),
    .Q(\hash.CA1.k_i2[19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[1]$_SDFF_PP0_  (.D(_01012_),
    .Q(\hash.CA1.k_i2[1] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[20]$_SDFF_PP1_  (.D(_01013_),
    .Q(\hash.CA1.k_i2[20] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[21]$_SDFF_PP1_  (.D(_01014_),
    .Q(\hash.CA1.k_i2[21] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[22]$_SDFF_PP0_  (.D(_01015_),
    .Q(\hash.CA1.k_i2[22] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[23]$_SDFF_PP0_  (.D(_01016_),
    .Q(\hash.CA1.k_i2[23] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[24]$_SDFF_PP1_  (.D(_01017_),
    .Q(\hash.CA1.k_i2[24] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[25]$_SDFF_PP0_  (.D(_01018_),
    .Q(\hash.CA1.k_i2[25] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[26]$_SDFF_PP0_  (.D(_01019_),
    .Q(\hash.CA1.k_i2[26] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[27]$_SDFF_PP0_  (.D(_01020_),
    .Q(\hash.CA1.k_i2[27] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[28]$_SDFF_PP1_  (.D(_01021_),
    .Q(\hash.CA1.k_i2[28] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[29]$_SDFF_PP1_  (.D(_01022_),
    .Q(\hash.CA1.k_i2[29] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[2]$_SDFF_PP0_  (.D(_01023_),
    .Q(\hash.CA1.k_i2[2] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[30]$_SDFF_PP1_  (.D(_01024_),
    .Q(\hash.CA1.k_i2[30] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[31]$_SDFF_PP0_  (.D(_01025_),
    .Q(\hash.CA1.k_i2[31] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[3]$_SDFF_PP0_  (.D(_01026_),
    .Q(\hash.CA1.k_i2[3] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[4]$_SDFF_PP1_  (.D(_01027_),
    .Q(\hash.CA1.k_i2[4] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[5]$_SDFF_PP0_  (.D(_01028_),
    .Q(\hash.CA1.k_i2[5] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[6]$_SDFF_PP0_  (.D(_01029_),
    .Q(\hash.CA1.k_i2[6] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[7]$_SDFF_PP1_  (.D(_01030_),
    .Q(\hash.CA1.k_i2[7] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[8]$_SDFF_PP0_  (.D(_01031_),
    .Q(\hash.CA1.k_i2[8] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[9]$_SDFF_PP0_  (.D(_01032_),
    .Q(\hash.CA1.k_i2[9] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \ready$_DFF_P_  (.D(ready_dash),
    .Q(net1041),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \ready_dash$_SDFF_PP0_  (.D(_01033_),
    .Q(ready_dash),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \reset_hash$_DFF_P_  (.D(net1044),
    .Q(reset_hash),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \reset_hash_dash$_DFF_P_  (.D(net540),
    .Q(\hash.reset ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][0]$_DFFE_PP_  (.D(_00129_),
    .DE(_00127_),
    .Q(\w[0][0] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][10]$_DFFE_PP_  (.D(_00130_),
    .DE(_00127_),
    .Q(\w[0][10] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][11]$_DFFE_PP_  (.D(_00131_),
    .DE(_00127_),
    .Q(\w[0][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][12]$_DFFE_PP_  (.D(_00132_),
    .DE(_00127_),
    .Q(\w[0][12] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][13]$_DFFE_PP_  (.D(_00133_),
    .DE(_00127_),
    .Q(\w[0][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][14]$_DFFE_PP_  (.D(_00134_),
    .DE(_00127_),
    .Q(\w[0][14] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][15]$_DFFE_PP_  (.D(_00135_),
    .DE(_00127_),
    .Q(\w[0][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][16]$_DFFE_PP_  (.D(_00136_),
    .DE(_00127_),
    .Q(\w[0][16] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][17]$_DFFE_PP_  (.D(_00137_),
    .DE(_00127_),
    .Q(\w[0][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][18]$_DFFE_PP_  (.D(_00138_),
    .DE(_00127_),
    .Q(\w[0][18] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][19]$_DFFE_PP_  (.D(_00139_),
    .DE(_00127_),
    .Q(\w[0][19] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][1]$_DFFE_PP_  (.D(_00140_),
    .DE(_00127_),
    .Q(\w[0][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][20]$_DFFE_PP_  (.D(_00141_),
    .DE(_00127_),
    .Q(\w[0][20] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][21]$_DFFE_PP_  (.D(_00142_),
    .DE(_00127_),
    .Q(\w[0][21] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][22]$_DFFE_PP_  (.D(_00143_),
    .DE(_00127_),
    .Q(\w[0][22] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][23]$_DFFE_PP_  (.D(_00144_),
    .DE(_00127_),
    .Q(\w[0][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][24]$_DFFE_PP_  (.D(_00145_),
    .DE(_00127_),
    .Q(\w[0][24] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][25]$_DFFE_PP_  (.D(_00146_),
    .DE(_00127_),
    .Q(\w[0][25] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][26]$_DFFE_PP_  (.D(_00147_),
    .DE(_00127_),
    .Q(\w[0][26] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][27]$_DFFE_PP_  (.D(_00148_),
    .DE(_00127_),
    .Q(\w[0][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][28]$_DFFE_PP_  (.D(_00149_),
    .DE(_00127_),
    .Q(\w[0][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][29]$_DFFE_PP_  (.D(_00150_),
    .DE(_00127_),
    .Q(\w[0][29] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][2]$_DFFE_PP_  (.D(_00151_),
    .DE(_00127_),
    .Q(\w[0][2] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][30]$_DFFE_PP_  (.D(_00152_),
    .DE(_00127_),
    .Q(\w[0][30] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][31]$_DFFE_PP_  (.D(_00153_),
    .DE(_00127_),
    .Q(\w[0][31] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][3]$_DFFE_PP_  (.D(_00154_),
    .DE(_00127_),
    .Q(\w[0][3] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][4]$_DFFE_PP_  (.D(_00155_),
    .DE(_00127_),
    .Q(\w[0][4] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][5]$_DFFE_PP_  (.D(_00156_),
    .DE(_00127_),
    .Q(\w[0][5] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][6]$_DFFE_PP_  (.D(_00157_),
    .DE(_00127_),
    .Q(\w[0][6] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][7]$_DFFE_PP_  (.D(_00158_),
    .DE(_00127_),
    .Q(\w[0][7] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][8]$_DFFE_PP_  (.D(_00159_),
    .DE(_00127_),
    .Q(\w[0][8] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][9]$_DFFE_PP_  (.D(_00160_),
    .DE(_00127_),
    .Q(\w[0][9] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][0]$_DFFE_PP_  (.D(_00161_),
    .DE(_00126_),
    .Q(\w[10][0] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][10]$_DFFE_PP_  (.D(_00162_),
    .DE(_00126_),
    .Q(\w[10][10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][11]$_DFFE_PP_  (.D(_00163_),
    .DE(_00126_),
    .Q(\w[10][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][12]$_DFFE_PP_  (.D(_00164_),
    .DE(_00126_),
    .Q(\w[10][12] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][13]$_DFFE_PP_  (.D(_00165_),
    .DE(_00126_),
    .Q(\w[10][13] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][14]$_DFFE_PP_  (.D(_00166_),
    .DE(_00126_),
    .Q(\w[10][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][15]$_DFFE_PP_  (.D(_00167_),
    .DE(_00126_),
    .Q(\w[10][15] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][16]$_DFFE_PP_  (.D(_00168_),
    .DE(_00126_),
    .Q(\w[10][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][17]$_DFFE_PP_  (.D(_00169_),
    .DE(_00126_),
    .Q(\w[10][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][18]$_DFFE_PP_  (.D(_00170_),
    .DE(_00126_),
    .Q(\w[10][18] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][19]$_DFFE_PP_  (.D(_00171_),
    .DE(_00126_),
    .Q(\w[10][19] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][1]$_DFFE_PP_  (.D(_00172_),
    .DE(_00126_),
    .Q(\w[10][1] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][20]$_DFFE_PP_  (.D(_00173_),
    .DE(_00126_),
    .Q(\w[10][20] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][21]$_DFFE_PP_  (.D(_00174_),
    .DE(_00126_),
    .Q(\w[10][21] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][22]$_DFFE_PP_  (.D(_00175_),
    .DE(_00126_),
    .Q(\w[10][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][23]$_DFFE_PP_  (.D(_00176_),
    .DE(_00126_),
    .Q(\w[10][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][24]$_DFFE_PP_  (.D(_00177_),
    .DE(_00126_),
    .Q(\w[10][24] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][25]$_DFFE_PP_  (.D(_00178_),
    .DE(_00126_),
    .Q(\w[10][25] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][26]$_DFFE_PP_  (.D(_00179_),
    .DE(_00126_),
    .Q(\w[10][26] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][27]$_DFFE_PP_  (.D(_00180_),
    .DE(_00126_),
    .Q(\w[10][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][28]$_DFFE_PP_  (.D(_00181_),
    .DE(_00126_),
    .Q(\w[10][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][29]$_DFFE_PP_  (.D(_00182_),
    .DE(_00126_),
    .Q(\w[10][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][2]$_DFFE_PP_  (.D(_00183_),
    .DE(_00126_),
    .Q(\w[10][2] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][30]$_DFFE_PP_  (.D(_00184_),
    .DE(_00126_),
    .Q(\w[10][30] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][31]$_DFFE_PP_  (.D(_00185_),
    .DE(_00126_),
    .Q(\w[10][31] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][3]$_DFFE_PP_  (.D(_00186_),
    .DE(_00126_),
    .Q(\w[10][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][4]$_DFFE_PP_  (.D(_00187_),
    .DE(_00126_),
    .Q(\w[10][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][5]$_DFFE_PP_  (.D(_00188_),
    .DE(_00126_),
    .Q(\w[10][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][6]$_DFFE_PP_  (.D(_00189_),
    .DE(_00126_),
    .Q(\w[10][6] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][7]$_DFFE_PP_  (.D(_00190_),
    .DE(_00126_),
    .Q(\w[10][7] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][8]$_DFFE_PP_  (.D(_00191_),
    .DE(_00126_),
    .Q(\w[10][8] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][9]$_DFFE_PP_  (.D(_00192_),
    .DE(_00126_),
    .Q(\w[10][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][0]$_DFFE_PP_  (.D(_00193_),
    .DE(_00095_),
    .Q(\w[11][0] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][10]$_DFFE_PP_  (.D(_00194_),
    .DE(_00095_),
    .Q(\w[11][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][11]$_DFFE_PP_  (.D(_00195_),
    .DE(_00095_),
    .Q(\w[11][11] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][12]$_DFFE_PP_  (.D(_00196_),
    .DE(_00095_),
    .Q(\w[11][12] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][13]$_DFFE_PP_  (.D(_00197_),
    .DE(_00095_),
    .Q(\w[11][13] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][14]$_DFFE_PP_  (.D(_00198_),
    .DE(_00095_),
    .Q(\w[11][14] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][15]$_DFFE_PP_  (.D(_00199_),
    .DE(_00095_),
    .Q(\w[11][15] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][16]$_DFFE_PP_  (.D(_00200_),
    .DE(_00095_),
    .Q(\w[11][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][17]$_DFFE_PP_  (.D(_00201_),
    .DE(_00095_),
    .Q(\w[11][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][18]$_DFFE_PP_  (.D(_00202_),
    .DE(_00095_),
    .Q(\w[11][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][19]$_DFFE_PP_  (.D(_00203_),
    .DE(_00095_),
    .Q(\w[11][19] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][1]$_DFFE_PP_  (.D(_00204_),
    .DE(_00095_),
    .Q(\w[11][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][20]$_DFFE_PP_  (.D(_00205_),
    .DE(_00095_),
    .Q(\w[11][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][21]$_DFFE_PP_  (.D(_00206_),
    .DE(_00095_),
    .Q(\w[11][21] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][22]$_DFFE_PP_  (.D(_00207_),
    .DE(_00095_),
    .Q(\w[11][22] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][23]$_DFFE_PP_  (.D(_00208_),
    .DE(_00095_),
    .Q(\w[11][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][24]$_DFFE_PP_  (.D(_00209_),
    .DE(_00095_),
    .Q(\w[11][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][25]$_DFFE_PP_  (.D(_00210_),
    .DE(_00095_),
    .Q(\w[11][25] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][26]$_DFFE_PP_  (.D(_00211_),
    .DE(_00095_),
    .Q(\w[11][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][27]$_DFFE_PP_  (.D(_00212_),
    .DE(_00095_),
    .Q(\w[11][27] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][28]$_DFFE_PP_  (.D(_00213_),
    .DE(_00095_),
    .Q(\w[11][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][29]$_DFFE_PP_  (.D(_00214_),
    .DE(_00095_),
    .Q(\w[11][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][2]$_DFFE_PP_  (.D(_00215_),
    .DE(_00095_),
    .Q(\w[11][2] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][30]$_DFFE_PP_  (.D(_00216_),
    .DE(_00095_),
    .Q(\w[11][30] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][31]$_DFFE_PP_  (.D(_00217_),
    .DE(_00095_),
    .Q(\w[11][31] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][3]$_DFFE_PP_  (.D(_00218_),
    .DE(_00095_),
    .Q(\w[11][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][4]$_DFFE_PP_  (.D(_00219_),
    .DE(_00095_),
    .Q(\w[11][4] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][5]$_DFFE_PP_  (.D(_00220_),
    .DE(_00095_),
    .Q(\w[11][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][6]$_DFFE_PP_  (.D(_00221_),
    .DE(_00095_),
    .Q(\w[11][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][7]$_DFFE_PP_  (.D(_00222_),
    .DE(_00095_),
    .Q(\w[11][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][8]$_DFFE_PP_  (.D(_00223_),
    .DE(_00095_),
    .Q(\w[11][8] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][9]$_DFFE_PP_  (.D(_00224_),
    .DE(_00095_),
    .Q(\w[11][9] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][0]$_DFFE_PP_  (.D(_00225_),
    .DE(_00125_),
    .Q(\w[12][0] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][10]$_DFFE_PP_  (.D(_00226_),
    .DE(_00125_),
    .Q(\w[12][10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][11]$_DFFE_PP_  (.D(_00227_),
    .DE(_00125_),
    .Q(\w[12][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][12]$_DFFE_PP_  (.D(_00228_),
    .DE(_00125_),
    .Q(\w[12][12] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][13]$_DFFE_PP_  (.D(_00229_),
    .DE(_00125_),
    .Q(\w[12][13] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][14]$_DFFE_PP_  (.D(_00230_),
    .DE(_00125_),
    .Q(\w[12][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][15]$_DFFE_PP_  (.D(_00231_),
    .DE(_00125_),
    .Q(\w[12][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][16]$_DFFE_PP_  (.D(_00232_),
    .DE(_00125_),
    .Q(\w[12][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][17]$_DFFE_PP_  (.D(_00233_),
    .DE(_00125_),
    .Q(\w[12][17] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][18]$_DFFE_PP_  (.D(_00234_),
    .DE(_00125_),
    .Q(\w[12][18] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][19]$_DFFE_PP_  (.D(_00235_),
    .DE(_00125_),
    .Q(\w[12][19] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][1]$_DFFE_PP_  (.D(_00236_),
    .DE(_00125_),
    .Q(\w[12][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][20]$_DFFE_PP_  (.D(_00237_),
    .DE(_00125_),
    .Q(\w[12][20] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][21]$_DFFE_PP_  (.D(_00238_),
    .DE(_00125_),
    .Q(\w[12][21] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][22]$_DFFE_PP_  (.D(_00239_),
    .DE(_00125_),
    .Q(\w[12][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][23]$_DFFE_PP_  (.D(_00240_),
    .DE(_00125_),
    .Q(\w[12][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][24]$_DFFE_PP_  (.D(_00241_),
    .DE(_00125_),
    .Q(\w[12][24] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][25]$_DFFE_PP_  (.D(_00242_),
    .DE(_00125_),
    .Q(\w[12][25] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][26]$_DFFE_PP_  (.D(_00243_),
    .DE(_00125_),
    .Q(\w[12][26] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][27]$_DFFE_PP_  (.D(_00244_),
    .DE(_00125_),
    .Q(\w[12][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][28]$_DFFE_PP_  (.D(_00245_),
    .DE(_00125_),
    .Q(\w[12][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][29]$_DFFE_PP_  (.D(_00246_),
    .DE(_00125_),
    .Q(\w[12][29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][2]$_DFFE_PP_  (.D(_00247_),
    .DE(_00125_),
    .Q(\w[12][2] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][30]$_DFFE_PP_  (.D(_00248_),
    .DE(_00125_),
    .Q(\w[12][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][31]$_DFFE_PP_  (.D(_00249_),
    .DE(_00125_),
    .Q(\w[12][31] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][3]$_DFFE_PP_  (.D(_00250_),
    .DE(_00125_),
    .Q(\w[12][3] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][4]$_DFFE_PP_  (.D(_00251_),
    .DE(_00125_),
    .Q(\w[12][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][5]$_DFFE_PP_  (.D(_00252_),
    .DE(_00125_),
    .Q(\w[12][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][6]$_DFFE_PP_  (.D(_00253_),
    .DE(_00125_),
    .Q(\w[12][6] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][7]$_DFFE_PP_  (.D(_00254_),
    .DE(_00125_),
    .Q(\w[12][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][8]$_DFFE_PP_  (.D(_00255_),
    .DE(_00125_),
    .Q(\w[12][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][9]$_DFFE_PP_  (.D(_00256_),
    .DE(_00125_),
    .Q(\w[12][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][0]$_DFFE_PP_  (.D(_00257_),
    .DE(_00094_),
    .Q(\w[13][0] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][10]$_DFFE_PP_  (.D(_00258_),
    .DE(_00094_),
    .Q(\w[13][10] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][11]$_DFFE_PP_  (.D(_00259_),
    .DE(_00094_),
    .Q(\w[13][11] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][12]$_DFFE_PP_  (.D(_00260_),
    .DE(_00094_),
    .Q(\w[13][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][13]$_DFFE_PP_  (.D(_00261_),
    .DE(_00094_),
    .Q(\w[13][13] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][14]$_DFFE_PP_  (.D(_00262_),
    .DE(_00094_),
    .Q(\w[13][14] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][15]$_DFFE_PP_  (.D(_00263_),
    .DE(_00094_),
    .Q(\w[13][15] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][16]$_DFFE_PP_  (.D(_00264_),
    .DE(_00094_),
    .Q(\w[13][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][17]$_DFFE_PP_  (.D(_00265_),
    .DE(_00094_),
    .Q(\w[13][17] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][18]$_DFFE_PP_  (.D(_00266_),
    .DE(_00094_),
    .Q(\w[13][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][19]$_DFFE_PP_  (.D(_00267_),
    .DE(_00094_),
    .Q(\w[13][19] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][1]$_DFFE_PP_  (.D(_00268_),
    .DE(_00094_),
    .Q(\w[13][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][20]$_DFFE_PP_  (.D(_00269_),
    .DE(_00094_),
    .Q(\w[13][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][21]$_DFFE_PP_  (.D(_00270_),
    .DE(_00094_),
    .Q(\w[13][21] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][22]$_DFFE_PP_  (.D(_00271_),
    .DE(_00094_),
    .Q(\w[13][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][23]$_DFFE_PP_  (.D(_00272_),
    .DE(_00094_),
    .Q(\w[13][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][24]$_DFFE_PP_  (.D(_00273_),
    .DE(_00094_),
    .Q(\w[13][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][25]$_DFFE_PP_  (.D(_00274_),
    .DE(_00094_),
    .Q(\w[13][25] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][26]$_DFFE_PP_  (.D(_00275_),
    .DE(_00094_),
    .Q(\w[13][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][27]$_DFFE_PP_  (.D(_00276_),
    .DE(_00094_),
    .Q(\w[13][27] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][28]$_DFFE_PP_  (.D(_00277_),
    .DE(_00094_),
    .Q(\w[13][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][29]$_DFFE_PP_  (.D(_00278_),
    .DE(_00094_),
    .Q(\w[13][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][2]$_DFFE_PP_  (.D(_00279_),
    .DE(_00094_),
    .Q(\w[13][2] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][30]$_DFFE_PP_  (.D(_00280_),
    .DE(_00094_),
    .Q(\w[13][30] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][31]$_DFFE_PP_  (.D(_00281_),
    .DE(_00094_),
    .Q(\w[13][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][3]$_DFFE_PP_  (.D(_00282_),
    .DE(_00094_),
    .Q(\w[13][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][4]$_DFFE_PP_  (.D(_00283_),
    .DE(_00094_),
    .Q(\w[13][4] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][5]$_DFFE_PP_  (.D(_00284_),
    .DE(_00094_),
    .Q(\w[13][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][6]$_DFFE_PP_  (.D(_00285_),
    .DE(_00094_),
    .Q(\w[13][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][7]$_DFFE_PP_  (.D(_00286_),
    .DE(_00094_),
    .Q(\w[13][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][8]$_DFFE_PP_  (.D(_00287_),
    .DE(_00094_),
    .Q(\w[13][8] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][9]$_DFFE_PP_  (.D(_00288_),
    .DE(_00094_),
    .Q(\w[13][9] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][0]$_DFFE_PP_  (.D(_00289_),
    .DE(_00124_),
    .Q(\w[14][0] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][10]$_DFFE_PP_  (.D(_00290_),
    .DE(_00124_),
    .Q(\w[14][10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][11]$_DFFE_PP_  (.D(_00291_),
    .DE(_00124_),
    .Q(\w[14][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][12]$_DFFE_PP_  (.D(_00292_),
    .DE(_00124_),
    .Q(\w[14][12] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][13]$_DFFE_PP_  (.D(_00293_),
    .DE(_00124_),
    .Q(\w[14][13] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][14]$_DFFE_PP_  (.D(_00294_),
    .DE(_00124_),
    .Q(\w[14][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][15]$_DFFE_PP_  (.D(_00295_),
    .DE(_00124_),
    .Q(\w[14][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][16]$_DFFE_PP_  (.D(_00296_),
    .DE(_00124_),
    .Q(\w[14][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][17]$_DFFE_PP_  (.D(_00297_),
    .DE(_00124_),
    .Q(\w[14][17] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][18]$_DFFE_PP_  (.D(_00298_),
    .DE(_00124_),
    .Q(\w[14][18] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][19]$_DFFE_PP_  (.D(_00299_),
    .DE(_00124_),
    .Q(\w[14][19] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][1]$_DFFE_PP_  (.D(_00300_),
    .DE(_00124_),
    .Q(\w[14][1] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][20]$_DFFE_PP_  (.D(_00301_),
    .DE(_00124_),
    .Q(\w[14][20] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][21]$_DFFE_PP_  (.D(_00302_),
    .DE(_00124_),
    .Q(\w[14][21] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][22]$_DFFE_PP_  (.D(_00303_),
    .DE(_00124_),
    .Q(\w[14][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][23]$_DFFE_PP_  (.D(_00304_),
    .DE(_00124_),
    .Q(\w[14][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][24]$_DFFE_PP_  (.D(_00305_),
    .DE(_00124_),
    .Q(\w[14][24] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][25]$_DFFE_PP_  (.D(_00306_),
    .DE(_00124_),
    .Q(\w[14][25] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][26]$_DFFE_PP_  (.D(_00307_),
    .DE(_00124_),
    .Q(\w[14][26] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][27]$_DFFE_PP_  (.D(_00308_),
    .DE(_00124_),
    .Q(\w[14][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][28]$_DFFE_PP_  (.D(_00309_),
    .DE(_00124_),
    .Q(\w[14][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][29]$_DFFE_PP_  (.D(_00310_),
    .DE(_00124_),
    .Q(\w[14][29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][2]$_DFFE_PP_  (.D(_00311_),
    .DE(_00124_),
    .Q(\w[14][2] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][30]$_DFFE_PP_  (.D(_00312_),
    .DE(_00124_),
    .Q(\w[14][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][31]$_DFFE_PP_  (.D(_00313_),
    .DE(_00124_),
    .Q(\w[14][31] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][3]$_DFFE_PP_  (.D(_00314_),
    .DE(_00124_),
    .Q(\w[14][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][4]$_DFFE_PP_  (.D(_00315_),
    .DE(_00124_),
    .Q(\w[14][4] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][5]$_DFFE_PP_  (.D(_00316_),
    .DE(_00124_),
    .Q(\w[14][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][6]$_DFFE_PP_  (.D(_00317_),
    .DE(_00124_),
    .Q(\w[14][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][7]$_DFFE_PP_  (.D(_00318_),
    .DE(_00124_),
    .Q(\w[14][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][8]$_DFFE_PP_  (.D(_00319_),
    .DE(_00124_),
    .Q(\w[14][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][9]$_DFFE_PP_  (.D(_00320_),
    .DE(_00124_),
    .Q(\w[14][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][0]$_DFFE_PP_  (.D(_00321_),
    .DE(_00093_),
    .Q(\w[15][0] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][10]$_DFFE_PP_  (.D(_00322_),
    .DE(_00093_),
    .Q(\w[15][10] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][11]$_DFFE_PP_  (.D(_00323_),
    .DE(_00093_),
    .Q(\w[15][11] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][12]$_DFFE_PP_  (.D(_00324_),
    .DE(_00093_),
    .Q(\w[15][12] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][13]$_DFFE_PP_  (.D(_00325_),
    .DE(_00093_),
    .Q(\w[15][13] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][14]$_DFFE_PP_  (.D(_00326_),
    .DE(_00093_),
    .Q(\w[15][14] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][15]$_DFFE_PP_  (.D(_00327_),
    .DE(_00093_),
    .Q(\w[15][15] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][16]$_DFFE_PP_  (.D(_00328_),
    .DE(_00093_),
    .Q(\w[15][16] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][17]$_DFFE_PP_  (.D(_00329_),
    .DE(_00093_),
    .Q(\w[15][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][18]$_DFFE_PP_  (.D(_00330_),
    .DE(_00093_),
    .Q(\w[15][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][19]$_DFFE_PP_  (.D(_00331_),
    .DE(_00093_),
    .Q(\w[15][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][1]$_DFFE_PP_  (.D(_00332_),
    .DE(_00093_),
    .Q(\w[15][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][20]$_DFFE_PP_  (.D(_00333_),
    .DE(_00093_),
    .Q(\w[15][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][21]$_DFFE_PP_  (.D(_00334_),
    .DE(_00093_),
    .Q(\w[15][21] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][22]$_DFFE_PP_  (.D(_00335_),
    .DE(_00093_),
    .Q(\w[15][22] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][23]$_DFFE_PP_  (.D(_00336_),
    .DE(_00093_),
    .Q(\w[15][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][24]$_DFFE_PP_  (.D(_00337_),
    .DE(_00093_),
    .Q(\w[15][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][25]$_DFFE_PP_  (.D(_00338_),
    .DE(_00093_),
    .Q(\w[15][25] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][26]$_DFFE_PP_  (.D(_00339_),
    .DE(_00093_),
    .Q(\w[15][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][27]$_DFFE_PP_  (.D(_00340_),
    .DE(_00093_),
    .Q(\w[15][27] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][28]$_DFFE_PP_  (.D(_00341_),
    .DE(_00093_),
    .Q(\w[15][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][29]$_DFFE_PP_  (.D(_00342_),
    .DE(_00093_),
    .Q(\w[15][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][2]$_DFFE_PP_  (.D(_00343_),
    .DE(_00093_),
    .Q(\w[15][2] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][30]$_DFFE_PP_  (.D(_00344_),
    .DE(_00093_),
    .Q(\w[15][30] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][31]$_DFFE_PP_  (.D(_00345_),
    .DE(_00093_),
    .Q(\w[15][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][3]$_DFFE_PP_  (.D(_00346_),
    .DE(_00093_),
    .Q(\w[15][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][4]$_DFFE_PP_  (.D(_00347_),
    .DE(_00093_),
    .Q(\w[15][4] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][5]$_DFFE_PP_  (.D(_00348_),
    .DE(_00093_),
    .Q(\w[15][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][6]$_DFFE_PP_  (.D(_00349_),
    .DE(_00093_),
    .Q(\w[15][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][7]$_DFFE_PP_  (.D(_00350_),
    .DE(_00093_),
    .Q(\w[15][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][8]$_DFFE_PP_  (.D(_00351_),
    .DE(_00093_),
    .Q(\w[15][8] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][9]$_DFFE_PP_  (.D(_00352_),
    .DE(_00093_),
    .Q(\w[15][9] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][0]$_SDFFCE_PN0P_  (.D(_01034_),
    .DE(_00123_),
    .Q(\w[16][0] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][10]$_SDFFCE_PN0P_  (.D(_01035_),
    .DE(_00123_),
    .Q(\w[16][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][11]$_SDFFCE_PN0P_  (.D(_01036_),
    .DE(_00123_),
    .Q(\w[16][11] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][12]$_SDFFCE_PN0P_  (.D(_01037_),
    .DE(_00123_),
    .Q(\w[16][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][13]$_SDFFCE_PN0P_  (.D(_01038_),
    .DE(_00123_),
    .Q(\w[16][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][14]$_SDFFCE_PN0P_  (.D(_01039_),
    .DE(_00123_),
    .Q(\w[16][14] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][15]$_SDFFCE_PN0P_  (.D(_01040_),
    .DE(_00123_),
    .Q(\w[16][15] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][16]$_SDFFCE_PN0P_  (.D(_01041_),
    .DE(_00123_),
    .Q(\w[16][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][17]$_SDFFCE_PN0P_  (.D(_01042_),
    .DE(_00123_),
    .Q(\w[16][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][18]$_SDFFCE_PN0P_  (.D(_01043_),
    .DE(_00123_),
    .Q(\w[16][18] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][19]$_SDFFCE_PN0P_  (.D(_01044_),
    .DE(_00123_),
    .Q(\w[16][19] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][1]$_SDFFCE_PN0P_  (.D(_01045_),
    .DE(_00123_),
    .Q(\w[16][1] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][20]$_SDFFCE_PN0P_  (.D(_01046_),
    .DE(_00123_),
    .Q(\w[16][20] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][21]$_SDFFCE_PN0P_  (.D(_01047_),
    .DE(_00123_),
    .Q(\w[16][21] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][22]$_SDFFCE_PN0P_  (.D(_01048_),
    .DE(_00123_),
    .Q(\w[16][22] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][23]$_SDFFCE_PN0P_  (.D(_01049_),
    .DE(_00123_),
    .Q(\w[16][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][24]$_SDFFCE_PN0P_  (.D(_01050_),
    .DE(_00123_),
    .Q(\w[16][24] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][25]$_SDFFCE_PN0P_  (.D(_01051_),
    .DE(_00123_),
    .Q(\w[16][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][26]$_SDFFCE_PN0P_  (.D(_01052_),
    .DE(_00123_),
    .Q(\w[16][26] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][27]$_SDFFCE_PN0P_  (.D(_01053_),
    .DE(_00123_),
    .Q(\w[16][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][28]$_SDFFCE_PN0P_  (.D(_01054_),
    .DE(_00123_),
    .Q(\w[16][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][29]$_SDFFCE_PN0P_  (.D(_01055_),
    .DE(_00123_),
    .Q(\w[16][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][2]$_SDFFCE_PN0P_  (.D(_01056_),
    .DE(_00123_),
    .Q(\w[16][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][30]$_SDFFCE_PN0P_  (.D(_01057_),
    .DE(_00123_),
    .Q(\w[16][30] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][31]$_SDFFCE_PN0P_  (.D(_01058_),
    .DE(_00123_),
    .Q(\w[16][31] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][3]$_SDFFCE_PN0P_  (.D(_01059_),
    .DE(_00123_),
    .Q(\w[16][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][4]$_SDFFCE_PN0P_  (.D(_01060_),
    .DE(_00123_),
    .Q(\w[16][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][5]$_SDFFCE_PN0P_  (.D(_01061_),
    .DE(_00123_),
    .Q(\w[16][5] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][6]$_SDFFCE_PN0P_  (.D(_01062_),
    .DE(_00123_),
    .Q(\w[16][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][7]$_SDFFCE_PN0P_  (.D(_01063_),
    .DE(_00123_),
    .Q(\w[16][7] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][8]$_SDFFCE_PN0P_  (.D(_01064_),
    .DE(_00123_),
    .Q(\w[16][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][9]$_SDFFCE_PN0P_  (.D(_01065_),
    .DE(_00123_),
    .Q(\w[16][9] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][0]$_SDFFCE_PN0P_  (.D(_01066_),
    .DE(_00092_),
    .Q(\w[17][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][10]$_SDFFCE_PN0P_  (.D(_01067_),
    .DE(_00092_),
    .Q(\w[17][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][11]$_SDFFCE_PN0P_  (.D(_01068_),
    .DE(_00092_),
    .Q(\w[17][11] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][12]$_SDFFCE_PN0P_  (.D(_01069_),
    .DE(_00092_),
    .Q(\w[17][12] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][13]$_SDFFCE_PN0P_  (.D(_01070_),
    .DE(_00092_),
    .Q(\w[17][13] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][14]$_SDFFCE_PN0P_  (.D(_01071_),
    .DE(_00092_),
    .Q(\w[17][14] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][15]$_SDFFCE_PN0P_  (.D(_01072_),
    .DE(_00092_),
    .Q(\w[17][15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][16]$_SDFFCE_PN0P_  (.D(_01073_),
    .DE(_00092_),
    .Q(\w[17][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][17]$_SDFFCE_PN0P_  (.D(_01074_),
    .DE(_00092_),
    .Q(\w[17][17] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][18]$_SDFFCE_PN0P_  (.D(_01075_),
    .DE(_00092_),
    .Q(\w[17][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][19]$_SDFFCE_PN0P_  (.D(_01076_),
    .DE(_00092_),
    .Q(\w[17][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][1]$_SDFFCE_PN0P_  (.D(_01077_),
    .DE(_00092_),
    .Q(\w[17][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][20]$_SDFFCE_PN0P_  (.D(_01078_),
    .DE(_00092_),
    .Q(\w[17][20] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][21]$_SDFFCE_PN0P_  (.D(_01079_),
    .DE(_00092_),
    .Q(\w[17][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][22]$_SDFFCE_PN0P_  (.D(_01080_),
    .DE(_00092_),
    .Q(\w[17][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][23]$_SDFFCE_PN0P_  (.D(_01081_),
    .DE(_00092_),
    .Q(\w[17][23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][24]$_SDFFCE_PN0P_  (.D(_01082_),
    .DE(_00092_),
    .Q(\w[17][24] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][25]$_SDFFCE_PN0P_  (.D(_01083_),
    .DE(_00092_),
    .Q(\w[17][25] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][26]$_SDFFCE_PN0P_  (.D(_01084_),
    .DE(_00092_),
    .Q(\w[17][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][27]$_SDFFCE_PN0P_  (.D(_01085_),
    .DE(_00092_),
    .Q(\w[17][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][28]$_SDFFCE_PN0P_  (.D(_01086_),
    .DE(_00092_),
    .Q(\w[17][28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][29]$_SDFFCE_PN0P_  (.D(_01087_),
    .DE(_00092_),
    .Q(\w[17][29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][2]$_SDFFCE_PN0P_  (.D(_01088_),
    .DE(_00092_),
    .Q(\w[17][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][30]$_SDFFCE_PN0P_  (.D(_01089_),
    .DE(_00092_),
    .Q(\w[17][30] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][31]$_SDFFCE_PN0P_  (.D(_01090_),
    .DE(_00092_),
    .Q(\w[17][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][3]$_SDFFCE_PN0P_  (.D(_01091_),
    .DE(_00092_),
    .Q(\w[17][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][4]$_SDFFCE_PN0P_  (.D(_01092_),
    .DE(_00092_),
    .Q(\w[17][4] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][5]$_SDFFCE_PN0P_  (.D(_01093_),
    .DE(_00092_),
    .Q(\w[17][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][6]$_SDFFCE_PN0P_  (.D(_01094_),
    .DE(_00092_),
    .Q(\w[17][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][7]$_SDFFCE_PN0P_  (.D(_01095_),
    .DE(_00092_),
    .Q(\w[17][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][8]$_SDFFCE_PN0P_  (.D(_01096_),
    .DE(_00092_),
    .Q(\w[17][8] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][9]$_SDFFCE_PN0P_  (.D(_01097_),
    .DE(_00092_),
    .Q(\w[17][9] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][0]$_SDFFCE_PN0P_  (.D(_01098_),
    .DE(_00122_),
    .Q(\w[18][0] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][10]$_SDFFCE_PN0P_  (.D(_01099_),
    .DE(_00122_),
    .Q(\w[18][10] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][11]$_SDFFCE_PN0P_  (.D(_01100_),
    .DE(_00122_),
    .Q(\w[18][11] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][12]$_SDFFCE_PN0P_  (.D(_01101_),
    .DE(_00122_),
    .Q(\w[18][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][13]$_SDFFCE_PN0P_  (.D(_01102_),
    .DE(_00122_),
    .Q(\w[18][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][14]$_SDFFCE_PN0P_  (.D(_01103_),
    .DE(_00122_),
    .Q(\w[18][14] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][15]$_SDFFCE_PN0P_  (.D(_01104_),
    .DE(_00122_),
    .Q(\w[18][15] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][16]$_SDFFCE_PN0P_  (.D(_01105_),
    .DE(_00122_),
    .Q(\w[18][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][17]$_SDFFCE_PN0P_  (.D(_01106_),
    .DE(_00122_),
    .Q(\w[18][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][18]$_SDFFCE_PN0P_  (.D(_01107_),
    .DE(_00122_),
    .Q(\w[18][18] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][19]$_SDFFCE_PN0P_  (.D(_01108_),
    .DE(_00122_),
    .Q(\w[18][19] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][1]$_SDFFCE_PN0P_  (.D(_01109_),
    .DE(_00122_),
    .Q(\w[18][1] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][20]$_SDFFCE_PN0P_  (.D(_01110_),
    .DE(_00122_),
    .Q(\w[18][20] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][21]$_SDFFCE_PN0P_  (.D(_01111_),
    .DE(_00122_),
    .Q(\w[18][21] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][22]$_SDFFCE_PN0P_  (.D(_01112_),
    .DE(_00122_),
    .Q(\w[18][22] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][23]$_SDFFCE_PN0P_  (.D(_01113_),
    .DE(_00122_),
    .Q(\w[18][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][24]$_SDFFCE_PN0P_  (.D(_01114_),
    .DE(_00122_),
    .Q(\w[18][24] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][25]$_SDFFCE_PN0P_  (.D(_01115_),
    .DE(_00122_),
    .Q(\w[18][25] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][26]$_SDFFCE_PN0P_  (.D(_01116_),
    .DE(_00122_),
    .Q(\w[18][26] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][27]$_SDFFCE_PN0P_  (.D(_01117_),
    .DE(_00122_),
    .Q(\w[18][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][28]$_SDFFCE_PN0P_  (.D(_01118_),
    .DE(_00122_),
    .Q(\w[18][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][29]$_SDFFCE_PN0P_  (.D(_01119_),
    .DE(_00122_),
    .Q(\w[18][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][2]$_SDFFCE_PN0P_  (.D(_01120_),
    .DE(_00122_),
    .Q(\w[18][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][30]$_SDFFCE_PN0P_  (.D(_01121_),
    .DE(_00122_),
    .Q(\w[18][30] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][31]$_SDFFCE_PN0P_  (.D(_01122_),
    .DE(_00122_),
    .Q(\w[18][31] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][3]$_SDFFCE_PN0P_  (.D(_01123_),
    .DE(_00122_),
    .Q(\w[18][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][4]$_SDFFCE_PN0P_  (.D(_01124_),
    .DE(_00122_),
    .Q(\w[18][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][5]$_SDFFCE_PN0P_  (.D(_01125_),
    .DE(_00122_),
    .Q(\w[18][5] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][6]$_SDFFCE_PN0P_  (.D(_01126_),
    .DE(_00122_),
    .Q(\w[18][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][7]$_SDFFCE_PN0P_  (.D(_01127_),
    .DE(_00122_),
    .Q(\w[18][7] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][8]$_SDFFCE_PN0P_  (.D(_01128_),
    .DE(_00122_),
    .Q(\w[18][8] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][9]$_SDFFCE_PN0P_  (.D(_01129_),
    .DE(_00122_),
    .Q(\w[18][9] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][0]$_SDFFCE_PN0P_  (.D(_01130_),
    .DE(_00091_),
    .Q(\w[19][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][10]$_SDFFCE_PN0P_  (.D(_01131_),
    .DE(_00091_),
    .Q(\w[19][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][11]$_SDFFCE_PN0P_  (.D(_01132_),
    .DE(_00091_),
    .Q(\w[19][11] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][12]$_SDFFCE_PN0P_  (.D(_01133_),
    .DE(_00091_),
    .Q(\w[19][12] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][13]$_SDFFCE_PN0P_  (.D(_01134_),
    .DE(_00091_),
    .Q(\w[19][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][14]$_SDFFCE_PN0P_  (.D(_01135_),
    .DE(_00091_),
    .Q(\w[19][14] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][15]$_SDFFCE_PN0P_  (.D(_01136_),
    .DE(_00091_),
    .Q(\w[19][15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][16]$_SDFFCE_PN0P_  (.D(_01137_),
    .DE(_00091_),
    .Q(\w[19][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][17]$_SDFFCE_PN0P_  (.D(_01138_),
    .DE(_00091_),
    .Q(\w[19][17] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][18]$_SDFFCE_PN0P_  (.D(_01139_),
    .DE(_00091_),
    .Q(\w[19][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][19]$_SDFFCE_PN0P_  (.D(_01140_),
    .DE(_00091_),
    .Q(\w[19][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][1]$_SDFFCE_PN0P_  (.D(_01141_),
    .DE(_00091_),
    .Q(\w[19][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][20]$_SDFFCE_PN0P_  (.D(_01142_),
    .DE(_00091_),
    .Q(\w[19][20] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][21]$_SDFFCE_PN0P_  (.D(_01143_),
    .DE(_00091_),
    .Q(\w[19][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][22]$_SDFFCE_PN0P_  (.D(_01144_),
    .DE(_00091_),
    .Q(\w[19][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][23]$_SDFFCE_PN0P_  (.D(_01145_),
    .DE(_00091_),
    .Q(\w[19][23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][24]$_SDFFCE_PN0P_  (.D(_01146_),
    .DE(_00091_),
    .Q(\w[19][24] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][25]$_SDFFCE_PN0P_  (.D(_01147_),
    .DE(_00091_),
    .Q(\w[19][25] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][26]$_SDFFCE_PN0P_  (.D(_01148_),
    .DE(_00091_),
    .Q(\w[19][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][27]$_SDFFCE_PN0P_  (.D(_01149_),
    .DE(_00091_),
    .Q(\w[19][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][28]$_SDFFCE_PN0P_  (.D(_01150_),
    .DE(_00091_),
    .Q(\w[19][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][29]$_SDFFCE_PN0P_  (.D(_01151_),
    .DE(_00091_),
    .Q(\w[19][29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][2]$_SDFFCE_PN0P_  (.D(_01152_),
    .DE(_00091_),
    .Q(\w[19][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][30]$_SDFFCE_PN0P_  (.D(_01153_),
    .DE(_00091_),
    .Q(\w[19][30] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][31]$_SDFFCE_PN0P_  (.D(_01154_),
    .DE(_00091_),
    .Q(\w[19][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][3]$_SDFFCE_PN0P_  (.D(_01155_),
    .DE(_00091_),
    .Q(\w[19][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][4]$_SDFFCE_PN0P_  (.D(_01156_),
    .DE(_00091_),
    .Q(\w[19][4] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][5]$_SDFFCE_PN0P_  (.D(_01157_),
    .DE(_00091_),
    .Q(\w[19][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][6]$_SDFFCE_PN0P_  (.D(_01158_),
    .DE(_00091_),
    .Q(\w[19][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][7]$_SDFFCE_PN0P_  (.D(_01159_),
    .DE(_00091_),
    .Q(\w[19][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][8]$_SDFFCE_PN0P_  (.D(_01160_),
    .DE(_00091_),
    .Q(\w[19][8] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][9]$_SDFFCE_PN0P_  (.D(_01161_),
    .DE(_00091_),
    .Q(\w[19][9] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][0]$_DFFE_PP_  (.D(_00353_),
    .DE(_00090_),
    .Q(\w[1][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][10]$_DFFE_PP_  (.D(_00354_),
    .DE(_00090_),
    .Q(\w[1][10] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][11]$_DFFE_PP_  (.D(_00355_),
    .DE(_00090_),
    .Q(\w[1][11] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][12]$_DFFE_PP_  (.D(_00356_),
    .DE(_00090_),
    .Q(\w[1][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][13]$_DFFE_PP_  (.D(_00357_),
    .DE(_00090_),
    .Q(\w[1][13] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][14]$_DFFE_PP_  (.D(_00358_),
    .DE(_00090_),
    .Q(\w[1][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][15]$_DFFE_PP_  (.D(_00359_),
    .DE(_00090_),
    .Q(\w[1][15] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][16]$_DFFE_PP_  (.D(_00360_),
    .DE(_00090_),
    .Q(\w[1][16] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][17]$_DFFE_PP_  (.D(_00361_),
    .DE(_00090_),
    .Q(\w[1][17] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][18]$_DFFE_PP_  (.D(_00362_),
    .DE(_00090_),
    .Q(\w[1][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][19]$_DFFE_PP_  (.D(_00363_),
    .DE(_00090_),
    .Q(\w[1][19] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][1]$_DFFE_PP_  (.D(_00364_),
    .DE(_00090_),
    .Q(\w[1][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][20]$_DFFE_PP_  (.D(_00365_),
    .DE(_00090_),
    .Q(\w[1][20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][21]$_DFFE_PP_  (.D(_00366_),
    .DE(_00090_),
    .Q(\w[1][21] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][22]$_DFFE_PP_  (.D(_00367_),
    .DE(_00090_),
    .Q(\w[1][22] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][23]$_DFFE_PP_  (.D(_00368_),
    .DE(_00090_),
    .Q(\w[1][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][24]$_DFFE_PP_  (.D(_00369_),
    .DE(_00090_),
    .Q(\w[1][24] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][25]$_DFFE_PP_  (.D(_00370_),
    .DE(_00090_),
    .Q(\w[1][25] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][26]$_DFFE_PP_  (.D(_00371_),
    .DE(_00090_),
    .Q(\w[1][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][27]$_DFFE_PP_  (.D(_00372_),
    .DE(_00090_),
    .Q(\w[1][27] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][28]$_DFFE_PP_  (.D(_00373_),
    .DE(_00090_),
    .Q(\w[1][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][29]$_DFFE_PP_  (.D(_00374_),
    .DE(_00090_),
    .Q(\w[1][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][2]$_DFFE_PP_  (.D(_00375_),
    .DE(_00090_),
    .Q(\w[1][2] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][30]$_DFFE_PP_  (.D(_00376_),
    .DE(_00090_),
    .Q(\w[1][30] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][31]$_DFFE_PP_  (.D(_00377_),
    .DE(_00090_),
    .Q(\w[1][31] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][3]$_DFFE_PP_  (.D(_00378_),
    .DE(_00090_),
    .Q(\w[1][3] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][4]$_DFFE_PP_  (.D(_00379_),
    .DE(_00090_),
    .Q(\w[1][4] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][5]$_DFFE_PP_  (.D(_00380_),
    .DE(_00090_),
    .Q(\w[1][5] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][6]$_DFFE_PP_  (.D(_00381_),
    .DE(_00090_),
    .Q(\w[1][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][7]$_DFFE_PP_  (.D(_00382_),
    .DE(_00090_),
    .Q(\w[1][7] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][8]$_DFFE_PP_  (.D(_00383_),
    .DE(_00090_),
    .Q(\w[1][8] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][9]$_DFFE_PP_  (.D(_00384_),
    .DE(_00090_),
    .Q(\w[1][9] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][0]$_SDFFCE_PN0P_  (.D(_01162_),
    .DE(_00121_),
    .Q(\w[20][0] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][10]$_SDFFCE_PN0P_  (.D(_01163_),
    .DE(_00121_),
    .Q(\w[20][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][11]$_SDFFCE_PN0P_  (.D(_01164_),
    .DE(_00121_),
    .Q(\w[20][11] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][12]$_SDFFCE_PN0P_  (.D(_01165_),
    .DE(_00121_),
    .Q(\w[20][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][13]$_SDFFCE_PN0P_  (.D(_01166_),
    .DE(_00121_),
    .Q(\w[20][13] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][14]$_SDFFCE_PN0P_  (.D(_01167_),
    .DE(_00121_),
    .Q(\w[20][14] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][15]$_SDFFCE_PN0P_  (.D(_01168_),
    .DE(_00121_),
    .Q(\w[20][15] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][16]$_SDFFCE_PN0P_  (.D(_01169_),
    .DE(_00121_),
    .Q(\w[20][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][17]$_SDFFCE_PN0P_  (.D(_01170_),
    .DE(_00121_),
    .Q(\w[20][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][18]$_SDFFCE_PN0P_  (.D(_01171_),
    .DE(_00121_),
    .Q(\w[20][18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][19]$_SDFFCE_PN0P_  (.D(_01172_),
    .DE(_00121_),
    .Q(\w[20][19] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][1]$_SDFFCE_PN0P_  (.D(_01173_),
    .DE(_00121_),
    .Q(\w[20][1] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][20]$_SDFFCE_PN0P_  (.D(_01174_),
    .DE(_00121_),
    .Q(\w[20][20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][21]$_SDFFCE_PN0P_  (.D(_01175_),
    .DE(_00121_),
    .Q(\w[20][21] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][22]$_SDFFCE_PN0P_  (.D(_01176_),
    .DE(_00121_),
    .Q(\w[20][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][23]$_SDFFCE_PN0P_  (.D(_01177_),
    .DE(_00121_),
    .Q(\w[20][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][24]$_SDFFCE_PN0P_  (.D(_01178_),
    .DE(_00121_),
    .Q(\w[20][24] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][25]$_SDFFCE_PN0P_  (.D(_01179_),
    .DE(_00121_),
    .Q(\w[20][25] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][26]$_SDFFCE_PN0P_  (.D(_01180_),
    .DE(_00121_),
    .Q(\w[20][26] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][27]$_SDFFCE_PN0P_  (.D(_01181_),
    .DE(_00121_),
    .Q(\w[20][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][28]$_SDFFCE_PN0P_  (.D(_01182_),
    .DE(_00121_),
    .Q(\w[20][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][29]$_SDFFCE_PN0P_  (.D(_01183_),
    .DE(_00121_),
    .Q(\w[20][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][2]$_SDFFCE_PN0P_  (.D(_01184_),
    .DE(_00121_),
    .Q(\w[20][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][30]$_SDFFCE_PN0P_  (.D(_01185_),
    .DE(_00121_),
    .Q(\w[20][30] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][31]$_SDFFCE_PN0P_  (.D(_01186_),
    .DE(_00121_),
    .Q(\w[20][31] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][3]$_SDFFCE_PN0P_  (.D(_01187_),
    .DE(_00121_),
    .Q(\w[20][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][4]$_SDFFCE_PN0P_  (.D(_01188_),
    .DE(_00121_),
    .Q(\w[20][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][5]$_SDFFCE_PN0P_  (.D(_01189_),
    .DE(_00121_),
    .Q(\w[20][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][6]$_SDFFCE_PN0P_  (.D(_01190_),
    .DE(_00121_),
    .Q(\w[20][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][7]$_SDFFCE_PN0P_  (.D(_01191_),
    .DE(_00121_),
    .Q(\w[20][7] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][8]$_SDFFCE_PN0P_  (.D(_01192_),
    .DE(_00121_),
    .Q(\w[20][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][9]$_SDFFCE_PN0P_  (.D(_01193_),
    .DE(_00121_),
    .Q(\w[20][9] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][0]$_SDFFCE_PN0P_  (.D(_01194_),
    .DE(_00089_),
    .Q(\w[21][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][10]$_SDFFCE_PN0P_  (.D(_01195_),
    .DE(_00089_),
    .Q(\w[21][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][11]$_SDFFCE_PN0P_  (.D(_01196_),
    .DE(_00089_),
    .Q(\w[21][11] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][12]$_SDFFCE_PN0P_  (.D(_01197_),
    .DE(_00089_),
    .Q(\w[21][12] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][13]$_SDFFCE_PN0P_  (.D(_01198_),
    .DE(_00089_),
    .Q(\w[21][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][14]$_SDFFCE_PN0P_  (.D(_01199_),
    .DE(_00089_),
    .Q(\w[21][14] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][15]$_SDFFCE_PN0P_  (.D(_01200_),
    .DE(_00089_),
    .Q(\w[21][15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][16]$_SDFFCE_PN0P_  (.D(_01201_),
    .DE(_00089_),
    .Q(\w[21][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][17]$_SDFFCE_PN0P_  (.D(_01202_),
    .DE(_00089_),
    .Q(\w[21][17] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][18]$_SDFFCE_PN0P_  (.D(_01203_),
    .DE(_00089_),
    .Q(\w[21][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][19]$_SDFFCE_PN0P_  (.D(_01204_),
    .DE(_00089_),
    .Q(\w[21][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][1]$_SDFFCE_PN0P_  (.D(_01205_),
    .DE(_00089_),
    .Q(\w[21][1] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][20]$_SDFFCE_PN0P_  (.D(_01206_),
    .DE(_00089_),
    .Q(\w[21][20] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][21]$_SDFFCE_PN0P_  (.D(_01207_),
    .DE(_00089_),
    .Q(\w[21][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][22]$_SDFFCE_PN0P_  (.D(_01208_),
    .DE(_00089_),
    .Q(\w[21][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][23]$_SDFFCE_PN0P_  (.D(_01209_),
    .DE(_00089_),
    .Q(\w[21][23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][24]$_SDFFCE_PN0P_  (.D(_01210_),
    .DE(_00089_),
    .Q(\w[21][24] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][25]$_SDFFCE_PN0P_  (.D(_01211_),
    .DE(_00089_),
    .Q(\w[21][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][26]$_SDFFCE_PN0P_  (.D(_01212_),
    .DE(_00089_),
    .Q(\w[21][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][27]$_SDFFCE_PN0P_  (.D(_01213_),
    .DE(_00089_),
    .Q(\w[21][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][28]$_SDFFCE_PN0P_  (.D(_01214_),
    .DE(_00089_),
    .Q(\w[21][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][29]$_SDFFCE_PN0P_  (.D(_01215_),
    .DE(_00089_),
    .Q(\w[21][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][2]$_SDFFCE_PN0P_  (.D(_01216_),
    .DE(_00089_),
    .Q(\w[21][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][30]$_SDFFCE_PN0P_  (.D(_01217_),
    .DE(_00089_),
    .Q(\w[21][30] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][31]$_SDFFCE_PN0P_  (.D(_01218_),
    .DE(_00089_),
    .Q(\w[21][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][3]$_SDFFCE_PN0P_  (.D(_01219_),
    .DE(_00089_),
    .Q(\w[21][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][4]$_SDFFCE_PN0P_  (.D(_01220_),
    .DE(_00089_),
    .Q(\w[21][4] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][5]$_SDFFCE_PN0P_  (.D(_01221_),
    .DE(_00089_),
    .Q(\w[21][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][6]$_SDFFCE_PN0P_  (.D(_01222_),
    .DE(_00089_),
    .Q(\w[21][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][7]$_SDFFCE_PN0P_  (.D(_01223_),
    .DE(_00089_),
    .Q(\w[21][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][8]$_SDFFCE_PN0P_  (.D(_01224_),
    .DE(_00089_),
    .Q(\w[21][8] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][9]$_SDFFCE_PN0P_  (.D(_01225_),
    .DE(_00089_),
    .Q(\w[21][9] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][0]$_SDFFCE_PN0P_  (.D(_01226_),
    .DE(_00120_),
    .Q(\w[22][0] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][10]$_SDFFCE_PN0P_  (.D(_01227_),
    .DE(_00120_),
    .Q(\w[22][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][11]$_SDFFCE_PN0P_  (.D(_01228_),
    .DE(_00120_),
    .Q(\w[22][11] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][12]$_SDFFCE_PN0P_  (.D(_01229_),
    .DE(_00120_),
    .Q(\w[22][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][13]$_SDFFCE_PN0P_  (.D(_01230_),
    .DE(_00120_),
    .Q(\w[22][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][14]$_SDFFCE_PN0P_  (.D(_01231_),
    .DE(_00120_),
    .Q(\w[22][14] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][15]$_SDFFCE_PN0P_  (.D(_01232_),
    .DE(_00120_),
    .Q(\w[22][15] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][16]$_SDFFCE_PN0P_  (.D(_01233_),
    .DE(_00120_),
    .Q(\w[22][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][17]$_SDFFCE_PN0P_  (.D(_01234_),
    .DE(_00120_),
    .Q(\w[22][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][18]$_SDFFCE_PN0P_  (.D(_01235_),
    .DE(_00120_),
    .Q(\w[22][18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][19]$_SDFFCE_PN0P_  (.D(_01236_),
    .DE(_00120_),
    .Q(\w[22][19] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][1]$_SDFFCE_PN0P_  (.D(_01237_),
    .DE(_00120_),
    .Q(\w[22][1] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][20]$_SDFFCE_PN0P_  (.D(_01238_),
    .DE(_00120_),
    .Q(\w[22][20] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][21]$_SDFFCE_PN0P_  (.D(_01239_),
    .DE(_00120_),
    .Q(\w[22][21] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][22]$_SDFFCE_PN0P_  (.D(_01240_),
    .DE(_00120_),
    .Q(\w[22][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][23]$_SDFFCE_PN0P_  (.D(_01241_),
    .DE(_00120_),
    .Q(\w[22][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][24]$_SDFFCE_PN0P_  (.D(_01242_),
    .DE(_00120_),
    .Q(\w[22][24] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][25]$_SDFFCE_PN0P_  (.D(_01243_),
    .DE(_00120_),
    .Q(\w[22][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][26]$_SDFFCE_PN0P_  (.D(_01244_),
    .DE(_00120_),
    .Q(\w[22][26] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][27]$_SDFFCE_PN0P_  (.D(_01245_),
    .DE(_00120_),
    .Q(\w[22][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][28]$_SDFFCE_PN0P_  (.D(_01246_),
    .DE(_00120_),
    .Q(\w[22][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][29]$_SDFFCE_PN0P_  (.D(_01247_),
    .DE(_00120_),
    .Q(\w[22][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][2]$_SDFFCE_PN0P_  (.D(_01248_),
    .DE(_00120_),
    .Q(\w[22][2] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][30]$_SDFFCE_PN0P_  (.D(_01249_),
    .DE(_00120_),
    .Q(\w[22][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][31]$_SDFFCE_PN0P_  (.D(_01250_),
    .DE(_00120_),
    .Q(\w[22][31] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][3]$_SDFFCE_PN0P_  (.D(_01251_),
    .DE(_00120_),
    .Q(\w[22][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][4]$_SDFFCE_PN0P_  (.D(_01252_),
    .DE(_00120_),
    .Q(\w[22][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][5]$_SDFFCE_PN0P_  (.D(_01253_),
    .DE(_00120_),
    .Q(\w[22][5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][6]$_SDFFCE_PN0P_  (.D(_01254_),
    .DE(_00120_),
    .Q(\w[22][6] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][7]$_SDFFCE_PN0P_  (.D(_01255_),
    .DE(_00120_),
    .Q(\w[22][7] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][8]$_SDFFCE_PN0P_  (.D(_01256_),
    .DE(_00120_),
    .Q(\w[22][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][9]$_SDFFCE_PN0P_  (.D(_01257_),
    .DE(_00120_),
    .Q(\w[22][9] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][0]$_SDFFCE_PN0P_  (.D(_01258_),
    .DE(net306),
    .Q(\w[23][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][10]$_SDFFCE_PN0P_  (.D(_01259_),
    .DE(net307),
    .Q(\w[23][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][11]$_SDFFCE_PN0P_  (.D(_01260_),
    .DE(net306),
    .Q(\w[23][11] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][12]$_SDFFCE_PN0P_  (.D(_01261_),
    .DE(net306),
    .Q(\w[23][12] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][13]$_SDFFCE_PN0P_  (.D(_01262_),
    .DE(net307),
    .Q(\w[23][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][14]$_SDFFCE_PN0P_  (.D(_01263_),
    .DE(net306),
    .Q(\w[23][14] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][15]$_SDFFCE_PN0P_  (.D(_01264_),
    .DE(_00088_),
    .Q(\w[23][15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][16]$_SDFFCE_PN0P_  (.D(_01265_),
    .DE(net306),
    .Q(\w[23][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][17]$_SDFFCE_PN0P_  (.D(_01266_),
    .DE(net306),
    .Q(\w[23][17] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][18]$_SDFFCE_PN0P_  (.D(_01267_),
    .DE(net307),
    .Q(\w[23][18] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][19]$_SDFFCE_PN0P_  (.D(_01268_),
    .DE(net306),
    .Q(\w[23][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][1]$_SDFFCE_PN0P_  (.D(_01269_),
    .DE(net306),
    .Q(\w[23][1] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][20]$_SDFFCE_PN0P_  (.D(_01270_),
    .DE(net307),
    .Q(\w[23][20] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][21]$_SDFFCE_PN0P_  (.D(_01271_),
    .DE(net307),
    .Q(\w[23][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][22]$_SDFFCE_PN0P_  (.D(_01272_),
    .DE(net306),
    .Q(\w[23][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][23]$_SDFFCE_PN0P_  (.D(_01273_),
    .DE(_00088_),
    .Q(\w[23][23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][24]$_SDFFCE_PN0P_  (.D(_01274_),
    .DE(_00088_),
    .Q(\w[23][24] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][25]$_SDFFCE_PN0P_  (.D(_01275_),
    .DE(net306),
    .Q(\w[23][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][26]$_SDFFCE_PN0P_  (.D(_01276_),
    .DE(_00088_),
    .Q(\w[23][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][27]$_SDFFCE_PN0P_  (.D(_01277_),
    .DE(net306),
    .Q(\w[23][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][28]$_SDFFCE_PN0P_  (.D(_01278_),
    .DE(_00088_),
    .Q(\w[23][28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][29]$_SDFFCE_PN0P_  (.D(_01279_),
    .DE(_00088_),
    .Q(\w[23][29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][2]$_SDFFCE_PN0P_  (.D(_01280_),
    .DE(net306),
    .Q(\w[23][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][30]$_SDFFCE_PN0P_  (.D(_01281_),
    .DE(_00088_),
    .Q(\w[23][30] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][31]$_SDFFCE_PN0P_  (.D(_01282_),
    .DE(net306),
    .Q(\w[23][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][3]$_SDFFCE_PN0P_  (.D(_01283_),
    .DE(net306),
    .Q(\w[23][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][4]$_SDFFCE_PN0P_  (.D(_01284_),
    .DE(net306),
    .Q(\w[23][4] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][5]$_SDFFCE_PN0P_  (.D(_01285_),
    .DE(net306),
    .Q(\w[23][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][6]$_SDFFCE_PN0P_  (.D(_01286_),
    .DE(_00088_),
    .Q(\w[23][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][7]$_SDFFCE_PN0P_  (.D(_01287_),
    .DE(_00088_),
    .Q(\w[23][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][8]$_SDFFCE_PN0P_  (.D(_01288_),
    .DE(net306),
    .Q(\w[23][8] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][9]$_SDFFCE_PN0P_  (.D(_01289_),
    .DE(net307),
    .Q(\w[23][9] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][0]$_SDFFCE_PN0P_  (.D(_01290_),
    .DE(_00119_),
    .Q(\w[24][0] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][10]$_SDFFCE_PN0P_  (.D(_01291_),
    .DE(_00119_),
    .Q(\w[24][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][11]$_SDFFCE_PN0P_  (.D(_01292_),
    .DE(_00119_),
    .Q(\w[24][11] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][12]$_SDFFCE_PN0P_  (.D(_01293_),
    .DE(_00119_),
    .Q(\w[24][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][13]$_SDFFCE_PN0P_  (.D(_01294_),
    .DE(_00119_),
    .Q(\w[24][13] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][14]$_SDFFCE_PN0P_  (.D(_01295_),
    .DE(_00119_),
    .Q(\w[24][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][15]$_SDFFCE_PN0P_  (.D(_01296_),
    .DE(_00119_),
    .Q(\w[24][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][16]$_SDFFCE_PN0P_  (.D(_01297_),
    .DE(_00119_),
    .Q(\w[24][16] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][17]$_SDFFCE_PN0P_  (.D(_01298_),
    .DE(_00119_),
    .Q(\w[24][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][18]$_SDFFCE_PN0P_  (.D(_01299_),
    .DE(_00119_),
    .Q(\w[24][18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][19]$_SDFFCE_PN0P_  (.D(_01300_),
    .DE(_00119_),
    .Q(\w[24][19] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][1]$_SDFFCE_PN0P_  (.D(_01301_),
    .DE(_00119_),
    .Q(\w[24][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][20]$_SDFFCE_PN0P_  (.D(_01302_),
    .DE(_00119_),
    .Q(\w[24][20] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][21]$_SDFFCE_PN0P_  (.D(_01303_),
    .DE(_00119_),
    .Q(\w[24][21] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][22]$_SDFFCE_PN0P_  (.D(_01304_),
    .DE(_00119_),
    .Q(\w[24][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][23]$_SDFFCE_PN0P_  (.D(_01305_),
    .DE(_00119_),
    .Q(\w[24][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][24]$_SDFFCE_PN0P_  (.D(_01306_),
    .DE(_00119_),
    .Q(\w[24][24] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][25]$_SDFFCE_PN0P_  (.D(_01307_),
    .DE(_00119_),
    .Q(\w[24][25] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][26]$_SDFFCE_PN0P_  (.D(_01308_),
    .DE(_00119_),
    .Q(\w[24][26] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][27]$_SDFFCE_PN0P_  (.D(_01309_),
    .DE(_00119_),
    .Q(\w[24][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][28]$_SDFFCE_PN0P_  (.D(_01310_),
    .DE(_00119_),
    .Q(\w[24][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][29]$_SDFFCE_PN0P_  (.D(_01311_),
    .DE(_00119_),
    .Q(\w[24][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][2]$_SDFFCE_PN0P_  (.D(_01312_),
    .DE(_00119_),
    .Q(\w[24][2] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][30]$_SDFFCE_PN0P_  (.D(_01313_),
    .DE(_00119_),
    .Q(\w[24][30] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][31]$_SDFFCE_PN0P_  (.D(_01314_),
    .DE(_00119_),
    .Q(\w[24][31] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][3]$_SDFFCE_PN0P_  (.D(_01315_),
    .DE(_00119_),
    .Q(\w[24][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][4]$_SDFFCE_PN0P_  (.D(_01316_),
    .DE(_00119_),
    .Q(\w[24][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][5]$_SDFFCE_PN0P_  (.D(_01317_),
    .DE(_00119_),
    .Q(\w[24][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][6]$_SDFFCE_PN0P_  (.D(_01318_),
    .DE(_00119_),
    .Q(\w[24][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][7]$_SDFFCE_PN0P_  (.D(_01319_),
    .DE(_00119_),
    .Q(\w[24][7] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][8]$_SDFFCE_PN0P_  (.D(_01320_),
    .DE(_00119_),
    .Q(\w[24][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][9]$_SDFFCE_PN0P_  (.D(_01321_),
    .DE(_00119_),
    .Q(\w[24][9] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][0]$_SDFFCE_PN0P_  (.D(_01322_),
    .DE(_00087_),
    .Q(\w[25][0] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][10]$_SDFFCE_PN0P_  (.D(_01323_),
    .DE(_00087_),
    .Q(\w[25][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][11]$_SDFFCE_PN0P_  (.D(_01324_),
    .DE(_00087_),
    .Q(\w[25][11] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][12]$_SDFFCE_PN0P_  (.D(_01325_),
    .DE(_00087_),
    .Q(\w[25][12] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][13]$_SDFFCE_PN0P_  (.D(_01326_),
    .DE(_00087_),
    .Q(\w[25][13] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][14]$_SDFFCE_PN0P_  (.D(_01327_),
    .DE(_00087_),
    .Q(\w[25][14] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][15]$_SDFFCE_PN0P_  (.D(_01328_),
    .DE(_00087_),
    .Q(\w[25][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][16]$_SDFFCE_PN0P_  (.D(_01329_),
    .DE(_00087_),
    .Q(\w[25][16] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][17]$_SDFFCE_PN0P_  (.D(_01330_),
    .DE(_00087_),
    .Q(\w[25][17] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][18]$_SDFFCE_PN0P_  (.D(_01331_),
    .DE(_00087_),
    .Q(\w[25][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][19]$_SDFFCE_PN0P_  (.D(_01332_),
    .DE(_00087_),
    .Q(\w[25][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][1]$_SDFFCE_PN0P_  (.D(_01333_),
    .DE(_00087_),
    .Q(\w[25][1] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][20]$_SDFFCE_PN0P_  (.D(_01334_),
    .DE(_00087_),
    .Q(\w[25][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][21]$_SDFFCE_PN0P_  (.D(_01335_),
    .DE(_00087_),
    .Q(\w[25][21] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][22]$_SDFFCE_PN0P_  (.D(_01336_),
    .DE(_00087_),
    .Q(\w[25][22] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][23]$_SDFFCE_PN0P_  (.D(_01337_),
    .DE(_00087_),
    .Q(\w[25][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][24]$_SDFFCE_PN0P_  (.D(_01338_),
    .DE(_00087_),
    .Q(\w[25][24] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][25]$_SDFFCE_PN0P_  (.D(_01339_),
    .DE(_00087_),
    .Q(\w[25][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][26]$_SDFFCE_PN0P_  (.D(_01340_),
    .DE(_00087_),
    .Q(\w[25][26] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][27]$_SDFFCE_PN0P_  (.D(_01341_),
    .DE(_00087_),
    .Q(\w[25][27] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][28]$_SDFFCE_PN0P_  (.D(_01342_),
    .DE(_00087_),
    .Q(\w[25][28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][29]$_SDFFCE_PN0P_  (.D(_01343_),
    .DE(_00087_),
    .Q(\w[25][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][2]$_SDFFCE_PN0P_  (.D(_01344_),
    .DE(_00087_),
    .Q(\w[25][2] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][30]$_SDFFCE_PN0P_  (.D(_01345_),
    .DE(_00087_),
    .Q(\w[25][30] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][31]$_SDFFCE_PN0P_  (.D(_01346_),
    .DE(_00087_),
    .Q(\w[25][31] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][3]$_SDFFCE_PN0P_  (.D(_01347_),
    .DE(_00087_),
    .Q(\w[25][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][4]$_SDFFCE_PN0P_  (.D(_01348_),
    .DE(_00087_),
    .Q(\w[25][4] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][5]$_SDFFCE_PN0P_  (.D(_01349_),
    .DE(_00087_),
    .Q(\w[25][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][6]$_SDFFCE_PN0P_  (.D(_01350_),
    .DE(_00087_),
    .Q(\w[25][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][7]$_SDFFCE_PN0P_  (.D(_01351_),
    .DE(_00087_),
    .Q(\w[25][7] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][8]$_SDFFCE_PN0P_  (.D(_01352_),
    .DE(_00087_),
    .Q(\w[25][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][9]$_SDFFCE_PN0P_  (.D(_01353_),
    .DE(_00087_),
    .Q(\w[25][9] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][0]$_SDFFCE_PN0P_  (.D(_01354_),
    .DE(_00118_),
    .Q(\w[26][0] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][10]$_SDFFCE_PN0P_  (.D(_01355_),
    .DE(_00118_),
    .Q(\w[26][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][11]$_SDFFCE_PN0P_  (.D(_01356_),
    .DE(_00118_),
    .Q(\w[26][11] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][12]$_SDFFCE_PN0P_  (.D(_01357_),
    .DE(_00118_),
    .Q(\w[26][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][13]$_SDFFCE_PN0P_  (.D(_01358_),
    .DE(_00118_),
    .Q(\w[26][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][14]$_SDFFCE_PN0P_  (.D(_01359_),
    .DE(_00118_),
    .Q(\w[26][14] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][15]$_SDFFCE_PN0P_  (.D(_01360_),
    .DE(_00118_),
    .Q(\w[26][15] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][16]$_SDFFCE_PN0P_  (.D(_01361_),
    .DE(_00118_),
    .Q(\w[26][16] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][17]$_SDFFCE_PN0P_  (.D(_01362_),
    .DE(_00118_),
    .Q(\w[26][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][18]$_SDFFCE_PN0P_  (.D(_01363_),
    .DE(_00118_),
    .Q(\w[26][18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][19]$_SDFFCE_PN0P_  (.D(_01364_),
    .DE(_00118_),
    .Q(\w[26][19] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][1]$_SDFFCE_PN0P_  (.D(_01365_),
    .DE(_00118_),
    .Q(\w[26][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][20]$_SDFFCE_PN0P_  (.D(_01366_),
    .DE(_00118_),
    .Q(\w[26][20] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][21]$_SDFFCE_PN0P_  (.D(_01367_),
    .DE(_00118_),
    .Q(\w[26][21] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][22]$_SDFFCE_PN0P_  (.D(_01368_),
    .DE(_00118_),
    .Q(\w[26][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][23]$_SDFFCE_PN0P_  (.D(_01369_),
    .DE(_00118_),
    .Q(\w[26][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][24]$_SDFFCE_PN0P_  (.D(_01370_),
    .DE(_00118_),
    .Q(\w[26][24] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][25]$_SDFFCE_PN0P_  (.D(_01371_),
    .DE(_00118_),
    .Q(\w[26][25] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][26]$_SDFFCE_PN0P_  (.D(_01372_),
    .DE(_00118_),
    .Q(\w[26][26] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][27]$_SDFFCE_PN0P_  (.D(_01373_),
    .DE(_00118_),
    .Q(\w[26][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][28]$_SDFFCE_PN0P_  (.D(_01374_),
    .DE(_00118_),
    .Q(\w[26][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][29]$_SDFFCE_PN0P_  (.D(_01375_),
    .DE(_00118_),
    .Q(\w[26][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][2]$_SDFFCE_PN0P_  (.D(_01376_),
    .DE(_00118_),
    .Q(\w[26][2] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][30]$_SDFFCE_PN0P_  (.D(_01377_),
    .DE(_00118_),
    .Q(\w[26][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][31]$_SDFFCE_PN0P_  (.D(_01378_),
    .DE(_00118_),
    .Q(\w[26][31] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][3]$_SDFFCE_PN0P_  (.D(_01379_),
    .DE(_00118_),
    .Q(\w[26][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][4]$_SDFFCE_PN0P_  (.D(_01380_),
    .DE(_00118_),
    .Q(\w[26][4] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][5]$_SDFFCE_PN0P_  (.D(_01381_),
    .DE(_00118_),
    .Q(\w[26][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][6]$_SDFFCE_PN0P_  (.D(_01382_),
    .DE(_00118_),
    .Q(\w[26][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][7]$_SDFFCE_PN0P_  (.D(_01383_),
    .DE(_00118_),
    .Q(\w[26][7] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][8]$_SDFFCE_PN0P_  (.D(_01384_),
    .DE(_00118_),
    .Q(\w[26][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][9]$_SDFFCE_PN0P_  (.D(_01385_),
    .DE(_00118_),
    .Q(\w[26][9] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][0]$_SDFFCE_PN0P_  (.D(_01386_),
    .DE(_00086_),
    .Q(\w[27][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][10]$_SDFFCE_PN0P_  (.D(_01387_),
    .DE(_00086_),
    .Q(\w[27][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][11]$_SDFFCE_PN0P_  (.D(_01388_),
    .DE(_00086_),
    .Q(\w[27][11] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][12]$_SDFFCE_PN0P_  (.D(_01389_),
    .DE(_00086_),
    .Q(\w[27][12] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][13]$_SDFFCE_PN0P_  (.D(_01390_),
    .DE(_00086_),
    .Q(\w[27][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][14]$_SDFFCE_PN0P_  (.D(_01391_),
    .DE(_00086_),
    .Q(\w[27][14] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][15]$_SDFFCE_PN0P_  (.D(_01392_),
    .DE(_00086_),
    .Q(\w[27][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][16]$_SDFFCE_PN0P_  (.D(_01393_),
    .DE(_00086_),
    .Q(\w[27][16] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][17]$_SDFFCE_PN0P_  (.D(_01394_),
    .DE(_00086_),
    .Q(\w[27][17] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][18]$_SDFFCE_PN0P_  (.D(_01395_),
    .DE(_00086_),
    .Q(\w[27][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][19]$_SDFFCE_PN0P_  (.D(_01396_),
    .DE(_00086_),
    .Q(\w[27][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][1]$_SDFFCE_PN0P_  (.D(_01397_),
    .DE(_00086_),
    .Q(\w[27][1] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][20]$_SDFFCE_PN0P_  (.D(_01398_),
    .DE(_00086_),
    .Q(\w[27][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][21]$_SDFFCE_PN0P_  (.D(_01399_),
    .DE(_00086_),
    .Q(\w[27][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][22]$_SDFFCE_PN0P_  (.D(_01400_),
    .DE(_00086_),
    .Q(\w[27][22] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][23]$_SDFFCE_PN0P_  (.D(_01401_),
    .DE(_00086_),
    .Q(\w[27][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][24]$_SDFFCE_PN0P_  (.D(_01402_),
    .DE(_00086_),
    .Q(\w[27][24] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][25]$_SDFFCE_PN0P_  (.D(_01403_),
    .DE(_00086_),
    .Q(\w[27][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][26]$_SDFFCE_PN0P_  (.D(_01404_),
    .DE(_00086_),
    .Q(\w[27][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][27]$_SDFFCE_PN0P_  (.D(_01405_),
    .DE(_00086_),
    .Q(\w[27][27] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][28]$_SDFFCE_PN0P_  (.D(_01406_),
    .DE(_00086_),
    .Q(\w[27][28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][29]$_SDFFCE_PN0P_  (.D(_01407_),
    .DE(_00086_),
    .Q(\w[27][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][2]$_SDFFCE_PN0P_  (.D(_01408_),
    .DE(_00086_),
    .Q(\w[27][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][30]$_SDFFCE_PN0P_  (.D(_01409_),
    .DE(_00086_),
    .Q(\w[27][30] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][31]$_SDFFCE_PN0P_  (.D(_01410_),
    .DE(_00086_),
    .Q(\w[27][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][3]$_SDFFCE_PN0P_  (.D(_01411_),
    .DE(_00086_),
    .Q(\w[27][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][4]$_SDFFCE_PN0P_  (.D(_01412_),
    .DE(_00086_),
    .Q(\w[27][4] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][5]$_SDFFCE_PN0P_  (.D(_01413_),
    .DE(_00086_),
    .Q(\w[27][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][6]$_SDFFCE_PN0P_  (.D(_01414_),
    .DE(_00086_),
    .Q(\w[27][6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][7]$_SDFFCE_PN0P_  (.D(_01415_),
    .DE(_00086_),
    .Q(\w[27][7] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][8]$_SDFFCE_PN0P_  (.D(_01416_),
    .DE(_00086_),
    .Q(\w[27][8] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][9]$_SDFFCE_PN0P_  (.D(_01417_),
    .DE(_00086_),
    .Q(\w[27][9] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][0]$_SDFFCE_PN0P_  (.D(_01418_),
    .DE(_00117_),
    .Q(\w[28][0] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][10]$_SDFFCE_PN0P_  (.D(_01419_),
    .DE(_00117_),
    .Q(\w[28][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][11]$_SDFFCE_PN0P_  (.D(_01420_),
    .DE(_00117_),
    .Q(\w[28][11] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][12]$_SDFFCE_PN0P_  (.D(_01421_),
    .DE(_00117_),
    .Q(\w[28][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][13]$_SDFFCE_PN0P_  (.D(_01422_),
    .DE(_00117_),
    .Q(\w[28][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][14]$_SDFFCE_PN0P_  (.D(_01423_),
    .DE(_00117_),
    .Q(\w[28][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][15]$_SDFFCE_PN0P_  (.D(_01424_),
    .DE(_00117_),
    .Q(\w[28][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][16]$_SDFFCE_PN0P_  (.D(_01425_),
    .DE(_00117_),
    .Q(\w[28][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][17]$_SDFFCE_PN0P_  (.D(_01426_),
    .DE(_00117_),
    .Q(\w[28][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][18]$_SDFFCE_PN0P_  (.D(_01427_),
    .DE(_00117_),
    .Q(\w[28][18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][19]$_SDFFCE_PN0P_  (.D(_01428_),
    .DE(_00117_),
    .Q(\w[28][19] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][1]$_SDFFCE_PN0P_  (.D(_01429_),
    .DE(_00117_),
    .Q(\w[28][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][20]$_SDFFCE_PN0P_  (.D(_01430_),
    .DE(_00117_),
    .Q(\w[28][20] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][21]$_SDFFCE_PN0P_  (.D(_01431_),
    .DE(_00117_),
    .Q(\w[28][21] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][22]$_SDFFCE_PN0P_  (.D(_01432_),
    .DE(_00117_),
    .Q(\w[28][22] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][23]$_SDFFCE_PN0P_  (.D(_01433_),
    .DE(_00117_),
    .Q(\w[28][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][24]$_SDFFCE_PN0P_  (.D(_01434_),
    .DE(_00117_),
    .Q(\w[28][24] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][25]$_SDFFCE_PN0P_  (.D(_01435_),
    .DE(_00117_),
    .Q(\w[28][25] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][26]$_SDFFCE_PN0P_  (.D(_01436_),
    .DE(_00117_),
    .Q(\w[28][26] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][27]$_SDFFCE_PN0P_  (.D(_01437_),
    .DE(_00117_),
    .Q(\w[28][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][28]$_SDFFCE_PN0P_  (.D(_01438_),
    .DE(_00117_),
    .Q(\w[28][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][29]$_SDFFCE_PN0P_  (.D(_01439_),
    .DE(_00117_),
    .Q(\w[28][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][2]$_SDFFCE_PN0P_  (.D(_01440_),
    .DE(_00117_),
    .Q(\w[28][2] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][30]$_SDFFCE_PN0P_  (.D(_01441_),
    .DE(_00117_),
    .Q(\w[28][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][31]$_SDFFCE_PN0P_  (.D(_01442_),
    .DE(_00117_),
    .Q(\w[28][31] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][3]$_SDFFCE_PN0P_  (.D(_01443_),
    .DE(_00117_),
    .Q(\w[28][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][4]$_SDFFCE_PN0P_  (.D(_01444_),
    .DE(_00117_),
    .Q(\w[28][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][5]$_SDFFCE_PN0P_  (.D(_01445_),
    .DE(_00117_),
    .Q(\w[28][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][6]$_SDFFCE_PN0P_  (.D(_01446_),
    .DE(_00117_),
    .Q(\w[28][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][7]$_SDFFCE_PN0P_  (.D(_01447_),
    .DE(_00117_),
    .Q(\w[28][7] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][8]$_SDFFCE_PN0P_  (.D(_01448_),
    .DE(_00117_),
    .Q(\w[28][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][9]$_SDFFCE_PN0P_  (.D(_01449_),
    .DE(_00117_),
    .Q(\w[28][9] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][0]$_SDFFCE_PN0P_  (.D(_01450_),
    .DE(_00085_),
    .Q(\w[29][0] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][10]$_SDFFCE_PN0P_  (.D(_01451_),
    .DE(_00085_),
    .Q(\w[29][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][11]$_SDFFCE_PN0P_  (.D(_01452_),
    .DE(_00085_),
    .Q(\w[29][11] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][12]$_SDFFCE_PN0P_  (.D(_01453_),
    .DE(_00085_),
    .Q(\w[29][12] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][13]$_SDFFCE_PN0P_  (.D(_01454_),
    .DE(_00085_),
    .Q(\w[29][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][14]$_SDFFCE_PN0P_  (.D(_01455_),
    .DE(_00085_),
    .Q(\w[29][14] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][15]$_SDFFCE_PN0P_  (.D(_01456_),
    .DE(_00085_),
    .Q(\w[29][15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][16]$_SDFFCE_PN0P_  (.D(_01457_),
    .DE(_00085_),
    .Q(\w[29][16] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][17]$_SDFFCE_PN0P_  (.D(_01458_),
    .DE(_00085_),
    .Q(\w[29][17] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][18]$_SDFFCE_PN0P_  (.D(_01459_),
    .DE(_00085_),
    .Q(\w[29][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][19]$_SDFFCE_PN0P_  (.D(_01460_),
    .DE(_00085_),
    .Q(\w[29][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][1]$_SDFFCE_PN0P_  (.D(_01461_),
    .DE(_00085_),
    .Q(\w[29][1] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][20]$_SDFFCE_PN0P_  (.D(_01462_),
    .DE(_00085_),
    .Q(\w[29][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][21]$_SDFFCE_PN0P_  (.D(_01463_),
    .DE(_00085_),
    .Q(\w[29][21] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][22]$_SDFFCE_PN0P_  (.D(_01464_),
    .DE(_00085_),
    .Q(\w[29][22] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][23]$_SDFFCE_PN0P_  (.D(_01465_),
    .DE(_00085_),
    .Q(\w[29][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][24]$_SDFFCE_PN0P_  (.D(_01466_),
    .DE(_00085_),
    .Q(\w[29][24] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][25]$_SDFFCE_PN0P_  (.D(_01467_),
    .DE(_00085_),
    .Q(\w[29][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][26]$_SDFFCE_PN0P_  (.D(_01468_),
    .DE(_00085_),
    .Q(\w[29][26] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][27]$_SDFFCE_PN0P_  (.D(_01469_),
    .DE(_00085_),
    .Q(\w[29][27] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][28]$_SDFFCE_PN0P_  (.D(_01470_),
    .DE(_00085_),
    .Q(\w[29][28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][29]$_SDFFCE_PN0P_  (.D(_01471_),
    .DE(_00085_),
    .Q(\w[29][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][2]$_SDFFCE_PN0P_  (.D(_01472_),
    .DE(_00085_),
    .Q(\w[29][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][30]$_SDFFCE_PN0P_  (.D(_01473_),
    .DE(_00085_),
    .Q(\w[29][30] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][31]$_SDFFCE_PN0P_  (.D(_01474_),
    .DE(_00085_),
    .Q(\w[29][31] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][3]$_SDFFCE_PN0P_  (.D(_01475_),
    .DE(_00085_),
    .Q(\w[29][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][4]$_SDFFCE_PN0P_  (.D(_01476_),
    .DE(_00085_),
    .Q(\w[29][4] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][5]$_SDFFCE_PN0P_  (.D(_01477_),
    .DE(_00085_),
    .Q(\w[29][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][6]$_SDFFCE_PN0P_  (.D(_01478_),
    .DE(_00085_),
    .Q(\w[29][6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][7]$_SDFFCE_PN0P_  (.D(_01479_),
    .DE(_00085_),
    .Q(\w[29][7] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][8]$_SDFFCE_PN0P_  (.D(_01480_),
    .DE(_00085_),
    .Q(\w[29][8] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][9]$_SDFFCE_PN0P_  (.D(_01481_),
    .DE(_00085_),
    .Q(\w[29][9] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][0]$_DFFE_PP_  (.D(_00385_),
    .DE(_00116_),
    .Q(\w[2][0] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][10]$_DFFE_PP_  (.D(_00386_),
    .DE(_00116_),
    .Q(\w[2][10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][11]$_DFFE_PP_  (.D(_00387_),
    .DE(_00116_),
    .Q(\w[2][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][12]$_DFFE_PP_  (.D(_00388_),
    .DE(_00116_),
    .Q(\w[2][12] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][13]$_DFFE_PP_  (.D(_00389_),
    .DE(_00116_),
    .Q(\w[2][13] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][14]$_DFFE_PP_  (.D(_00390_),
    .DE(_00116_),
    .Q(\w[2][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][15]$_DFFE_PP_  (.D(_00391_),
    .DE(_00116_),
    .Q(\w[2][15] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][16]$_DFFE_PP_  (.D(_00392_),
    .DE(_00116_),
    .Q(\w[2][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][17]$_DFFE_PP_  (.D(_00393_),
    .DE(_00116_),
    .Q(\w[2][17] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][18]$_DFFE_PP_  (.D(_00394_),
    .DE(_00116_),
    .Q(\w[2][18] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][19]$_DFFE_PP_  (.D(_00395_),
    .DE(_00116_),
    .Q(\w[2][19] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][1]$_DFFE_PP_  (.D(_00396_),
    .DE(_00116_),
    .Q(\w[2][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][20]$_DFFE_PP_  (.D(_00397_),
    .DE(_00116_),
    .Q(\w[2][20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][21]$_DFFE_PP_  (.D(_00398_),
    .DE(_00116_),
    .Q(\w[2][21] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][22]$_DFFE_PP_  (.D(_00399_),
    .DE(_00116_),
    .Q(\w[2][22] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][23]$_DFFE_PP_  (.D(_00400_),
    .DE(_00116_),
    .Q(\w[2][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][24]$_DFFE_PP_  (.D(_00401_),
    .DE(_00116_),
    .Q(\w[2][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][25]$_DFFE_PP_  (.D(_00402_),
    .DE(_00116_),
    .Q(\w[2][25] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][26]$_DFFE_PP_  (.D(_00403_),
    .DE(_00116_),
    .Q(\w[2][26] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][27]$_DFFE_PP_  (.D(_00404_),
    .DE(_00116_),
    .Q(\w[2][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][28]$_DFFE_PP_  (.D(_00405_),
    .DE(_00116_),
    .Q(\w[2][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][29]$_DFFE_PP_  (.D(_00406_),
    .DE(_00116_),
    .Q(\w[2][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][2]$_DFFE_PP_  (.D(_00407_),
    .DE(_00116_),
    .Q(\w[2][2] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][30]$_DFFE_PP_  (.D(_00408_),
    .DE(_00116_),
    .Q(\w[2][30] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][31]$_DFFE_PP_  (.D(_00409_),
    .DE(_00116_),
    .Q(\w[2][31] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][3]$_DFFE_PP_  (.D(_00410_),
    .DE(_00116_),
    .Q(\w[2][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][4]$_DFFE_PP_  (.D(_00411_),
    .DE(_00116_),
    .Q(\w[2][4] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][5]$_DFFE_PP_  (.D(_00412_),
    .DE(_00116_),
    .Q(\w[2][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][6]$_DFFE_PP_  (.D(_00413_),
    .DE(_00116_),
    .Q(\w[2][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][7]$_DFFE_PP_  (.D(_00414_),
    .DE(_00116_),
    .Q(\w[2][7] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][8]$_DFFE_PP_  (.D(_00415_),
    .DE(_00116_),
    .Q(\w[2][8] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][9]$_DFFE_PP_  (.D(_00416_),
    .DE(_00116_),
    .Q(\w[2][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][0]$_SDFFCE_PN0P_  (.D(_01482_),
    .DE(_00115_),
    .Q(\w[30][0] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][10]$_SDFFCE_PN0P_  (.D(_01483_),
    .DE(_00115_),
    .Q(\w[30][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][11]$_SDFFCE_PN0P_  (.D(_01484_),
    .DE(_00115_),
    .Q(\w[30][11] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][12]$_SDFFCE_PN0P_  (.D(_01485_),
    .DE(_00115_),
    .Q(\w[30][12] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][13]$_SDFFCE_PN0P_  (.D(_01486_),
    .DE(_00115_),
    .Q(\w[30][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][14]$_SDFFCE_PN0P_  (.D(_01487_),
    .DE(_00115_),
    .Q(\w[30][14] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][15]$_SDFFCE_PN0P_  (.D(_01488_),
    .DE(_00115_),
    .Q(\w[30][15] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][16]$_SDFFCE_PN0P_  (.D(_01489_),
    .DE(_00115_),
    .Q(\w[30][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][17]$_SDFFCE_PN0P_  (.D(_01490_),
    .DE(_00115_),
    .Q(\w[30][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][18]$_SDFFCE_PN0P_  (.D(_01491_),
    .DE(_00115_),
    .Q(\w[30][18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][19]$_SDFFCE_PN0P_  (.D(_01492_),
    .DE(_00115_),
    .Q(\w[30][19] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][1]$_SDFFCE_PN0P_  (.D(_01493_),
    .DE(_00115_),
    .Q(\w[30][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][20]$_SDFFCE_PN0P_  (.D(_01494_),
    .DE(_00115_),
    .Q(\w[30][20] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][21]$_SDFFCE_PN0P_  (.D(_01495_),
    .DE(_00115_),
    .Q(\w[30][21] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][22]$_SDFFCE_PN0P_  (.D(_01496_),
    .DE(_00115_),
    .Q(\w[30][22] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][23]$_SDFFCE_PN0P_  (.D(_01497_),
    .DE(_00115_),
    .Q(\w[30][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][24]$_SDFFCE_PN0P_  (.D(_01498_),
    .DE(_00115_),
    .Q(\w[30][24] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][25]$_SDFFCE_PN0P_  (.D(_01499_),
    .DE(_00115_),
    .Q(\w[30][25] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][26]$_SDFFCE_PN0P_  (.D(_01500_),
    .DE(_00115_),
    .Q(\w[30][26] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][27]$_SDFFCE_PN0P_  (.D(_01501_),
    .DE(_00115_),
    .Q(\w[30][27] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][28]$_SDFFCE_PN0P_  (.D(_01502_),
    .DE(_00115_),
    .Q(\w[30][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][29]$_SDFFCE_PN0P_  (.D(_01503_),
    .DE(_00115_),
    .Q(\w[30][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][2]$_SDFFCE_PN0P_  (.D(_01504_),
    .DE(_00115_),
    .Q(\w[30][2] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][30]$_SDFFCE_PN0P_  (.D(_01505_),
    .DE(_00115_),
    .Q(\w[30][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][31]$_SDFFCE_PN0P_  (.D(_01506_),
    .DE(_00115_),
    .Q(\w[30][31] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][3]$_SDFFCE_PN0P_  (.D(_01507_),
    .DE(_00115_),
    .Q(\w[30][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][4]$_SDFFCE_PN0P_  (.D(_01508_),
    .DE(_00115_),
    .Q(\w[30][4] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][5]$_SDFFCE_PN0P_  (.D(_01509_),
    .DE(_00115_),
    .Q(\w[30][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][6]$_SDFFCE_PN0P_  (.D(_01510_),
    .DE(_00115_),
    .Q(\w[30][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][7]$_SDFFCE_PN0P_  (.D(_01511_),
    .DE(_00115_),
    .Q(\w[30][7] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][8]$_SDFFCE_PN0P_  (.D(_01512_),
    .DE(_00115_),
    .Q(\w[30][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][9]$_SDFFCE_PN0P_  (.D(_01513_),
    .DE(_00115_),
    .Q(\w[30][9] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][0]$_SDFFCE_PN0P_  (.D(_01514_),
    .DE(_00084_),
    .Q(\w[31][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][10]$_SDFFCE_PN0P_  (.D(_01515_),
    .DE(_00084_),
    .Q(\w[31][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][11]$_SDFFCE_PN0P_  (.D(_01516_),
    .DE(_00084_),
    .Q(\w[31][11] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][12]$_SDFFCE_PN0P_  (.D(_01517_),
    .DE(_00084_),
    .Q(\w[31][12] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][13]$_SDFFCE_PN0P_  (.D(_01518_),
    .DE(_00084_),
    .Q(\w[31][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][14]$_SDFFCE_PN0P_  (.D(_01519_),
    .DE(_00084_),
    .Q(\w[31][14] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][15]$_SDFFCE_PN0P_  (.D(_01520_),
    .DE(_00084_),
    .Q(\w[31][15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][16]$_SDFFCE_PN0P_  (.D(_01521_),
    .DE(_00084_),
    .Q(\w[31][16] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][17]$_SDFFCE_PN0P_  (.D(_01522_),
    .DE(_00084_),
    .Q(\w[31][17] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][18]$_SDFFCE_PN0P_  (.D(_01523_),
    .DE(_00084_),
    .Q(\w[31][18] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][19]$_SDFFCE_PN0P_  (.D(_01524_),
    .DE(_00084_),
    .Q(\w[31][19] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][1]$_SDFFCE_PN0P_  (.D(_01525_),
    .DE(_00084_),
    .Q(\w[31][1] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][20]$_SDFFCE_PN0P_  (.D(_01526_),
    .DE(_00084_),
    .Q(\w[31][20] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][21]$_SDFFCE_PN0P_  (.D(_01527_),
    .DE(_00084_),
    .Q(\w[31][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][22]$_SDFFCE_PN0P_  (.D(_01528_),
    .DE(_00084_),
    .Q(\w[31][22] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][23]$_SDFFCE_PN0P_  (.D(_01529_),
    .DE(_00084_),
    .Q(\w[31][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][24]$_SDFFCE_PN0P_  (.D(_01530_),
    .DE(_00084_),
    .Q(\w[31][24] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][25]$_SDFFCE_PN0P_  (.D(_01531_),
    .DE(_00084_),
    .Q(\w[31][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][26]$_SDFFCE_PN0P_  (.D(_01532_),
    .DE(_00084_),
    .Q(\w[31][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][27]$_SDFFCE_PN0P_  (.D(_01533_),
    .DE(_00084_),
    .Q(\w[31][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][28]$_SDFFCE_PN0P_  (.D(_01534_),
    .DE(_00084_),
    .Q(\w[31][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][29]$_SDFFCE_PN0P_  (.D(_01535_),
    .DE(_00084_),
    .Q(\w[31][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][2]$_SDFFCE_PN0P_  (.D(_01536_),
    .DE(_00084_),
    .Q(\w[31][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][30]$_SDFFCE_PN0P_  (.D(_01537_),
    .DE(_00084_),
    .Q(\w[31][30] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][31]$_SDFFCE_PN0P_  (.D(_01538_),
    .DE(_00084_),
    .Q(\w[31][31] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][3]$_SDFFCE_PN0P_  (.D(_01539_),
    .DE(_00084_),
    .Q(\w[31][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][4]$_SDFFCE_PN0P_  (.D(_01540_),
    .DE(_00084_),
    .Q(\w[31][4] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][5]$_SDFFCE_PN0P_  (.D(_01541_),
    .DE(_00084_),
    .Q(\w[31][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][6]$_SDFFCE_PN0P_  (.D(_01542_),
    .DE(_00084_),
    .Q(\w[31][6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][7]$_SDFFCE_PN0P_  (.D(_01543_),
    .DE(_00084_),
    .Q(\w[31][7] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][8]$_SDFFCE_PN0P_  (.D(_01544_),
    .DE(_00084_),
    .Q(\w[31][8] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][9]$_SDFFCE_PN0P_  (.D(_01545_),
    .DE(_00084_),
    .Q(\w[31][9] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][0]$_SDFFCE_PN0P_  (.D(_01546_),
    .DE(_00114_),
    .Q(\w[32][0] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][10]$_SDFFCE_PN0P_  (.D(_01547_),
    .DE(_00114_),
    .Q(\w[32][10] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][11]$_SDFFCE_PN0P_  (.D(_01548_),
    .DE(_00114_),
    .Q(\w[32][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][12]$_SDFFCE_PN0P_  (.D(_01549_),
    .DE(_00114_),
    .Q(\w[32][12] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][13]$_SDFFCE_PN0P_  (.D(_01550_),
    .DE(_00114_),
    .Q(\w[32][13] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][14]$_SDFFCE_PN0P_  (.D(_01551_),
    .DE(_00114_),
    .Q(\w[32][14] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][15]$_SDFFCE_PN0P_  (.D(_01552_),
    .DE(_00114_),
    .Q(\w[32][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][16]$_SDFFCE_PN0P_  (.D(_01553_),
    .DE(_00114_),
    .Q(\w[32][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][17]$_SDFFCE_PN0P_  (.D(_01554_),
    .DE(_00114_),
    .Q(\w[32][17] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][18]$_SDFFCE_PN0P_  (.D(_01555_),
    .DE(_00114_),
    .Q(\w[32][18] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][19]$_SDFFCE_PN0P_  (.D(_01556_),
    .DE(_00114_),
    .Q(\w[32][19] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][1]$_SDFFCE_PN0P_  (.D(_01557_),
    .DE(_00114_),
    .Q(\w[32][1] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][20]$_SDFFCE_PN0P_  (.D(_01558_),
    .DE(_00114_),
    .Q(\w[32][20] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][21]$_SDFFCE_PN0P_  (.D(_01559_),
    .DE(_00114_),
    .Q(\w[32][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][22]$_SDFFCE_PN0P_  (.D(_01560_),
    .DE(_00114_),
    .Q(\w[32][22] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][23]$_SDFFCE_PN0P_  (.D(_01561_),
    .DE(_00114_),
    .Q(\w[32][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][24]$_SDFFCE_PN0P_  (.D(_01562_),
    .DE(_00114_),
    .Q(\w[32][24] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][25]$_SDFFCE_PN0P_  (.D(_01563_),
    .DE(_00114_),
    .Q(\w[32][25] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][26]$_SDFFCE_PN0P_  (.D(_01564_),
    .DE(_00114_),
    .Q(\w[32][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][27]$_SDFFCE_PN0P_  (.D(_01565_),
    .DE(_00114_),
    .Q(\w[32][27] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][28]$_SDFFCE_PN0P_  (.D(_01566_),
    .DE(_00114_),
    .Q(\w[32][28] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][29]$_SDFFCE_PN0P_  (.D(_01567_),
    .DE(_00114_),
    .Q(\w[32][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][2]$_SDFFCE_PN0P_  (.D(_01568_),
    .DE(_00114_),
    .Q(\w[32][2] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][30]$_SDFFCE_PN0P_  (.D(_01569_),
    .DE(_00114_),
    .Q(\w[32][30] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][31]$_SDFFCE_PN0P_  (.D(_01570_),
    .DE(_00114_),
    .Q(\w[32][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][3]$_SDFFCE_PN0P_  (.D(_01571_),
    .DE(_00114_),
    .Q(\w[32][3] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][4]$_SDFFCE_PN0P_  (.D(_01572_),
    .DE(_00114_),
    .Q(\w[32][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][5]$_SDFFCE_PN0P_  (.D(_01573_),
    .DE(_00114_),
    .Q(\w[32][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][6]$_SDFFCE_PN0P_  (.D(_01574_),
    .DE(_00114_),
    .Q(\w[32][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][7]$_SDFFCE_PN0P_  (.D(_01575_),
    .DE(_00114_),
    .Q(\w[32][7] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][8]$_SDFFCE_PN0P_  (.D(_01576_),
    .DE(_00114_),
    .Q(\w[32][8] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][9]$_SDFFCE_PN0P_  (.D(_01577_),
    .DE(_00114_),
    .Q(\w[32][9] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][0]$_SDFFCE_PN0P_  (.D(_01578_),
    .DE(_00083_),
    .Q(\w[33][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][10]$_SDFFCE_PN0P_  (.D(_01579_),
    .DE(_00083_),
    .Q(\w[33][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][11]$_SDFFCE_PN0P_  (.D(_01580_),
    .DE(_00083_),
    .Q(\w[33][11] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][12]$_SDFFCE_PN0P_  (.D(_01581_),
    .DE(_00083_),
    .Q(\w[33][12] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][13]$_SDFFCE_PN0P_  (.D(_01582_),
    .DE(_00083_),
    .Q(\w[33][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][14]$_SDFFCE_PN0P_  (.D(_01583_),
    .DE(_00083_),
    .Q(\w[33][14] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][15]$_SDFFCE_PN0P_  (.D(_01584_),
    .DE(_00083_),
    .Q(\w[33][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][16]$_SDFFCE_PN0P_  (.D(_01585_),
    .DE(_00083_),
    .Q(\w[33][16] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][17]$_SDFFCE_PN0P_  (.D(_01586_),
    .DE(_00083_),
    .Q(\w[33][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][18]$_SDFFCE_PN0P_  (.D(_01587_),
    .DE(_00083_),
    .Q(\w[33][18] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][19]$_SDFFCE_PN0P_  (.D(_01588_),
    .DE(_00083_),
    .Q(\w[33][19] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][1]$_SDFFCE_PN0P_  (.D(_01589_),
    .DE(_00083_),
    .Q(\w[33][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][20]$_SDFFCE_PN0P_  (.D(_01590_),
    .DE(_00083_),
    .Q(\w[33][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][21]$_SDFFCE_PN0P_  (.D(_01591_),
    .DE(_00083_),
    .Q(\w[33][21] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][22]$_SDFFCE_PN0P_  (.D(_01592_),
    .DE(_00083_),
    .Q(\w[33][22] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][23]$_SDFFCE_PN0P_  (.D(_01593_),
    .DE(_00083_),
    .Q(\w[33][23] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][24]$_SDFFCE_PN0P_  (.D(_01594_),
    .DE(_00083_),
    .Q(\w[33][24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][25]$_SDFFCE_PN0P_  (.D(_01595_),
    .DE(_00083_),
    .Q(\w[33][25] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][26]$_SDFFCE_PN0P_  (.D(_01596_),
    .DE(_00083_),
    .Q(\w[33][26] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][27]$_SDFFCE_PN0P_  (.D(_01597_),
    .DE(_00083_),
    .Q(\w[33][27] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][28]$_SDFFCE_PN0P_  (.D(_01598_),
    .DE(_00083_),
    .Q(\w[33][28] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][29]$_SDFFCE_PN0P_  (.D(_01599_),
    .DE(_00083_),
    .Q(\w[33][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][2]$_SDFFCE_PN0P_  (.D(_01600_),
    .DE(_00083_),
    .Q(\w[33][2] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][30]$_SDFFCE_PN0P_  (.D(_01601_),
    .DE(_00083_),
    .Q(\w[33][30] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][31]$_SDFFCE_PN0P_  (.D(_01602_),
    .DE(_00083_),
    .Q(\w[33][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][3]$_SDFFCE_PN0P_  (.D(_01603_),
    .DE(_00083_),
    .Q(\w[33][3] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][4]$_SDFFCE_PN0P_  (.D(_01604_),
    .DE(_00083_),
    .Q(\w[33][4] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][5]$_SDFFCE_PN0P_  (.D(_01605_),
    .DE(_00083_),
    .Q(\w[33][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][6]$_SDFFCE_PN0P_  (.D(_01606_),
    .DE(_00083_),
    .Q(\w[33][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][7]$_SDFFCE_PN0P_  (.D(_01607_),
    .DE(_00083_),
    .Q(\w[33][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][8]$_SDFFCE_PN0P_  (.D(_01608_),
    .DE(_00083_),
    .Q(\w[33][8] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][9]$_SDFFCE_PN0P_  (.D(_01609_),
    .DE(_00083_),
    .Q(\w[33][9] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][0]$_SDFFCE_PN0P_  (.D(_01610_),
    .DE(_00113_),
    .Q(\w[34][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][10]$_SDFFCE_PN0P_  (.D(_01611_),
    .DE(_00113_),
    .Q(\w[34][10] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][11]$_SDFFCE_PN0P_  (.D(_01612_),
    .DE(_00113_),
    .Q(\w[34][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][12]$_SDFFCE_PN0P_  (.D(_01613_),
    .DE(_00113_),
    .Q(\w[34][12] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][13]$_SDFFCE_PN0P_  (.D(_01614_),
    .DE(_00113_),
    .Q(\w[34][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][14]$_SDFFCE_PN0P_  (.D(_01615_),
    .DE(_00113_),
    .Q(\w[34][14] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][15]$_SDFFCE_PN0P_  (.D(_01616_),
    .DE(_00113_),
    .Q(\w[34][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][16]$_SDFFCE_PN0P_  (.D(_01617_),
    .DE(_00113_),
    .Q(\w[34][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][17]$_SDFFCE_PN0P_  (.D(_01618_),
    .DE(_00113_),
    .Q(\w[34][17] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][18]$_SDFFCE_PN0P_  (.D(_01619_),
    .DE(_00113_),
    .Q(\w[34][18] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][19]$_SDFFCE_PN0P_  (.D(_01620_),
    .DE(_00113_),
    .Q(\w[34][19] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][1]$_SDFFCE_PN0P_  (.D(_01621_),
    .DE(_00113_),
    .Q(\w[34][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][20]$_SDFFCE_PN0P_  (.D(_01622_),
    .DE(_00113_),
    .Q(\w[34][20] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][21]$_SDFFCE_PN0P_  (.D(_01623_),
    .DE(_00113_),
    .Q(\w[34][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][22]$_SDFFCE_PN0P_  (.D(_01624_),
    .DE(_00113_),
    .Q(\w[34][22] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][23]$_SDFFCE_PN0P_  (.D(_01625_),
    .DE(_00113_),
    .Q(\w[34][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][24]$_SDFFCE_PN0P_  (.D(_01626_),
    .DE(_00113_),
    .Q(\w[34][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][25]$_SDFFCE_PN0P_  (.D(_01627_),
    .DE(_00113_),
    .Q(\w[34][25] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][26]$_SDFFCE_PN0P_  (.D(_01628_),
    .DE(_00113_),
    .Q(\w[34][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][27]$_SDFFCE_PN0P_  (.D(_01629_),
    .DE(_00113_),
    .Q(\w[34][27] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][28]$_SDFFCE_PN0P_  (.D(_01630_),
    .DE(_00113_),
    .Q(\w[34][28] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][29]$_SDFFCE_PN0P_  (.D(_01631_),
    .DE(_00113_),
    .Q(\w[34][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][2]$_SDFFCE_PN0P_  (.D(_01632_),
    .DE(_00113_),
    .Q(\w[34][2] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][30]$_SDFFCE_PN0P_  (.D(_01633_),
    .DE(_00113_),
    .Q(\w[34][30] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][31]$_SDFFCE_PN0P_  (.D(_01634_),
    .DE(_00113_),
    .Q(\w[34][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][3]$_SDFFCE_PN0P_  (.D(_01635_),
    .DE(_00113_),
    .Q(\w[34][3] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][4]$_SDFFCE_PN0P_  (.D(_01636_),
    .DE(_00113_),
    .Q(\w[34][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][5]$_SDFFCE_PN0P_  (.D(_01637_),
    .DE(_00113_),
    .Q(\w[34][5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][6]$_SDFFCE_PN0P_  (.D(_01638_),
    .DE(_00113_),
    .Q(\w[34][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][7]$_SDFFCE_PN0P_  (.D(_01639_),
    .DE(_00113_),
    .Q(\w[34][7] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][8]$_SDFFCE_PN0P_  (.D(_01640_),
    .DE(_00113_),
    .Q(\w[34][8] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][9]$_SDFFCE_PN0P_  (.D(_01641_),
    .DE(_00113_),
    .Q(\w[34][9] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][0]$_SDFFCE_PN0P_  (.D(_01642_),
    .DE(_00082_),
    .Q(\w[35][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][10]$_SDFFCE_PN0P_  (.D(_01643_),
    .DE(_00082_),
    .Q(\w[35][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][11]$_SDFFCE_PN0P_  (.D(_01644_),
    .DE(_00082_),
    .Q(\w[35][11] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][12]$_SDFFCE_PN0P_  (.D(_01645_),
    .DE(_00082_),
    .Q(\w[35][12] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][13]$_SDFFCE_PN0P_  (.D(_01646_),
    .DE(_00082_),
    .Q(\w[35][13] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][14]$_SDFFCE_PN0P_  (.D(_01647_),
    .DE(_00082_),
    .Q(\w[35][14] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][15]$_SDFFCE_PN0P_  (.D(_01648_),
    .DE(_00082_),
    .Q(\w[35][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][16]$_SDFFCE_PN0P_  (.D(_01649_),
    .DE(_00082_),
    .Q(\w[35][16] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][17]$_SDFFCE_PN0P_  (.D(_01650_),
    .DE(_00082_),
    .Q(\w[35][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][18]$_SDFFCE_PN0P_  (.D(_01651_),
    .DE(_00082_),
    .Q(\w[35][18] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][19]$_SDFFCE_PN0P_  (.D(_01652_),
    .DE(_00082_),
    .Q(\w[35][19] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][1]$_SDFFCE_PN0P_  (.D(_01653_),
    .DE(_00082_),
    .Q(\w[35][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][20]$_SDFFCE_PN0P_  (.D(_01654_),
    .DE(_00082_),
    .Q(\w[35][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][21]$_SDFFCE_PN0P_  (.D(_01655_),
    .DE(_00082_),
    .Q(\w[35][21] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][22]$_SDFFCE_PN0P_  (.D(_01656_),
    .DE(_00082_),
    .Q(\w[35][22] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][23]$_SDFFCE_PN0P_  (.D(_01657_),
    .DE(_00082_),
    .Q(\w[35][23] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][24]$_SDFFCE_PN0P_  (.D(_01658_),
    .DE(_00082_),
    .Q(\w[35][24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][25]$_SDFFCE_PN0P_  (.D(_01659_),
    .DE(_00082_),
    .Q(\w[35][25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][26]$_SDFFCE_PN0P_  (.D(_01660_),
    .DE(_00082_),
    .Q(\w[35][26] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][27]$_SDFFCE_PN0P_  (.D(_01661_),
    .DE(_00082_),
    .Q(\w[35][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][28]$_SDFFCE_PN0P_  (.D(_01662_),
    .DE(_00082_),
    .Q(\w[35][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][29]$_SDFFCE_PN0P_  (.D(_01663_),
    .DE(_00082_),
    .Q(\w[35][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][2]$_SDFFCE_PN0P_  (.D(_01664_),
    .DE(_00082_),
    .Q(\w[35][2] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][30]$_SDFFCE_PN0P_  (.D(_01665_),
    .DE(_00082_),
    .Q(\w[35][30] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][31]$_SDFFCE_PN0P_  (.D(_01666_),
    .DE(_00082_),
    .Q(\w[35][31] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][3]$_SDFFCE_PN0P_  (.D(_01667_),
    .DE(_00082_),
    .Q(\w[35][3] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][4]$_SDFFCE_PN0P_  (.D(_01668_),
    .DE(_00082_),
    .Q(\w[35][4] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][5]$_SDFFCE_PN0P_  (.D(_01669_),
    .DE(_00082_),
    .Q(\w[35][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][6]$_SDFFCE_PN0P_  (.D(_01670_),
    .DE(_00082_),
    .Q(\w[35][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][7]$_SDFFCE_PN0P_  (.D(_01671_),
    .DE(_00082_),
    .Q(\w[35][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][8]$_SDFFCE_PN0P_  (.D(_01672_),
    .DE(_00082_),
    .Q(\w[35][8] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][9]$_SDFFCE_PN0P_  (.D(_01673_),
    .DE(_00082_),
    .Q(\w[35][9] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][0]$_SDFFCE_PN0P_  (.D(_01674_),
    .DE(_00112_),
    .Q(\w[36][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][10]$_SDFFCE_PN0P_  (.D(_01675_),
    .DE(_00112_),
    .Q(\w[36][10] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][11]$_SDFFCE_PN0P_  (.D(_01676_),
    .DE(_00112_),
    .Q(\w[36][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][12]$_SDFFCE_PN0P_  (.D(_01677_),
    .DE(_00112_),
    .Q(\w[36][12] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][13]$_SDFFCE_PN0P_  (.D(_01678_),
    .DE(_00112_),
    .Q(\w[36][13] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][14]$_SDFFCE_PN0P_  (.D(_01679_),
    .DE(_00112_),
    .Q(\w[36][14] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][15]$_SDFFCE_PN0P_  (.D(_01680_),
    .DE(_00112_),
    .Q(\w[36][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][16]$_SDFFCE_PN0P_  (.D(_01681_),
    .DE(_00112_),
    .Q(\w[36][16] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][17]$_SDFFCE_PN0P_  (.D(_01682_),
    .DE(_00112_),
    .Q(\w[36][17] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][18]$_SDFFCE_PN0P_  (.D(_01683_),
    .DE(_00112_),
    .Q(\w[36][18] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][19]$_SDFFCE_PN0P_  (.D(_01684_),
    .DE(_00112_),
    .Q(\w[36][19] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][1]$_SDFFCE_PN0P_  (.D(_01685_),
    .DE(_00112_),
    .Q(\w[36][1] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][20]$_SDFFCE_PN0P_  (.D(_01686_),
    .DE(_00112_),
    .Q(\w[36][20] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][21]$_SDFFCE_PN0P_  (.D(_01687_),
    .DE(_00112_),
    .Q(\w[36][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][22]$_SDFFCE_PN0P_  (.D(_01688_),
    .DE(_00112_),
    .Q(\w[36][22] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][23]$_SDFFCE_PN0P_  (.D(_01689_),
    .DE(_00112_),
    .Q(\w[36][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][24]$_SDFFCE_PN0P_  (.D(_01690_),
    .DE(_00112_),
    .Q(\w[36][24] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][25]$_SDFFCE_PN0P_  (.D(_01691_),
    .DE(_00112_),
    .Q(\w[36][25] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][26]$_SDFFCE_PN0P_  (.D(_01692_),
    .DE(_00112_),
    .Q(\w[36][26] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][27]$_SDFFCE_PN0P_  (.D(_01693_),
    .DE(_00112_),
    .Q(\w[36][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][28]$_SDFFCE_PN0P_  (.D(_01694_),
    .DE(_00112_),
    .Q(\w[36][28] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][29]$_SDFFCE_PN0P_  (.D(_01695_),
    .DE(_00112_),
    .Q(\w[36][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][2]$_SDFFCE_PN0P_  (.D(_01696_),
    .DE(_00112_),
    .Q(\w[36][2] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][30]$_SDFFCE_PN0P_  (.D(_01697_),
    .DE(_00112_),
    .Q(\w[36][30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][31]$_SDFFCE_PN0P_  (.D(_01698_),
    .DE(_00112_),
    .Q(\w[36][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][3]$_SDFFCE_PN0P_  (.D(_01699_),
    .DE(_00112_),
    .Q(\w[36][3] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][4]$_SDFFCE_PN0P_  (.D(_01700_),
    .DE(_00112_),
    .Q(\w[36][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][5]$_SDFFCE_PN0P_  (.D(_01701_),
    .DE(_00112_),
    .Q(\w[36][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][6]$_SDFFCE_PN0P_  (.D(_01702_),
    .DE(_00112_),
    .Q(\w[36][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][7]$_SDFFCE_PN0P_  (.D(_01703_),
    .DE(_00112_),
    .Q(\w[36][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][8]$_SDFFCE_PN0P_  (.D(_01704_),
    .DE(_00112_),
    .Q(\w[36][8] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][9]$_SDFFCE_PN0P_  (.D(_01705_),
    .DE(_00112_),
    .Q(\w[36][9] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][0]$_SDFFCE_PN0P_  (.D(_01706_),
    .DE(_00081_),
    .Q(\w[37][0] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][10]$_SDFFCE_PN0P_  (.D(_01707_),
    .DE(_00081_),
    .Q(\w[37][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][11]$_SDFFCE_PN0P_  (.D(_01708_),
    .DE(_00081_),
    .Q(\w[37][11] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][12]$_SDFFCE_PN0P_  (.D(_01709_),
    .DE(_00081_),
    .Q(\w[37][12] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][13]$_SDFFCE_PN0P_  (.D(_01710_),
    .DE(_00081_),
    .Q(\w[37][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][14]$_SDFFCE_PN0P_  (.D(_01711_),
    .DE(_00081_),
    .Q(\w[37][14] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][15]$_SDFFCE_PN0P_  (.D(_01712_),
    .DE(_00081_),
    .Q(\w[37][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][16]$_SDFFCE_PN0P_  (.D(_01713_),
    .DE(_00081_),
    .Q(\w[37][16] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][17]$_SDFFCE_PN0P_  (.D(_01714_),
    .DE(_00081_),
    .Q(\w[37][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][18]$_SDFFCE_PN0P_  (.D(_01715_),
    .DE(_00081_),
    .Q(\w[37][18] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][19]$_SDFFCE_PN0P_  (.D(_01716_),
    .DE(_00081_),
    .Q(\w[37][19] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][1]$_SDFFCE_PN0P_  (.D(_01717_),
    .DE(_00081_),
    .Q(\w[37][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][20]$_SDFFCE_PN0P_  (.D(_01718_),
    .DE(_00081_),
    .Q(\w[37][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][21]$_SDFFCE_PN0P_  (.D(_01719_),
    .DE(_00081_),
    .Q(\w[37][21] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][22]$_SDFFCE_PN0P_  (.D(_01720_),
    .DE(_00081_),
    .Q(\w[37][22] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][23]$_SDFFCE_PN0P_  (.D(_01721_),
    .DE(_00081_),
    .Q(\w[37][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][24]$_SDFFCE_PN0P_  (.D(_01722_),
    .DE(_00081_),
    .Q(\w[37][24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][25]$_SDFFCE_PN0P_  (.D(_01723_),
    .DE(_00081_),
    .Q(\w[37][25] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][26]$_SDFFCE_PN0P_  (.D(_01724_),
    .DE(_00081_),
    .Q(\w[37][26] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][27]$_SDFFCE_PN0P_  (.D(_01725_),
    .DE(_00081_),
    .Q(\w[37][27] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][28]$_SDFFCE_PN0P_  (.D(_01726_),
    .DE(_00081_),
    .Q(\w[37][28] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][29]$_SDFFCE_PN0P_  (.D(_01727_),
    .DE(_00081_),
    .Q(\w[37][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][2]$_SDFFCE_PN0P_  (.D(_01728_),
    .DE(_00081_),
    .Q(\w[37][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][30]$_SDFFCE_PN0P_  (.D(_01729_),
    .DE(_00081_),
    .Q(\w[37][30] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][31]$_SDFFCE_PN0P_  (.D(_01730_),
    .DE(_00081_),
    .Q(\w[37][31] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][3]$_SDFFCE_PN0P_  (.D(_01731_),
    .DE(_00081_),
    .Q(\w[37][3] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][4]$_SDFFCE_PN0P_  (.D(_01732_),
    .DE(_00081_),
    .Q(\w[37][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][5]$_SDFFCE_PN0P_  (.D(_01733_),
    .DE(_00081_),
    .Q(\w[37][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][6]$_SDFFCE_PN0P_  (.D(_01734_),
    .DE(_00081_),
    .Q(\w[37][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][7]$_SDFFCE_PN0P_  (.D(_01735_),
    .DE(_00081_),
    .Q(\w[37][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][8]$_SDFFCE_PN0P_  (.D(_01736_),
    .DE(_00081_),
    .Q(\w[37][8] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][9]$_SDFFCE_PN0P_  (.D(_01737_),
    .DE(_00081_),
    .Q(\w[37][9] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][0]$_SDFFCE_PN0P_  (.D(_01738_),
    .DE(_00111_),
    .Q(\w[38][0] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][10]$_SDFFCE_PN0P_  (.D(_01739_),
    .DE(_00111_),
    .Q(\w[38][10] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][11]$_SDFFCE_PN0P_  (.D(_01740_),
    .DE(_00111_),
    .Q(\w[38][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][12]$_SDFFCE_PN0P_  (.D(_01741_),
    .DE(_00111_),
    .Q(\w[38][12] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][13]$_SDFFCE_PN0P_  (.D(_01742_),
    .DE(_00111_),
    .Q(\w[38][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][14]$_SDFFCE_PN0P_  (.D(_01743_),
    .DE(_00111_),
    .Q(\w[38][14] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][15]$_SDFFCE_PN0P_  (.D(_01744_),
    .DE(_00111_),
    .Q(\w[38][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][16]$_SDFFCE_PN0P_  (.D(_01745_),
    .DE(_00111_),
    .Q(\w[38][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][17]$_SDFFCE_PN0P_  (.D(_01746_),
    .DE(_00111_),
    .Q(\w[38][17] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][18]$_SDFFCE_PN0P_  (.D(_01747_),
    .DE(_00111_),
    .Q(\w[38][18] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][19]$_SDFFCE_PN0P_  (.D(_01748_),
    .DE(_00111_),
    .Q(\w[38][19] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][1]$_SDFFCE_PN0P_  (.D(_01749_),
    .DE(_00111_),
    .Q(\w[38][1] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][20]$_SDFFCE_PN0P_  (.D(_01750_),
    .DE(_00111_),
    .Q(\w[38][20] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][21]$_SDFFCE_PN0P_  (.D(_01751_),
    .DE(_00111_),
    .Q(\w[38][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][22]$_SDFFCE_PN0P_  (.D(_01752_),
    .DE(_00111_),
    .Q(\w[38][22] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][23]$_SDFFCE_PN0P_  (.D(_01753_),
    .DE(_00111_),
    .Q(\w[38][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][24]$_SDFFCE_PN0P_  (.D(_01754_),
    .DE(_00111_),
    .Q(\w[38][24] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][25]$_SDFFCE_PN0P_  (.D(_01755_),
    .DE(_00111_),
    .Q(\w[38][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][26]$_SDFFCE_PN0P_  (.D(_01756_),
    .DE(_00111_),
    .Q(\w[38][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][27]$_SDFFCE_PN0P_  (.D(_01757_),
    .DE(_00111_),
    .Q(\w[38][27] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][28]$_SDFFCE_PN0P_  (.D(_01758_),
    .DE(_00111_),
    .Q(\w[38][28] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][29]$_SDFFCE_PN0P_  (.D(_01759_),
    .DE(_00111_),
    .Q(\w[38][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][2]$_SDFFCE_PN0P_  (.D(_01760_),
    .DE(_00111_),
    .Q(\w[38][2] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][30]$_SDFFCE_PN0P_  (.D(_01761_),
    .DE(_00111_),
    .Q(\w[38][30] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][31]$_SDFFCE_PN0P_  (.D(_01762_),
    .DE(_00111_),
    .Q(\w[38][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][3]$_SDFFCE_PN0P_  (.D(_01763_),
    .DE(_00111_),
    .Q(\w[38][3] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][4]$_SDFFCE_PN0P_  (.D(_01764_),
    .DE(_00111_),
    .Q(\w[38][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][5]$_SDFFCE_PN0P_  (.D(_01765_),
    .DE(_00111_),
    .Q(\w[38][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][6]$_SDFFCE_PN0P_  (.D(_01766_),
    .DE(_00111_),
    .Q(\w[38][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][7]$_SDFFCE_PN0P_  (.D(_01767_),
    .DE(_00111_),
    .Q(\w[38][7] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][8]$_SDFFCE_PN0P_  (.D(_01768_),
    .DE(_00111_),
    .Q(\w[38][8] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][9]$_SDFFCE_PN0P_  (.D(_01769_),
    .DE(_00111_),
    .Q(\w[38][9] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][0]$_SDFFCE_PN0P_  (.D(_01770_),
    .DE(net303),
    .Q(\w[39][0] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][10]$_SDFFCE_PN0P_  (.D(_01771_),
    .DE(net304),
    .Q(\w[39][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][11]$_SDFFCE_PN0P_  (.D(_01772_),
    .DE(net304),
    .Q(\w[39][11] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][12]$_SDFFCE_PN0P_  (.D(_01773_),
    .DE(net304),
    .Q(\w[39][12] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][13]$_SDFFCE_PN0P_  (.D(_01774_),
    .DE(net304),
    .Q(\w[39][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][14]$_SDFFCE_PN0P_  (.D(_01775_),
    .DE(net303),
    .Q(\w[39][14] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][15]$_SDFFCE_PN0P_  (.D(_01776_),
    .DE(net305),
    .Q(\w[39][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][16]$_SDFFCE_PN0P_  (.D(_01777_),
    .DE(net303),
    .Q(\w[39][16] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][17]$_SDFFCE_PN0P_  (.D(_01778_),
    .DE(net303),
    .Q(\w[39][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][18]$_SDFFCE_PN0P_  (.D(_01779_),
    .DE(net303),
    .Q(\w[39][18] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][19]$_SDFFCE_PN0P_  (.D(_01780_),
    .DE(net304),
    .Q(\w[39][19] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][1]$_SDFFCE_PN0P_  (.D(_01781_),
    .DE(net303),
    .Q(\w[39][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][20]$_SDFFCE_PN0P_  (.D(_01782_),
    .DE(_00080_),
    .Q(\w[39][20] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][21]$_SDFFCE_PN0P_  (.D(_01783_),
    .DE(net304),
    .Q(\w[39][21] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][22]$_SDFFCE_PN0P_  (.D(_01784_),
    .DE(net303),
    .Q(\w[39][22] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][23]$_SDFFCE_PN0P_  (.D(_01785_),
    .DE(net304),
    .Q(\w[39][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][24]$_SDFFCE_PN0P_  (.D(_01786_),
    .DE(net305),
    .Q(\w[39][24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][25]$_SDFFCE_PN0P_  (.D(_01787_),
    .DE(net303),
    .Q(\w[39][25] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][26]$_SDFFCE_PN0P_  (.D(_01788_),
    .DE(net305),
    .Q(\w[39][26] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][27]$_SDFFCE_PN0P_  (.D(_01789_),
    .DE(net304),
    .Q(\w[39][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][28]$_SDFFCE_PN0P_  (.D(_01790_),
    .DE(net305),
    .Q(\w[39][28] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][29]$_SDFFCE_PN0P_  (.D(_01791_),
    .DE(net305),
    .Q(\w[39][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][2]$_SDFFCE_PN0P_  (.D(_01792_),
    .DE(net303),
    .Q(\w[39][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][30]$_SDFFCE_PN0P_  (.D(_01793_),
    .DE(_00080_),
    .Q(\w[39][30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][31]$_SDFFCE_PN0P_  (.D(_01794_),
    .DE(net303),
    .Q(\w[39][31] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][3]$_SDFFCE_PN0P_  (.D(_01795_),
    .DE(net305),
    .Q(\w[39][3] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][4]$_SDFFCE_PN0P_  (.D(_01796_),
    .DE(net303),
    .Q(\w[39][4] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][5]$_SDFFCE_PN0P_  (.D(_01797_),
    .DE(net305),
    .Q(\w[39][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][6]$_SDFFCE_PN0P_  (.D(_01798_),
    .DE(_00080_),
    .Q(\w[39][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][7]$_SDFFCE_PN0P_  (.D(_01799_),
    .DE(_00080_),
    .Q(\w[39][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][8]$_SDFFCE_PN0P_  (.D(_01800_),
    .DE(net304),
    .Q(\w[39][8] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][9]$_SDFFCE_PN0P_  (.D(_01801_),
    .DE(_00080_),
    .Q(\w[39][9] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][0]$_DFFE_PP_  (.D(_00417_),
    .DE(_00079_),
    .Q(\w[3][0] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][10]$_DFFE_PP_  (.D(_00418_),
    .DE(_00079_),
    .Q(\w[3][10] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][11]$_DFFE_PP_  (.D(_00419_),
    .DE(_00079_),
    .Q(\w[3][11] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][12]$_DFFE_PP_  (.D(_00420_),
    .DE(_00079_),
    .Q(\w[3][12] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][13]$_DFFE_PP_  (.D(_00421_),
    .DE(_00079_),
    .Q(\w[3][13] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][14]$_DFFE_PP_  (.D(_00422_),
    .DE(_00079_),
    .Q(\w[3][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][15]$_DFFE_PP_  (.D(_00423_),
    .DE(_00079_),
    .Q(\w[3][15] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][16]$_DFFE_PP_  (.D(_00424_),
    .DE(_00079_),
    .Q(\w[3][16] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][17]$_DFFE_PP_  (.D(_00425_),
    .DE(_00079_),
    .Q(\w[3][17] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][18]$_DFFE_PP_  (.D(_00426_),
    .DE(_00079_),
    .Q(\w[3][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][19]$_DFFE_PP_  (.D(_00427_),
    .DE(_00079_),
    .Q(\w[3][19] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][1]$_DFFE_PP_  (.D(_00428_),
    .DE(_00079_),
    .Q(\w[3][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][20]$_DFFE_PP_  (.D(_00429_),
    .DE(_00079_),
    .Q(\w[3][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][21]$_DFFE_PP_  (.D(_00430_),
    .DE(_00079_),
    .Q(\w[3][21] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][22]$_DFFE_PP_  (.D(_00431_),
    .DE(_00079_),
    .Q(\w[3][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][23]$_DFFE_PP_  (.D(_00432_),
    .DE(_00079_),
    .Q(\w[3][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][24]$_DFFE_PP_  (.D(_00433_),
    .DE(_00079_),
    .Q(\w[3][24] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][25]$_DFFE_PP_  (.D(_00434_),
    .DE(_00079_),
    .Q(\w[3][25] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][26]$_DFFE_PP_  (.D(_00435_),
    .DE(_00079_),
    .Q(\w[3][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][27]$_DFFE_PP_  (.D(_00436_),
    .DE(_00079_),
    .Q(\w[3][27] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][28]$_DFFE_PP_  (.D(_00437_),
    .DE(_00079_),
    .Q(\w[3][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][29]$_DFFE_PP_  (.D(_00438_),
    .DE(_00079_),
    .Q(\w[3][29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][2]$_DFFE_PP_  (.D(_00439_),
    .DE(_00079_),
    .Q(\w[3][2] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][30]$_DFFE_PP_  (.D(_00440_),
    .DE(_00079_),
    .Q(\w[3][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][31]$_DFFE_PP_  (.D(_00441_),
    .DE(_00079_),
    .Q(\w[3][31] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][3]$_DFFE_PP_  (.D(_00442_),
    .DE(_00079_),
    .Q(\w[3][3] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][4]$_DFFE_PP_  (.D(_00443_),
    .DE(_00079_),
    .Q(\w[3][4] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][5]$_DFFE_PP_  (.D(_00444_),
    .DE(_00079_),
    .Q(\w[3][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][6]$_DFFE_PP_  (.D(_00445_),
    .DE(_00079_),
    .Q(\w[3][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][7]$_DFFE_PP_  (.D(_00446_),
    .DE(_00079_),
    .Q(\w[3][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][8]$_DFFE_PP_  (.D(_00447_),
    .DE(_00079_),
    .Q(\w[3][8] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][9]$_DFFE_PP_  (.D(_00448_),
    .DE(_00079_),
    .Q(\w[3][9] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][0]$_SDFFCE_PN0P_  (.D(_01802_),
    .DE(_00110_),
    .Q(\w[40][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][10]$_SDFFCE_PN0P_  (.D(_01803_),
    .DE(_00110_),
    .Q(\w[40][10] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][11]$_SDFFCE_PN0P_  (.D(_01804_),
    .DE(_00110_),
    .Q(\w[40][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][12]$_SDFFCE_PN0P_  (.D(_01805_),
    .DE(_00110_),
    .Q(\w[40][12] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][13]$_SDFFCE_PN0P_  (.D(_01806_),
    .DE(_00110_),
    .Q(\w[40][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][14]$_SDFFCE_PN0P_  (.D(_01807_),
    .DE(_00110_),
    .Q(\w[40][14] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][15]$_SDFFCE_PN0P_  (.D(_01808_),
    .DE(_00110_),
    .Q(\w[40][15] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][16]$_SDFFCE_PN0P_  (.D(_01809_),
    .DE(_00110_),
    .Q(\w[40][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][17]$_SDFFCE_PN0P_  (.D(_01810_),
    .DE(_00110_),
    .Q(\w[40][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][18]$_SDFFCE_PN0P_  (.D(_01811_),
    .DE(_00110_),
    .Q(\w[40][18] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][19]$_SDFFCE_PN0P_  (.D(_01812_),
    .DE(_00110_),
    .Q(\w[40][19] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][1]$_SDFFCE_PN0P_  (.D(_01813_),
    .DE(_00110_),
    .Q(\w[40][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][20]$_SDFFCE_PN0P_  (.D(_01814_),
    .DE(_00110_),
    .Q(\w[40][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][21]$_SDFFCE_PN0P_  (.D(_01815_),
    .DE(_00110_),
    .Q(\w[40][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][22]$_SDFFCE_PN0P_  (.D(_01816_),
    .DE(_00110_),
    .Q(\w[40][22] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][23]$_SDFFCE_PN0P_  (.D(_01817_),
    .DE(_00110_),
    .Q(\w[40][23] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][24]$_SDFFCE_PN0P_  (.D(_01818_),
    .DE(_00110_),
    .Q(\w[40][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][25]$_SDFFCE_PN0P_  (.D(_01819_),
    .DE(_00110_),
    .Q(\w[40][25] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][26]$_SDFFCE_PN0P_  (.D(_01820_),
    .DE(_00110_),
    .Q(\w[40][26] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][27]$_SDFFCE_PN0P_  (.D(_01821_),
    .DE(_00110_),
    .Q(\w[40][27] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][28]$_SDFFCE_PN0P_  (.D(_01822_),
    .DE(_00110_),
    .Q(\w[40][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][29]$_SDFFCE_PN0P_  (.D(_01823_),
    .DE(_00110_),
    .Q(\w[40][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][2]$_SDFFCE_PN0P_  (.D(_01824_),
    .DE(_00110_),
    .Q(\w[40][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][30]$_SDFFCE_PN0P_  (.D(_01825_),
    .DE(_00110_),
    .Q(\w[40][30] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][31]$_SDFFCE_PN0P_  (.D(_01826_),
    .DE(_00110_),
    .Q(\w[40][31] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][3]$_SDFFCE_PN0P_  (.D(_01827_),
    .DE(_00110_),
    .Q(\w[40][3] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][4]$_SDFFCE_PN0P_  (.D(_01828_),
    .DE(_00110_),
    .Q(\w[40][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][5]$_SDFFCE_PN0P_  (.D(_01829_),
    .DE(_00110_),
    .Q(\w[40][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][6]$_SDFFCE_PN0P_  (.D(_01830_),
    .DE(_00110_),
    .Q(\w[40][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][7]$_SDFFCE_PN0P_  (.D(_01831_),
    .DE(_00110_),
    .Q(\w[40][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][8]$_SDFFCE_PN0P_  (.D(_01832_),
    .DE(_00110_),
    .Q(\w[40][8] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][9]$_SDFFCE_PN0P_  (.D(_01833_),
    .DE(_00110_),
    .Q(\w[40][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][0]$_SDFFCE_PN0P_  (.D(_01834_),
    .DE(_00078_),
    .Q(\w[41][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][10]$_SDFFCE_PN0P_  (.D(_01835_),
    .DE(_00078_),
    .Q(\w[41][10] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][11]$_SDFFCE_PN0P_  (.D(_01836_),
    .DE(_00078_),
    .Q(\w[41][11] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][12]$_SDFFCE_PN0P_  (.D(_01837_),
    .DE(_00078_),
    .Q(\w[41][12] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][13]$_SDFFCE_PN0P_  (.D(_01838_),
    .DE(_00078_),
    .Q(\w[41][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][14]$_SDFFCE_PN0P_  (.D(_01839_),
    .DE(_00078_),
    .Q(\w[41][14] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][15]$_SDFFCE_PN0P_  (.D(_01840_),
    .DE(_00078_),
    .Q(\w[41][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][16]$_SDFFCE_PN0P_  (.D(_01841_),
    .DE(_00078_),
    .Q(\w[41][16] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][17]$_SDFFCE_PN0P_  (.D(_01842_),
    .DE(_00078_),
    .Q(\w[41][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][18]$_SDFFCE_PN0P_  (.D(_01843_),
    .DE(_00078_),
    .Q(\w[41][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][19]$_SDFFCE_PN0P_  (.D(_01844_),
    .DE(_00078_),
    .Q(\w[41][19] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][1]$_SDFFCE_PN0P_  (.D(_01845_),
    .DE(_00078_),
    .Q(\w[41][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][20]$_SDFFCE_PN0P_  (.D(_01846_),
    .DE(_00078_),
    .Q(\w[41][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][21]$_SDFFCE_PN0P_  (.D(_01847_),
    .DE(_00078_),
    .Q(\w[41][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][22]$_SDFFCE_PN0P_  (.D(_01848_),
    .DE(_00078_),
    .Q(\w[41][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][23]$_SDFFCE_PN0P_  (.D(_01849_),
    .DE(_00078_),
    .Q(\w[41][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][24]$_SDFFCE_PN0P_  (.D(_01850_),
    .DE(_00078_),
    .Q(\w[41][24] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][25]$_SDFFCE_PN0P_  (.D(_01851_),
    .DE(_00078_),
    .Q(\w[41][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][26]$_SDFFCE_PN0P_  (.D(_01852_),
    .DE(_00078_),
    .Q(\w[41][26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][27]$_SDFFCE_PN0P_  (.D(_01853_),
    .DE(_00078_),
    .Q(\w[41][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][28]$_SDFFCE_PN0P_  (.D(_01854_),
    .DE(_00078_),
    .Q(\w[41][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][29]$_SDFFCE_PN0P_  (.D(_01855_),
    .DE(_00078_),
    .Q(\w[41][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][2]$_SDFFCE_PN0P_  (.D(_01856_),
    .DE(_00078_),
    .Q(\w[41][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][30]$_SDFFCE_PN0P_  (.D(_01857_),
    .DE(_00078_),
    .Q(\w[41][30] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][31]$_SDFFCE_PN0P_  (.D(_01858_),
    .DE(_00078_),
    .Q(\w[41][31] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][3]$_SDFFCE_PN0P_  (.D(_01859_),
    .DE(_00078_),
    .Q(\w[41][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][4]$_SDFFCE_PN0P_  (.D(_01860_),
    .DE(_00078_),
    .Q(\w[41][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][5]$_SDFFCE_PN0P_  (.D(_01861_),
    .DE(_00078_),
    .Q(\w[41][5] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][6]$_SDFFCE_PN0P_  (.D(_01862_),
    .DE(_00078_),
    .Q(\w[41][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][7]$_SDFFCE_PN0P_  (.D(_01863_),
    .DE(_00078_),
    .Q(\w[41][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][8]$_SDFFCE_PN0P_  (.D(_01864_),
    .DE(_00078_),
    .Q(\w[41][8] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][9]$_SDFFCE_PN0P_  (.D(_01865_),
    .DE(_00078_),
    .Q(\w[41][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][0]$_SDFFCE_PN0P_  (.D(_01866_),
    .DE(_00109_),
    .Q(\w[42][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][10]$_SDFFCE_PN0P_  (.D(_01867_),
    .DE(_00109_),
    .Q(\w[42][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][11]$_SDFFCE_PN0P_  (.D(_01868_),
    .DE(_00109_),
    .Q(\w[42][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][12]$_SDFFCE_PN0P_  (.D(_01869_),
    .DE(_00109_),
    .Q(\w[42][12] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][13]$_SDFFCE_PN0P_  (.D(_01870_),
    .DE(_00109_),
    .Q(\w[42][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][14]$_SDFFCE_PN0P_  (.D(_01871_),
    .DE(_00109_),
    .Q(\w[42][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][15]$_SDFFCE_PN0P_  (.D(_01872_),
    .DE(_00109_),
    .Q(\w[42][15] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][16]$_SDFFCE_PN0P_  (.D(_01873_),
    .DE(_00109_),
    .Q(\w[42][16] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][17]$_SDFFCE_PN0P_  (.D(_01874_),
    .DE(_00109_),
    .Q(\w[42][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][18]$_SDFFCE_PN0P_  (.D(_01875_),
    .DE(_00109_),
    .Q(\w[42][18] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][19]$_SDFFCE_PN0P_  (.D(_01876_),
    .DE(_00109_),
    .Q(\w[42][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][1]$_SDFFCE_PN0P_  (.D(_01877_),
    .DE(_00109_),
    .Q(\w[42][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][20]$_SDFFCE_PN0P_  (.D(_01878_),
    .DE(_00109_),
    .Q(\w[42][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][21]$_SDFFCE_PN0P_  (.D(_01879_),
    .DE(_00109_),
    .Q(\w[42][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][22]$_SDFFCE_PN0P_  (.D(_01880_),
    .DE(_00109_),
    .Q(\w[42][22] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][23]$_SDFFCE_PN0P_  (.D(_01881_),
    .DE(_00109_),
    .Q(\w[42][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][24]$_SDFFCE_PN0P_  (.D(_01882_),
    .DE(_00109_),
    .Q(\w[42][24] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][25]$_SDFFCE_PN0P_  (.D(_01883_),
    .DE(_00109_),
    .Q(\w[42][25] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][26]$_SDFFCE_PN0P_  (.D(_01884_),
    .DE(_00109_),
    .Q(\w[42][26] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][27]$_SDFFCE_PN0P_  (.D(_01885_),
    .DE(_00109_),
    .Q(\w[42][27] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][28]$_SDFFCE_PN0P_  (.D(_01886_),
    .DE(_00109_),
    .Q(\w[42][28] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][29]$_SDFFCE_PN0P_  (.D(_01887_),
    .DE(_00109_),
    .Q(\w[42][29] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][2]$_SDFFCE_PN0P_  (.D(_01888_),
    .DE(_00109_),
    .Q(\w[42][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][30]$_SDFFCE_PN0P_  (.D(_01889_),
    .DE(_00109_),
    .Q(\w[42][30] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][31]$_SDFFCE_PN0P_  (.D(_01890_),
    .DE(_00109_),
    .Q(\w[42][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][3]$_SDFFCE_PN0P_  (.D(_01891_),
    .DE(_00109_),
    .Q(\w[42][3] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][4]$_SDFFCE_PN0P_  (.D(_01892_),
    .DE(_00109_),
    .Q(\w[42][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][5]$_SDFFCE_PN0P_  (.D(_01893_),
    .DE(_00109_),
    .Q(\w[42][5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][6]$_SDFFCE_PN0P_  (.D(_01894_),
    .DE(_00109_),
    .Q(\w[42][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][7]$_SDFFCE_PN0P_  (.D(_01895_),
    .DE(_00109_),
    .Q(\w[42][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][8]$_SDFFCE_PN0P_  (.D(_01896_),
    .DE(_00109_),
    .Q(\w[42][8] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][9]$_SDFFCE_PN0P_  (.D(_01897_),
    .DE(_00109_),
    .Q(\w[42][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][0]$_SDFFCE_PN0P_  (.D(_01898_),
    .DE(_00077_),
    .Q(\w[43][0] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][10]$_SDFFCE_PN0P_  (.D(_01899_),
    .DE(_00077_),
    .Q(\w[43][10] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][11]$_SDFFCE_PN0P_  (.D(_01900_),
    .DE(_00077_),
    .Q(\w[43][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][12]$_SDFFCE_PN0P_  (.D(_01901_),
    .DE(_00077_),
    .Q(\w[43][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][13]$_SDFFCE_PN0P_  (.D(_01902_),
    .DE(_00077_),
    .Q(\w[43][13] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][14]$_SDFFCE_PN0P_  (.D(_01903_),
    .DE(_00077_),
    .Q(\w[43][14] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][15]$_SDFFCE_PN0P_  (.D(_01904_),
    .DE(_00077_),
    .Q(\w[43][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][16]$_SDFFCE_PN0P_  (.D(_01905_),
    .DE(_00077_),
    .Q(\w[43][16] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][17]$_SDFFCE_PN0P_  (.D(_01906_),
    .DE(_00077_),
    .Q(\w[43][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][18]$_SDFFCE_PN0P_  (.D(_01907_),
    .DE(_00077_),
    .Q(\w[43][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][19]$_SDFFCE_PN0P_  (.D(_01908_),
    .DE(_00077_),
    .Q(\w[43][19] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][1]$_SDFFCE_PN0P_  (.D(_01909_),
    .DE(_00077_),
    .Q(\w[43][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][20]$_SDFFCE_PN0P_  (.D(_01910_),
    .DE(_00077_),
    .Q(\w[43][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][21]$_SDFFCE_PN0P_  (.D(_01911_),
    .DE(_00077_),
    .Q(\w[43][21] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][22]$_SDFFCE_PN0P_  (.D(_01912_),
    .DE(_00077_),
    .Q(\w[43][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][23]$_SDFFCE_PN0P_  (.D(_01913_),
    .DE(_00077_),
    .Q(\w[43][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][24]$_SDFFCE_PN0P_  (.D(_01914_),
    .DE(_00077_),
    .Q(\w[43][24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][25]$_SDFFCE_PN0P_  (.D(_01915_),
    .DE(_00077_),
    .Q(\w[43][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][26]$_SDFFCE_PN0P_  (.D(_01916_),
    .DE(_00077_),
    .Q(\w[43][26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][27]$_SDFFCE_PN0P_  (.D(_01917_),
    .DE(_00077_),
    .Q(\w[43][27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][28]$_SDFFCE_PN0P_  (.D(_01918_),
    .DE(_00077_),
    .Q(\w[43][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][29]$_SDFFCE_PN0P_  (.D(_01919_),
    .DE(_00077_),
    .Q(\w[43][29] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][2]$_SDFFCE_PN0P_  (.D(_01920_),
    .DE(_00077_),
    .Q(\w[43][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][30]$_SDFFCE_PN0P_  (.D(_01921_),
    .DE(_00077_),
    .Q(\w[43][30] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][31]$_SDFFCE_PN0P_  (.D(_01922_),
    .DE(_00077_),
    .Q(\w[43][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][3]$_SDFFCE_PN0P_  (.D(_01923_),
    .DE(_00077_),
    .Q(\w[43][3] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][4]$_SDFFCE_PN0P_  (.D(_01924_),
    .DE(_00077_),
    .Q(\w[43][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][5]$_SDFFCE_PN0P_  (.D(_01925_),
    .DE(_00077_),
    .Q(\w[43][5] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][6]$_SDFFCE_PN0P_  (.D(_01926_),
    .DE(_00077_),
    .Q(\w[43][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][7]$_SDFFCE_PN0P_  (.D(_01927_),
    .DE(_00077_),
    .Q(\w[43][7] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][8]$_SDFFCE_PN0P_  (.D(_01928_),
    .DE(_00077_),
    .Q(\w[43][8] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][9]$_SDFFCE_PN0P_  (.D(_01929_),
    .DE(_00077_),
    .Q(\w[43][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][0]$_SDFFCE_PN0P_  (.D(_01930_),
    .DE(_00108_),
    .Q(\w[44][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][10]$_SDFFCE_PN0P_  (.D(_01931_),
    .DE(_00108_),
    .Q(\w[44][10] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][11]$_SDFFCE_PN0P_  (.D(_01932_),
    .DE(_00108_),
    .Q(\w[44][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][12]$_SDFFCE_PN0P_  (.D(_01933_),
    .DE(_00108_),
    .Q(\w[44][12] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][13]$_SDFFCE_PN0P_  (.D(_01934_),
    .DE(_00108_),
    .Q(\w[44][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][14]$_SDFFCE_PN0P_  (.D(_01935_),
    .DE(_00108_),
    .Q(\w[44][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][15]$_SDFFCE_PN0P_  (.D(_01936_),
    .DE(_00108_),
    .Q(\w[44][15] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][16]$_SDFFCE_PN0P_  (.D(_01937_),
    .DE(_00108_),
    .Q(\w[44][16] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][17]$_SDFFCE_PN0P_  (.D(_01938_),
    .DE(_00108_),
    .Q(\w[44][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][18]$_SDFFCE_PN0P_  (.D(_01939_),
    .DE(_00108_),
    .Q(\w[44][18] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][19]$_SDFFCE_PN0P_  (.D(_01940_),
    .DE(_00108_),
    .Q(\w[44][19] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][1]$_SDFFCE_PN0P_  (.D(_01941_),
    .DE(_00108_),
    .Q(\w[44][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][20]$_SDFFCE_PN0P_  (.D(_01942_),
    .DE(_00108_),
    .Q(\w[44][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][21]$_SDFFCE_PN0P_  (.D(_01943_),
    .DE(_00108_),
    .Q(\w[44][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][22]$_SDFFCE_PN0P_  (.D(_01944_),
    .DE(_00108_),
    .Q(\w[44][22] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][23]$_SDFFCE_PN0P_  (.D(_01945_),
    .DE(_00108_),
    .Q(\w[44][23] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][24]$_SDFFCE_PN0P_  (.D(_01946_),
    .DE(_00108_),
    .Q(\w[44][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][25]$_SDFFCE_PN0P_  (.D(_01947_),
    .DE(_00108_),
    .Q(\w[44][25] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][26]$_SDFFCE_PN0P_  (.D(_01948_),
    .DE(_00108_),
    .Q(\w[44][26] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][27]$_SDFFCE_PN0P_  (.D(_01949_),
    .DE(_00108_),
    .Q(\w[44][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][28]$_SDFFCE_PN0P_  (.D(_01950_),
    .DE(_00108_),
    .Q(\w[44][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][29]$_SDFFCE_PN0P_  (.D(_01951_),
    .DE(_00108_),
    .Q(\w[44][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][2]$_SDFFCE_PN0P_  (.D(_01952_),
    .DE(_00108_),
    .Q(\w[44][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][30]$_SDFFCE_PN0P_  (.D(_01953_),
    .DE(_00108_),
    .Q(\w[44][30] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][31]$_SDFFCE_PN0P_  (.D(_01954_),
    .DE(_00108_),
    .Q(\w[44][31] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][3]$_SDFFCE_PN0P_  (.D(_01955_),
    .DE(_00108_),
    .Q(\w[44][3] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][4]$_SDFFCE_PN0P_  (.D(_01956_),
    .DE(_00108_),
    .Q(\w[44][4] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][5]$_SDFFCE_PN0P_  (.D(_01957_),
    .DE(_00108_),
    .Q(\w[44][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][6]$_SDFFCE_PN0P_  (.D(_01958_),
    .DE(_00108_),
    .Q(\w[44][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][7]$_SDFFCE_PN0P_  (.D(_01959_),
    .DE(_00108_),
    .Q(\w[44][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][8]$_SDFFCE_PN0P_  (.D(_01960_),
    .DE(_00108_),
    .Q(\w[44][8] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][9]$_SDFFCE_PN0P_  (.D(_01961_),
    .DE(_00108_),
    .Q(\w[44][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][0]$_SDFFCE_PN0P_  (.D(_01962_),
    .DE(_00076_),
    .Q(\w[45][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][10]$_SDFFCE_PN0P_  (.D(_01963_),
    .DE(_00076_),
    .Q(\w[45][10] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][11]$_SDFFCE_PN0P_  (.D(_01964_),
    .DE(_00076_),
    .Q(\w[45][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][12]$_SDFFCE_PN0P_  (.D(_01965_),
    .DE(_00076_),
    .Q(\w[45][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][13]$_SDFFCE_PN0P_  (.D(_01966_),
    .DE(_00076_),
    .Q(\w[45][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][14]$_SDFFCE_PN0P_  (.D(_01967_),
    .DE(_00076_),
    .Q(\w[45][14] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][15]$_SDFFCE_PN0P_  (.D(_01968_),
    .DE(_00076_),
    .Q(\w[45][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][16]$_SDFFCE_PN0P_  (.D(_01969_),
    .DE(_00076_),
    .Q(\w[45][16] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][17]$_SDFFCE_PN0P_  (.D(_01970_),
    .DE(_00076_),
    .Q(\w[45][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][18]$_SDFFCE_PN0P_  (.D(_01971_),
    .DE(_00076_),
    .Q(\w[45][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][19]$_SDFFCE_PN0P_  (.D(_01972_),
    .DE(_00076_),
    .Q(\w[45][19] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][1]$_SDFFCE_PN0P_  (.D(_01973_),
    .DE(_00076_),
    .Q(\w[45][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][20]$_SDFFCE_PN0P_  (.D(_01974_),
    .DE(_00076_),
    .Q(\w[45][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][21]$_SDFFCE_PN0P_  (.D(_01975_),
    .DE(_00076_),
    .Q(\w[45][21] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][22]$_SDFFCE_PN0P_  (.D(_01976_),
    .DE(_00076_),
    .Q(\w[45][22] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][23]$_SDFFCE_PN0P_  (.D(_01977_),
    .DE(_00076_),
    .Q(\w[45][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][24]$_SDFFCE_PN0P_  (.D(_01978_),
    .DE(_00076_),
    .Q(\w[45][24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][25]$_SDFFCE_PN0P_  (.D(_01979_),
    .DE(_00076_),
    .Q(\w[45][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][26]$_SDFFCE_PN0P_  (.D(_01980_),
    .DE(_00076_),
    .Q(\w[45][26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][27]$_SDFFCE_PN0P_  (.D(_01981_),
    .DE(_00076_),
    .Q(\w[45][27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][28]$_SDFFCE_PN0P_  (.D(_01982_),
    .DE(_00076_),
    .Q(\w[45][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][29]$_SDFFCE_PN0P_  (.D(_01983_),
    .DE(_00076_),
    .Q(\w[45][29] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][2]$_SDFFCE_PN0P_  (.D(_01984_),
    .DE(_00076_),
    .Q(\w[45][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][30]$_SDFFCE_PN0P_  (.D(_01985_),
    .DE(_00076_),
    .Q(\w[45][30] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][31]$_SDFFCE_PN0P_  (.D(_01986_),
    .DE(_00076_),
    .Q(\w[45][31] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][3]$_SDFFCE_PN0P_  (.D(_01987_),
    .DE(_00076_),
    .Q(\w[45][3] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][4]$_SDFFCE_PN0P_  (.D(_01988_),
    .DE(_00076_),
    .Q(\w[45][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][5]$_SDFFCE_PN0P_  (.D(_01989_),
    .DE(_00076_),
    .Q(\w[45][5] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][6]$_SDFFCE_PN0P_  (.D(_01990_),
    .DE(_00076_),
    .Q(\w[45][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][7]$_SDFFCE_PN0P_  (.D(_01991_),
    .DE(_00076_),
    .Q(\w[45][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][8]$_SDFFCE_PN0P_  (.D(_01992_),
    .DE(_00076_),
    .Q(\w[45][8] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][9]$_SDFFCE_PN0P_  (.D(_01993_),
    .DE(_00076_),
    .Q(\w[45][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][0]$_SDFFCE_PN0P_  (.D(_01994_),
    .DE(_00107_),
    .Q(\w[46][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][10]$_SDFFCE_PN0P_  (.D(_01995_),
    .DE(_00107_),
    .Q(\w[46][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][11]$_SDFFCE_PN0P_  (.D(_01996_),
    .DE(_00107_),
    .Q(\w[46][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][12]$_SDFFCE_PN0P_  (.D(_01997_),
    .DE(_00107_),
    .Q(\w[46][12] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][13]$_SDFFCE_PN0P_  (.D(_01998_),
    .DE(_00107_),
    .Q(\w[46][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][14]$_SDFFCE_PN0P_  (.D(_01999_),
    .DE(_00107_),
    .Q(\w[46][14] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][15]$_SDFFCE_PN0P_  (.D(_02000_),
    .DE(_00107_),
    .Q(\w[46][15] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][16]$_SDFFCE_PN0P_  (.D(_02001_),
    .DE(_00107_),
    .Q(\w[46][16] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][17]$_SDFFCE_PN0P_  (.D(_02002_),
    .DE(_00107_),
    .Q(\w[46][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][18]$_SDFFCE_PN0P_  (.D(_02003_),
    .DE(_00107_),
    .Q(\w[46][18] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][19]$_SDFFCE_PN0P_  (.D(_02004_),
    .DE(_00107_),
    .Q(\w[46][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][1]$_SDFFCE_PN0P_  (.D(_02005_),
    .DE(_00107_),
    .Q(\w[46][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][20]$_SDFFCE_PN0P_  (.D(_02006_),
    .DE(_00107_),
    .Q(\w[46][20] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][21]$_SDFFCE_PN0P_  (.D(_02007_),
    .DE(_00107_),
    .Q(\w[46][21] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][22]$_SDFFCE_PN0P_  (.D(_02008_),
    .DE(_00107_),
    .Q(\w[46][22] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][23]$_SDFFCE_PN0P_  (.D(_02009_),
    .DE(_00107_),
    .Q(\w[46][23] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][24]$_SDFFCE_PN0P_  (.D(_02010_),
    .DE(_00107_),
    .Q(\w[46][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][25]$_SDFFCE_PN0P_  (.D(_02011_),
    .DE(_00107_),
    .Q(\w[46][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][26]$_SDFFCE_PN0P_  (.D(_02012_),
    .DE(_00107_),
    .Q(\w[46][26] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][27]$_SDFFCE_PN0P_  (.D(_02013_),
    .DE(_00107_),
    .Q(\w[46][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][28]$_SDFFCE_PN0P_  (.D(_02014_),
    .DE(_00107_),
    .Q(\w[46][28] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][29]$_SDFFCE_PN0P_  (.D(_02015_),
    .DE(_00107_),
    .Q(\w[46][29] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][2]$_SDFFCE_PN0P_  (.D(_02016_),
    .DE(_00107_),
    .Q(\w[46][2] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][30]$_SDFFCE_PN0P_  (.D(_02017_),
    .DE(_00107_),
    .Q(\w[46][30] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][31]$_SDFFCE_PN0P_  (.D(_02018_),
    .DE(_00107_),
    .Q(\w[46][31] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][3]$_SDFFCE_PN0P_  (.D(_02019_),
    .DE(_00107_),
    .Q(\w[46][3] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][4]$_SDFFCE_PN0P_  (.D(_02020_),
    .DE(_00107_),
    .Q(\w[46][4] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][5]$_SDFFCE_PN0P_  (.D(_02021_),
    .DE(_00107_),
    .Q(\w[46][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][6]$_SDFFCE_PN0P_  (.D(_02022_),
    .DE(_00107_),
    .Q(\w[46][6] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][7]$_SDFFCE_PN0P_  (.D(_02023_),
    .DE(_00107_),
    .Q(\w[46][7] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][8]$_SDFFCE_PN0P_  (.D(_02024_),
    .DE(_00107_),
    .Q(\w[46][8] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][9]$_SDFFCE_PN0P_  (.D(_02025_),
    .DE(_00107_),
    .Q(\w[46][9] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][0]$_SDFFCE_PN0P_  (.D(_02026_),
    .DE(_00075_),
    .Q(\w[47][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][10]$_SDFFCE_PN0P_  (.D(_02027_),
    .DE(_00075_),
    .Q(\w[47][10] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][11]$_SDFFCE_PN0P_  (.D(_02028_),
    .DE(_00075_),
    .Q(\w[47][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][12]$_SDFFCE_PN0P_  (.D(_02029_),
    .DE(_00075_),
    .Q(\w[47][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][13]$_SDFFCE_PN0P_  (.D(_02030_),
    .DE(_00075_),
    .Q(\w[47][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][14]$_SDFFCE_PN0P_  (.D(_02031_),
    .DE(_00075_),
    .Q(\w[47][14] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][15]$_SDFFCE_PN0P_  (.D(_02032_),
    .DE(_00075_),
    .Q(\w[47][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][16]$_SDFFCE_PN0P_  (.D(_02033_),
    .DE(_00075_),
    .Q(\w[47][16] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][17]$_SDFFCE_PN0P_  (.D(_02034_),
    .DE(_00075_),
    .Q(\w[47][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][18]$_SDFFCE_PN0P_  (.D(_02035_),
    .DE(_00075_),
    .Q(\w[47][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][19]$_SDFFCE_PN0P_  (.D(_02036_),
    .DE(_00075_),
    .Q(\w[47][19] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][1]$_SDFFCE_PN0P_  (.D(_02037_),
    .DE(_00075_),
    .Q(\w[47][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][20]$_SDFFCE_PN0P_  (.D(_02038_),
    .DE(_00075_),
    .Q(\w[47][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][21]$_SDFFCE_PN0P_  (.D(_02039_),
    .DE(_00075_),
    .Q(\w[47][21] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][22]$_SDFFCE_PN0P_  (.D(_02040_),
    .DE(_00075_),
    .Q(\w[47][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][23]$_SDFFCE_PN0P_  (.D(_02041_),
    .DE(_00075_),
    .Q(\w[47][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][24]$_SDFFCE_PN0P_  (.D(_02042_),
    .DE(_00075_),
    .Q(\w[47][24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][25]$_SDFFCE_PN0P_  (.D(_02043_),
    .DE(_00075_),
    .Q(\w[47][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][26]$_SDFFCE_PN0P_  (.D(_02044_),
    .DE(_00075_),
    .Q(\w[47][26] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][27]$_SDFFCE_PN0P_  (.D(_02045_),
    .DE(_00075_),
    .Q(\w[47][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][28]$_SDFFCE_PN0P_  (.D(_02046_),
    .DE(_00075_),
    .Q(\w[47][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][29]$_SDFFCE_PN0P_  (.D(_02047_),
    .DE(_00075_),
    .Q(\w[47][29] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][2]$_SDFFCE_PN0P_  (.D(_02048_),
    .DE(_00075_),
    .Q(\w[47][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][30]$_SDFFCE_PN0P_  (.D(_02049_),
    .DE(_00075_),
    .Q(\w[47][30] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][31]$_SDFFCE_PN0P_  (.D(_02050_),
    .DE(_00075_),
    .Q(\w[47][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][3]$_SDFFCE_PN0P_  (.D(_02051_),
    .DE(_00075_),
    .Q(\w[47][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][4]$_SDFFCE_PN0P_  (.D(_02052_),
    .DE(_00075_),
    .Q(\w[47][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][5]$_SDFFCE_PN0P_  (.D(_02053_),
    .DE(_00075_),
    .Q(\w[47][5] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][6]$_SDFFCE_PN0P_  (.D(_02054_),
    .DE(_00075_),
    .Q(\w[47][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][7]$_SDFFCE_PN0P_  (.D(_02055_),
    .DE(_00075_),
    .Q(\w[47][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][8]$_SDFFCE_PN0P_  (.D(_02056_),
    .DE(_00075_),
    .Q(\w[47][8] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][9]$_SDFFCE_PN0P_  (.D(_02057_),
    .DE(_00075_),
    .Q(\w[47][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][0]$_SDFFCE_PN0P_  (.D(_02058_),
    .DE(_00106_),
    .Q(\w[48][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][10]$_SDFFCE_PN0P_  (.D(_02059_),
    .DE(_00106_),
    .Q(\w[48][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][11]$_SDFFCE_PN0P_  (.D(_02060_),
    .DE(_00106_),
    .Q(\w[48][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][12]$_SDFFCE_PN0P_  (.D(_02061_),
    .DE(_00106_),
    .Q(\w[48][12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][13]$_SDFFCE_PN0P_  (.D(_02062_),
    .DE(_00106_),
    .Q(\w[48][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][14]$_SDFFCE_PN0P_  (.D(_02063_),
    .DE(_00106_),
    .Q(\w[48][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][15]$_SDFFCE_PN0P_  (.D(_02064_),
    .DE(_00106_),
    .Q(\w[48][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][16]$_SDFFCE_PN0P_  (.D(_02065_),
    .DE(_00106_),
    .Q(\w[48][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][17]$_SDFFCE_PN0P_  (.D(_02066_),
    .DE(_00106_),
    .Q(\w[48][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][18]$_SDFFCE_PN0P_  (.D(_02067_),
    .DE(_00106_),
    .Q(\w[48][18] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][19]$_SDFFCE_PN0P_  (.D(_02068_),
    .DE(_00106_),
    .Q(\w[48][19] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][1]$_SDFFCE_PN0P_  (.D(_02069_),
    .DE(_00106_),
    .Q(\w[48][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][20]$_SDFFCE_PN0P_  (.D(_02070_),
    .DE(_00106_),
    .Q(\w[48][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][21]$_SDFFCE_PN0P_  (.D(_02071_),
    .DE(_00106_),
    .Q(\w[48][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][22]$_SDFFCE_PN0P_  (.D(_02072_),
    .DE(_00106_),
    .Q(\w[48][22] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][23]$_SDFFCE_PN0P_  (.D(_02073_),
    .DE(_00106_),
    .Q(\w[48][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][24]$_SDFFCE_PN0P_  (.D(_02074_),
    .DE(_00106_),
    .Q(\w[48][24] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][25]$_SDFFCE_PN0P_  (.D(_02075_),
    .DE(_00106_),
    .Q(\w[48][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][26]$_SDFFCE_PN0P_  (.D(_02076_),
    .DE(_00106_),
    .Q(\w[48][26] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][27]$_SDFFCE_PN0P_  (.D(_02077_),
    .DE(_00106_),
    .Q(\w[48][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][28]$_SDFFCE_PN0P_  (.D(_02078_),
    .DE(_00106_),
    .Q(\w[48][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][29]$_SDFFCE_PN0P_  (.D(_02079_),
    .DE(_00106_),
    .Q(\w[48][29] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][2]$_SDFFCE_PN0P_  (.D(_02080_),
    .DE(_00106_),
    .Q(\w[48][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][30]$_SDFFCE_PN0P_  (.D(_02081_),
    .DE(_00106_),
    .Q(\w[48][30] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][31]$_SDFFCE_PN0P_  (.D(_02082_),
    .DE(_00106_),
    .Q(\w[48][31] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][3]$_SDFFCE_PN0P_  (.D(_02083_),
    .DE(_00106_),
    .Q(\w[48][3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][4]$_SDFFCE_PN0P_  (.D(_02084_),
    .DE(_00106_),
    .Q(\w[48][4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][5]$_SDFFCE_PN0P_  (.D(_02085_),
    .DE(_00106_),
    .Q(\w[48][5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][6]$_SDFFCE_PN0P_  (.D(_02086_),
    .DE(_00106_),
    .Q(\w[48][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][7]$_SDFFCE_PN0P_  (.D(_02087_),
    .DE(_00106_),
    .Q(\w[48][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][8]$_SDFFCE_PN0P_  (.D(_02088_),
    .DE(_00106_),
    .Q(\w[48][8] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][9]$_SDFFCE_PN0P_  (.D(_02089_),
    .DE(_00106_),
    .Q(\w[48][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][0]$_SDFFCE_PN0P_  (.D(_02090_),
    .DE(_00074_),
    .Q(\w[49][0] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][10]$_SDFFCE_PN0P_  (.D(_02091_),
    .DE(_00074_),
    .Q(\w[49][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][11]$_SDFFCE_PN0P_  (.D(_02092_),
    .DE(_00074_),
    .Q(\w[49][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][12]$_SDFFCE_PN0P_  (.D(_02093_),
    .DE(_00074_),
    .Q(\w[49][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][13]$_SDFFCE_PN0P_  (.D(_02094_),
    .DE(_00074_),
    .Q(\w[49][13] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][14]$_SDFFCE_PN0P_  (.D(_02095_),
    .DE(_00074_),
    .Q(\w[49][14] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][15]$_SDFFCE_PN0P_  (.D(_02096_),
    .DE(_00074_),
    .Q(\w[49][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][16]$_SDFFCE_PN0P_  (.D(_02097_),
    .DE(_00074_),
    .Q(\w[49][16] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][17]$_SDFFCE_PN0P_  (.D(_02098_),
    .DE(_00074_),
    .Q(\w[49][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][18]$_SDFFCE_PN0P_  (.D(_02099_),
    .DE(_00074_),
    .Q(\w[49][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][19]$_SDFFCE_PN0P_  (.D(_02100_),
    .DE(_00074_),
    .Q(\w[49][19] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][1]$_SDFFCE_PN0P_  (.D(_02101_),
    .DE(_00074_),
    .Q(\w[49][1] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][20]$_SDFFCE_PN0P_  (.D(_02102_),
    .DE(_00074_),
    .Q(\w[49][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][21]$_SDFFCE_PN0P_  (.D(_02103_),
    .DE(_00074_),
    .Q(\w[49][21] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][22]$_SDFFCE_PN0P_  (.D(_02104_),
    .DE(_00074_),
    .Q(\w[49][22] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][23]$_SDFFCE_PN0P_  (.D(_02105_),
    .DE(_00074_),
    .Q(\w[49][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][24]$_SDFFCE_PN0P_  (.D(_02106_),
    .DE(_00074_),
    .Q(\w[49][24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][25]$_SDFFCE_PN0P_  (.D(_02107_),
    .DE(_00074_),
    .Q(\w[49][25] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][26]$_SDFFCE_PN0P_  (.D(_02108_),
    .DE(_00074_),
    .Q(\w[49][26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][27]$_SDFFCE_PN0P_  (.D(_02109_),
    .DE(_00074_),
    .Q(\w[49][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][28]$_SDFFCE_PN0P_  (.D(_02110_),
    .DE(_00074_),
    .Q(\w[49][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][29]$_SDFFCE_PN0P_  (.D(_02111_),
    .DE(_00074_),
    .Q(\w[49][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][2]$_SDFFCE_PN0P_  (.D(_02112_),
    .DE(_00074_),
    .Q(\w[49][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][30]$_SDFFCE_PN0P_  (.D(_02113_),
    .DE(_00074_),
    .Q(\w[49][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][31]$_SDFFCE_PN0P_  (.D(_02114_),
    .DE(_00074_),
    .Q(\w[49][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][3]$_SDFFCE_PN0P_  (.D(_02115_),
    .DE(_00074_),
    .Q(\w[49][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][4]$_SDFFCE_PN0P_  (.D(_02116_),
    .DE(_00074_),
    .Q(\w[49][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][5]$_SDFFCE_PN0P_  (.D(_02117_),
    .DE(_00074_),
    .Q(\w[49][5] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][6]$_SDFFCE_PN0P_  (.D(_02118_),
    .DE(_00074_),
    .Q(\w[49][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][7]$_SDFFCE_PN0P_  (.D(_02119_),
    .DE(_00074_),
    .Q(\w[49][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][8]$_SDFFCE_PN0P_  (.D(_02120_),
    .DE(_00074_),
    .Q(\w[49][8] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][9]$_SDFFCE_PN0P_  (.D(_02121_),
    .DE(_00074_),
    .Q(\w[49][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][0]$_DFFE_PP_  (.D(_00449_),
    .DE(_00105_),
    .Q(\w[4][0] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][10]$_DFFE_PP_  (.D(_00450_),
    .DE(_00105_),
    .Q(\w[4][10] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][11]$_DFFE_PP_  (.D(_00451_),
    .DE(_00105_),
    .Q(\w[4][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][12]$_DFFE_PP_  (.D(_00452_),
    .DE(_00105_),
    .Q(\w[4][12] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][13]$_DFFE_PP_  (.D(_00453_),
    .DE(_00105_),
    .Q(\w[4][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][14]$_DFFE_PP_  (.D(_00454_),
    .DE(_00105_),
    .Q(\w[4][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][15]$_DFFE_PP_  (.D(_00455_),
    .DE(_00105_),
    .Q(\w[4][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][16]$_DFFE_PP_  (.D(_00456_),
    .DE(_00105_),
    .Q(\w[4][16] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][17]$_DFFE_PP_  (.D(_00457_),
    .DE(_00105_),
    .Q(\w[4][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][18]$_DFFE_PP_  (.D(_00458_),
    .DE(_00105_),
    .Q(\w[4][18] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][19]$_DFFE_PP_  (.D(_00459_),
    .DE(_00105_),
    .Q(\w[4][19] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][1]$_DFFE_PP_  (.D(_00460_),
    .DE(_00105_),
    .Q(\w[4][1] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][20]$_DFFE_PP_  (.D(_00461_),
    .DE(_00105_),
    .Q(\w[4][20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][21]$_DFFE_PP_  (.D(_00462_),
    .DE(_00105_),
    .Q(\w[4][21] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][22]$_DFFE_PP_  (.D(_00463_),
    .DE(_00105_),
    .Q(\w[4][22] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][23]$_DFFE_PP_  (.D(_00464_),
    .DE(_00105_),
    .Q(\w[4][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][24]$_DFFE_PP_  (.D(_00465_),
    .DE(_00105_),
    .Q(\w[4][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][25]$_DFFE_PP_  (.D(_00466_),
    .DE(_00105_),
    .Q(\w[4][25] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][26]$_DFFE_PP_  (.D(_00467_),
    .DE(_00105_),
    .Q(\w[4][26] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][27]$_DFFE_PP_  (.D(_00468_),
    .DE(_00105_),
    .Q(\w[4][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][28]$_DFFE_PP_  (.D(_00469_),
    .DE(_00105_),
    .Q(\w[4][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][29]$_DFFE_PP_  (.D(_00470_),
    .DE(_00105_),
    .Q(\w[4][29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][2]$_DFFE_PP_  (.D(_00471_),
    .DE(_00105_),
    .Q(\w[4][2] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][30]$_DFFE_PP_  (.D(_00472_),
    .DE(_00105_),
    .Q(\w[4][30] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][31]$_DFFE_PP_  (.D(_00473_),
    .DE(_00105_),
    .Q(\w[4][31] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][3]$_DFFE_PP_  (.D(_00474_),
    .DE(_00105_),
    .Q(\w[4][3] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][4]$_DFFE_PP_  (.D(_00475_),
    .DE(_00105_),
    .Q(\w[4][4] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][5]$_DFFE_PP_  (.D(_00476_),
    .DE(_00105_),
    .Q(\w[4][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][6]$_DFFE_PP_  (.D(_00477_),
    .DE(_00105_),
    .Q(\w[4][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][7]$_DFFE_PP_  (.D(_00478_),
    .DE(_00105_),
    .Q(\w[4][7] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][8]$_DFFE_PP_  (.D(_00479_),
    .DE(_00105_),
    .Q(\w[4][8] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][9]$_DFFE_PP_  (.D(_00480_),
    .DE(_00105_),
    .Q(\w[4][9] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][0]$_SDFFCE_PN0P_  (.D(_02122_),
    .DE(_00104_),
    .Q(\w[50][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][10]$_SDFFCE_PN0P_  (.D(_02123_),
    .DE(_00104_),
    .Q(\w[50][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][11]$_SDFFCE_PN0P_  (.D(_02124_),
    .DE(_00104_),
    .Q(\w[50][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][12]$_SDFFCE_PN0P_  (.D(_02125_),
    .DE(_00104_),
    .Q(\w[50][12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][13]$_SDFFCE_PN0P_  (.D(_02126_),
    .DE(_00104_),
    .Q(\w[50][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][14]$_SDFFCE_PN0P_  (.D(_02127_),
    .DE(_00104_),
    .Q(\w[50][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][15]$_SDFFCE_PN0P_  (.D(_02128_),
    .DE(_00104_),
    .Q(\w[50][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][16]$_SDFFCE_PN0P_  (.D(_02129_),
    .DE(_00104_),
    .Q(\w[50][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][17]$_SDFFCE_PN0P_  (.D(_02130_),
    .DE(_00104_),
    .Q(\w[50][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][18]$_SDFFCE_PN0P_  (.D(_02131_),
    .DE(_00104_),
    .Q(\w[50][18] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][19]$_SDFFCE_PN0P_  (.D(_02132_),
    .DE(_00104_),
    .Q(\w[50][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][1]$_SDFFCE_PN0P_  (.D(_02133_),
    .DE(_00104_),
    .Q(\w[50][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][20]$_SDFFCE_PN0P_  (.D(_02134_),
    .DE(_00104_),
    .Q(\w[50][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][21]$_SDFFCE_PN0P_  (.D(_02135_),
    .DE(_00104_),
    .Q(\w[50][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][22]$_SDFFCE_PN0P_  (.D(_02136_),
    .DE(_00104_),
    .Q(\w[50][22] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][23]$_SDFFCE_PN0P_  (.D(_02137_),
    .DE(_00104_),
    .Q(\w[50][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][24]$_SDFFCE_PN0P_  (.D(_02138_),
    .DE(_00104_),
    .Q(\w[50][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][25]$_SDFFCE_PN0P_  (.D(_02139_),
    .DE(_00104_),
    .Q(\w[50][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][26]$_SDFFCE_PN0P_  (.D(_02140_),
    .DE(_00104_),
    .Q(\w[50][26] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][27]$_SDFFCE_PN0P_  (.D(_02141_),
    .DE(_00104_),
    .Q(\w[50][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][28]$_SDFFCE_PN0P_  (.D(_02142_),
    .DE(_00104_),
    .Q(\w[50][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][29]$_SDFFCE_PN0P_  (.D(_02143_),
    .DE(_00104_),
    .Q(\w[50][29] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][2]$_SDFFCE_PN0P_  (.D(_02144_),
    .DE(_00104_),
    .Q(\w[50][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][30]$_SDFFCE_PN0P_  (.D(_02145_),
    .DE(_00104_),
    .Q(\w[50][30] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][31]$_SDFFCE_PN0P_  (.D(_02146_),
    .DE(_00104_),
    .Q(\w[50][31] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][3]$_SDFFCE_PN0P_  (.D(_02147_),
    .DE(_00104_),
    .Q(\w[50][3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][4]$_SDFFCE_PN0P_  (.D(_02148_),
    .DE(_00104_),
    .Q(\w[50][4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][5]$_SDFFCE_PN0P_  (.D(_02149_),
    .DE(_00104_),
    .Q(\w[50][5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][6]$_SDFFCE_PN0P_  (.D(_02150_),
    .DE(_00104_),
    .Q(\w[50][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][7]$_SDFFCE_PN0P_  (.D(_02151_),
    .DE(_00104_),
    .Q(\w[50][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][8]$_SDFFCE_PN0P_  (.D(_02152_),
    .DE(_00104_),
    .Q(\w[50][8] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][9]$_SDFFCE_PN0P_  (.D(_02153_),
    .DE(_00104_),
    .Q(\w[50][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][0]$_SDFFCE_PN0P_  (.D(_02154_),
    .DE(_00073_),
    .Q(\w[51][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][10]$_SDFFCE_PN0P_  (.D(_02155_),
    .DE(_00073_),
    .Q(\w[51][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][11]$_SDFFCE_PN0P_  (.D(_02156_),
    .DE(_00073_),
    .Q(\w[51][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][12]$_SDFFCE_PN0P_  (.D(_02157_),
    .DE(_00073_),
    .Q(\w[51][12] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][13]$_SDFFCE_PN0P_  (.D(_02158_),
    .DE(_00073_),
    .Q(\w[51][13] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][14]$_SDFFCE_PN0P_  (.D(_02159_),
    .DE(_00073_),
    .Q(\w[51][14] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][15]$_SDFFCE_PN0P_  (.D(_02160_),
    .DE(_00073_),
    .Q(\w[51][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][16]$_SDFFCE_PN0P_  (.D(_02161_),
    .DE(_00073_),
    .Q(\w[51][16] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][17]$_SDFFCE_PN0P_  (.D(_02162_),
    .DE(_00073_),
    .Q(\w[51][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][18]$_SDFFCE_PN0P_  (.D(_02163_),
    .DE(_00073_),
    .Q(\w[51][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][19]$_SDFFCE_PN0P_  (.D(_02164_),
    .DE(_00073_),
    .Q(\w[51][19] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][1]$_SDFFCE_PN0P_  (.D(_02165_),
    .DE(_00073_),
    .Q(\w[51][1] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][20]$_SDFFCE_PN0P_  (.D(_02166_),
    .DE(_00073_),
    .Q(\w[51][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][21]$_SDFFCE_PN0P_  (.D(_02167_),
    .DE(_00073_),
    .Q(\w[51][21] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][22]$_SDFFCE_PN0P_  (.D(_02168_),
    .DE(_00073_),
    .Q(\w[51][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][23]$_SDFFCE_PN0P_  (.D(_02169_),
    .DE(_00073_),
    .Q(\w[51][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][24]$_SDFFCE_PN0P_  (.D(_02170_),
    .DE(_00073_),
    .Q(\w[51][24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][25]$_SDFFCE_PN0P_  (.D(_02171_),
    .DE(_00073_),
    .Q(\w[51][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][26]$_SDFFCE_PN0P_  (.D(_02172_),
    .DE(_00073_),
    .Q(\w[51][26] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][27]$_SDFFCE_PN0P_  (.D(_02173_),
    .DE(_00073_),
    .Q(\w[51][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][28]$_SDFFCE_PN0P_  (.D(_02174_),
    .DE(_00073_),
    .Q(\w[51][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][29]$_SDFFCE_PN0P_  (.D(_02175_),
    .DE(_00073_),
    .Q(\w[51][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][2]$_SDFFCE_PN0P_  (.D(_02176_),
    .DE(_00073_),
    .Q(\w[51][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][30]$_SDFFCE_PN0P_  (.D(_02177_),
    .DE(_00073_),
    .Q(\w[51][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][31]$_SDFFCE_PN0P_  (.D(_02178_),
    .DE(_00073_),
    .Q(\w[51][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][3]$_SDFFCE_PN0P_  (.D(_02179_),
    .DE(_00073_),
    .Q(\w[51][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][4]$_SDFFCE_PN0P_  (.D(_02180_),
    .DE(_00073_),
    .Q(\w[51][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][5]$_SDFFCE_PN0P_  (.D(_02181_),
    .DE(_00073_),
    .Q(\w[51][5] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][6]$_SDFFCE_PN0P_  (.D(_02182_),
    .DE(_00073_),
    .Q(\w[51][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][7]$_SDFFCE_PN0P_  (.D(_02183_),
    .DE(_00073_),
    .Q(\w[51][7] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][8]$_SDFFCE_PN0P_  (.D(_02184_),
    .DE(_00073_),
    .Q(\w[51][8] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][9]$_SDFFCE_PN0P_  (.D(_02185_),
    .DE(_00073_),
    .Q(\w[51][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][0]$_SDFFCE_PN0P_  (.D(_02186_),
    .DE(_00103_),
    .Q(\w[52][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][10]$_SDFFCE_PN0P_  (.D(_02187_),
    .DE(_00103_),
    .Q(\w[52][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][11]$_SDFFCE_PN0P_  (.D(_02188_),
    .DE(_00103_),
    .Q(\w[52][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][12]$_SDFFCE_PN0P_  (.D(_02189_),
    .DE(_00103_),
    .Q(\w[52][12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][13]$_SDFFCE_PN0P_  (.D(_02190_),
    .DE(_00103_),
    .Q(\w[52][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][14]$_SDFFCE_PN0P_  (.D(_02191_),
    .DE(_00103_),
    .Q(\w[52][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][15]$_SDFFCE_PN0P_  (.D(_02192_),
    .DE(_00103_),
    .Q(\w[52][15] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][16]$_SDFFCE_PN0P_  (.D(_02193_),
    .DE(_00103_),
    .Q(\w[52][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][17]$_SDFFCE_PN0P_  (.D(_02194_),
    .DE(_00103_),
    .Q(\w[52][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][18]$_SDFFCE_PN0P_  (.D(_02195_),
    .DE(_00103_),
    .Q(\w[52][18] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][19]$_SDFFCE_PN0P_  (.D(_02196_),
    .DE(_00103_),
    .Q(\w[52][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][1]$_SDFFCE_PN0P_  (.D(_02197_),
    .DE(_00103_),
    .Q(\w[52][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][20]$_SDFFCE_PN0P_  (.D(_02198_),
    .DE(_00103_),
    .Q(\w[52][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][21]$_SDFFCE_PN0P_  (.D(_02199_),
    .DE(_00103_),
    .Q(\w[52][21] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][22]$_SDFFCE_PN0P_  (.D(_02200_),
    .DE(_00103_),
    .Q(\w[52][22] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][23]$_SDFFCE_PN0P_  (.D(_02201_),
    .DE(_00103_),
    .Q(\w[52][23] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][24]$_SDFFCE_PN0P_  (.D(_02202_),
    .DE(_00103_),
    .Q(\w[52][24] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][25]$_SDFFCE_PN0P_  (.D(_02203_),
    .DE(_00103_),
    .Q(\w[52][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][26]$_SDFFCE_PN0P_  (.D(_02204_),
    .DE(_00103_),
    .Q(\w[52][26] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][27]$_SDFFCE_PN0P_  (.D(_02205_),
    .DE(_00103_),
    .Q(\w[52][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][28]$_SDFFCE_PN0P_  (.D(_02206_),
    .DE(_00103_),
    .Q(\w[52][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][29]$_SDFFCE_PN0P_  (.D(_02207_),
    .DE(_00103_),
    .Q(\w[52][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][2]$_SDFFCE_PN0P_  (.D(_02208_),
    .DE(_00103_),
    .Q(\w[52][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][30]$_SDFFCE_PN0P_  (.D(_02209_),
    .DE(_00103_),
    .Q(\w[52][30] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][31]$_SDFFCE_PN0P_  (.D(_02210_),
    .DE(_00103_),
    .Q(\w[52][31] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][3]$_SDFFCE_PN0P_  (.D(_02211_),
    .DE(_00103_),
    .Q(\w[52][3] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][4]$_SDFFCE_PN0P_  (.D(_02212_),
    .DE(_00103_),
    .Q(\w[52][4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][5]$_SDFFCE_PN0P_  (.D(_02213_),
    .DE(_00103_),
    .Q(\w[52][5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][6]$_SDFFCE_PN0P_  (.D(_02214_),
    .DE(_00103_),
    .Q(\w[52][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][7]$_SDFFCE_PN0P_  (.D(_02215_),
    .DE(_00103_),
    .Q(\w[52][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][8]$_SDFFCE_PN0P_  (.D(_02216_),
    .DE(_00103_),
    .Q(\w[52][8] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][9]$_SDFFCE_PN0P_  (.D(_02217_),
    .DE(_00103_),
    .Q(\w[52][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][0]$_SDFFCE_PN0P_  (.D(_02218_),
    .DE(_00072_),
    .Q(\w[53][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][10]$_SDFFCE_PN0P_  (.D(_02219_),
    .DE(_00072_),
    .Q(\w[53][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][11]$_SDFFCE_PN0P_  (.D(_02220_),
    .DE(_00072_),
    .Q(\w[53][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][12]$_SDFFCE_PN0P_  (.D(_02221_),
    .DE(_00072_),
    .Q(\w[53][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][13]$_SDFFCE_PN0P_  (.D(_02222_),
    .DE(_00072_),
    .Q(\w[53][13] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][14]$_SDFFCE_PN0P_  (.D(_02223_),
    .DE(_00072_),
    .Q(\w[53][14] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][15]$_SDFFCE_PN0P_  (.D(_02224_),
    .DE(_00072_),
    .Q(\w[53][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][16]$_SDFFCE_PN0P_  (.D(_02225_),
    .DE(_00072_),
    .Q(\w[53][16] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][17]$_SDFFCE_PN0P_  (.D(_02226_),
    .DE(_00072_),
    .Q(\w[53][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][18]$_SDFFCE_PN0P_  (.D(_02227_),
    .DE(_00072_),
    .Q(\w[53][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][19]$_SDFFCE_PN0P_  (.D(_02228_),
    .DE(_00072_),
    .Q(\w[53][19] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][1]$_SDFFCE_PN0P_  (.D(_02229_),
    .DE(_00072_),
    .Q(\w[53][1] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][20]$_SDFFCE_PN0P_  (.D(_02230_),
    .DE(_00072_),
    .Q(\w[53][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][21]$_SDFFCE_PN0P_  (.D(_02231_),
    .DE(_00072_),
    .Q(\w[53][21] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][22]$_SDFFCE_PN0P_  (.D(_02232_),
    .DE(_00072_),
    .Q(\w[53][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][23]$_SDFFCE_PN0P_  (.D(_02233_),
    .DE(_00072_),
    .Q(\w[53][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][24]$_SDFFCE_PN0P_  (.D(_02234_),
    .DE(_00072_),
    .Q(\w[53][24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][25]$_SDFFCE_PN0P_  (.D(_02235_),
    .DE(_00072_),
    .Q(\w[53][25] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][26]$_SDFFCE_PN0P_  (.D(_02236_),
    .DE(_00072_),
    .Q(\w[53][26] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][27]$_SDFFCE_PN0P_  (.D(_02237_),
    .DE(_00072_),
    .Q(\w[53][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][28]$_SDFFCE_PN0P_  (.D(_02238_),
    .DE(_00072_),
    .Q(\w[53][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][29]$_SDFFCE_PN0P_  (.D(_02239_),
    .DE(_00072_),
    .Q(\w[53][29] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][2]$_SDFFCE_PN0P_  (.D(_02240_),
    .DE(_00072_),
    .Q(\w[53][2] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][30]$_SDFFCE_PN0P_  (.D(_02241_),
    .DE(_00072_),
    .Q(\w[53][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][31]$_SDFFCE_PN0P_  (.D(_02242_),
    .DE(_00072_),
    .Q(\w[53][31] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][3]$_SDFFCE_PN0P_  (.D(_02243_),
    .DE(_00072_),
    .Q(\w[53][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][4]$_SDFFCE_PN0P_  (.D(_02244_),
    .DE(_00072_),
    .Q(\w[53][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][5]$_SDFFCE_PN0P_  (.D(_02245_),
    .DE(_00072_),
    .Q(\w[53][5] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][6]$_SDFFCE_PN0P_  (.D(_02246_),
    .DE(_00072_),
    .Q(\w[53][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][7]$_SDFFCE_PN0P_  (.D(_02247_),
    .DE(_00072_),
    .Q(\w[53][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][8]$_SDFFCE_PN0P_  (.D(_02248_),
    .DE(_00072_),
    .Q(\w[53][8] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][9]$_SDFFCE_PN0P_  (.D(_02249_),
    .DE(_00072_),
    .Q(\w[53][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][0]$_SDFFCE_PN0P_  (.D(_02250_),
    .DE(_00102_),
    .Q(\w[54][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][10]$_SDFFCE_PN0P_  (.D(_02251_),
    .DE(_00102_),
    .Q(\w[54][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][11]$_SDFFCE_PN0P_  (.D(_02252_),
    .DE(_00102_),
    .Q(\w[54][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][12]$_SDFFCE_PN0P_  (.D(_02253_),
    .DE(_00102_),
    .Q(\w[54][12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][13]$_SDFFCE_PN0P_  (.D(_02254_),
    .DE(_00102_),
    .Q(\w[54][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][14]$_SDFFCE_PN0P_  (.D(_02255_),
    .DE(_00102_),
    .Q(\w[54][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][15]$_SDFFCE_PN0P_  (.D(_02256_),
    .DE(_00102_),
    .Q(\w[54][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][16]$_SDFFCE_PN0P_  (.D(_02257_),
    .DE(_00102_),
    .Q(\w[54][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][17]$_SDFFCE_PN0P_  (.D(_02258_),
    .DE(_00102_),
    .Q(\w[54][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][18]$_SDFFCE_PN0P_  (.D(_02259_),
    .DE(_00102_),
    .Q(\w[54][18] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][19]$_SDFFCE_PN0P_  (.D(_02260_),
    .DE(_00102_),
    .Q(\w[54][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][1]$_SDFFCE_PN0P_  (.D(_02261_),
    .DE(_00102_),
    .Q(\w[54][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][20]$_SDFFCE_PN0P_  (.D(_02262_),
    .DE(_00102_),
    .Q(\w[54][20] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][21]$_SDFFCE_PN0P_  (.D(_02263_),
    .DE(_00102_),
    .Q(\w[54][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][22]$_SDFFCE_PN0P_  (.D(_02264_),
    .DE(_00102_),
    .Q(\w[54][22] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][23]$_SDFFCE_PN0P_  (.D(_02265_),
    .DE(_00102_),
    .Q(\w[54][23] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][24]$_SDFFCE_PN0P_  (.D(_02266_),
    .DE(_00102_),
    .Q(\w[54][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][25]$_SDFFCE_PN0P_  (.D(_02267_),
    .DE(_00102_),
    .Q(\w[54][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][26]$_SDFFCE_PN0P_  (.D(_02268_),
    .DE(_00102_),
    .Q(\w[54][26] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][27]$_SDFFCE_PN0P_  (.D(_02269_),
    .DE(_00102_),
    .Q(\w[54][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][28]$_SDFFCE_PN0P_  (.D(_02270_),
    .DE(_00102_),
    .Q(\w[54][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][29]$_SDFFCE_PN0P_  (.D(_02271_),
    .DE(_00102_),
    .Q(\w[54][29] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][2]$_SDFFCE_PN0P_  (.D(_02272_),
    .DE(_00102_),
    .Q(\w[54][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][30]$_SDFFCE_PN0P_  (.D(_02273_),
    .DE(_00102_),
    .Q(\w[54][30] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][31]$_SDFFCE_PN0P_  (.D(_02274_),
    .DE(_00102_),
    .Q(\w[54][31] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][3]$_SDFFCE_PN0P_  (.D(_02275_),
    .DE(_00102_),
    .Q(\w[54][3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][4]$_SDFFCE_PN0P_  (.D(_02276_),
    .DE(_00102_),
    .Q(\w[54][4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][5]$_SDFFCE_PN0P_  (.D(_02277_),
    .DE(_00102_),
    .Q(\w[54][5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][6]$_SDFFCE_PN0P_  (.D(_02278_),
    .DE(_00102_),
    .Q(\w[54][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][7]$_SDFFCE_PN0P_  (.D(_02279_),
    .DE(_00102_),
    .Q(\w[54][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][8]$_SDFFCE_PN0P_  (.D(_02280_),
    .DE(_00102_),
    .Q(\w[54][8] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][9]$_SDFFCE_PN0P_  (.D(_02281_),
    .DE(_00102_),
    .Q(\w[54][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][0]$_SDFFCE_PN0P_  (.D(_02282_),
    .DE(net302),
    .Q(\w[55][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][10]$_SDFFCE_PN0P_  (.D(_02283_),
    .DE(_00071_),
    .Q(\w[55][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][11]$_SDFFCE_PN0P_  (.D(_02284_),
    .DE(_00071_),
    .Q(\w[55][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][12]$_SDFFCE_PN0P_  (.D(_02285_),
    .DE(net301),
    .Q(\w[55][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][13]$_SDFFCE_PN0P_  (.D(_02286_),
    .DE(_00071_),
    .Q(\w[55][13] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][14]$_SDFFCE_PN0P_  (.D(_02287_),
    .DE(net301),
    .Q(\w[55][14] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][15]$_SDFFCE_PN0P_  (.D(_02288_),
    .DE(net302),
    .Q(\w[55][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][16]$_SDFFCE_PN0P_  (.D(_02289_),
    .DE(net301),
    .Q(\w[55][16] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][17]$_SDFFCE_PN0P_  (.D(_02290_),
    .DE(net301),
    .Q(\w[55][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][18]$_SDFFCE_PN0P_  (.D(_02291_),
    .DE(net301),
    .Q(\w[55][18] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][19]$_SDFFCE_PN0P_  (.D(_02292_),
    .DE(net301),
    .Q(\w[55][19] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][1]$_SDFFCE_PN0P_  (.D(_02293_),
    .DE(net302),
    .Q(\w[55][1] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][20]$_SDFFCE_PN0P_  (.D(_02294_),
    .DE(_00071_),
    .Q(\w[55][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][21]$_SDFFCE_PN0P_  (.D(_02295_),
    .DE(net301),
    .Q(\w[55][21] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][22]$_SDFFCE_PN0P_  (.D(_02296_),
    .DE(net301),
    .Q(\w[55][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][23]$_SDFFCE_PN0P_  (.D(_02297_),
    .DE(net301),
    .Q(\w[55][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][24]$_SDFFCE_PN0P_  (.D(_02298_),
    .DE(net302),
    .Q(\w[55][24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][25]$_SDFFCE_PN0P_  (.D(_02299_),
    .DE(net301),
    .Q(\w[55][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][26]$_SDFFCE_PN0P_  (.D(_02300_),
    .DE(net302),
    .Q(\w[55][26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][27]$_SDFFCE_PN0P_  (.D(_02301_),
    .DE(net301),
    .Q(\w[55][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][28]$_SDFFCE_PN0P_  (.D(_02302_),
    .DE(net302),
    .Q(\w[55][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][29]$_SDFFCE_PN0P_  (.D(_02303_),
    .DE(net302),
    .Q(\w[55][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][2]$_SDFFCE_PN0P_  (.D(_02304_),
    .DE(net301),
    .Q(\w[55][2] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][30]$_SDFFCE_PN0P_  (.D(_02305_),
    .DE(_00071_),
    .Q(\w[55][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][31]$_SDFFCE_PN0P_  (.D(_02306_),
    .DE(net302),
    .Q(\w[55][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][3]$_SDFFCE_PN0P_  (.D(_02307_),
    .DE(net302),
    .Q(\w[55][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][4]$_SDFFCE_PN0P_  (.D(_02308_),
    .DE(net301),
    .Q(\w[55][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][5]$_SDFFCE_PN0P_  (.D(_02309_),
    .DE(net302),
    .Q(\w[55][5] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][6]$_SDFFCE_PN0P_  (.D(_02310_),
    .DE(_00071_),
    .Q(\w[55][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][7]$_SDFFCE_PN0P_  (.D(_02311_),
    .DE(_00071_),
    .Q(\w[55][7] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][8]$_SDFFCE_PN0P_  (.D(_02312_),
    .DE(net301),
    .Q(\w[55][8] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][9]$_SDFFCE_PN0P_  (.D(_02313_),
    .DE(_00071_),
    .Q(\w[55][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][0]$_SDFFCE_PN0P_  (.D(_02314_),
    .DE(_00101_),
    .Q(\w[56][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][10]$_SDFFCE_PN0P_  (.D(_02315_),
    .DE(_00101_),
    .Q(\w[56][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][11]$_SDFFCE_PN0P_  (.D(_02316_),
    .DE(_00101_),
    .Q(\w[56][11] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][12]$_SDFFCE_PN0P_  (.D(_02317_),
    .DE(_00101_),
    .Q(\w[56][12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][13]$_SDFFCE_PN0P_  (.D(_02318_),
    .DE(_00101_),
    .Q(\w[56][13] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][14]$_SDFFCE_PN0P_  (.D(_02319_),
    .DE(_00101_),
    .Q(\w[56][14] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][15]$_SDFFCE_PN0P_  (.D(_02320_),
    .DE(_00101_),
    .Q(\w[56][15] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][16]$_SDFFCE_PN0P_  (.D(_02321_),
    .DE(_00101_),
    .Q(\w[56][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][17]$_SDFFCE_PN0P_  (.D(_02322_),
    .DE(_00101_),
    .Q(\w[56][17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][18]$_SDFFCE_PN0P_  (.D(_02323_),
    .DE(_00101_),
    .Q(\w[56][18] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][19]$_SDFFCE_PN0P_  (.D(_02324_),
    .DE(_00101_),
    .Q(\w[56][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][1]$_SDFFCE_PN0P_  (.D(_02325_),
    .DE(_00101_),
    .Q(\w[56][1] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][20]$_SDFFCE_PN0P_  (.D(_02326_),
    .DE(_00101_),
    .Q(\w[56][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][21]$_SDFFCE_PN0P_  (.D(_02327_),
    .DE(_00101_),
    .Q(\w[56][21] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][22]$_SDFFCE_PN0P_  (.D(_02328_),
    .DE(_00101_),
    .Q(\w[56][22] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][23]$_SDFFCE_PN0P_  (.D(_02329_),
    .DE(_00101_),
    .Q(\w[56][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][24]$_SDFFCE_PN0P_  (.D(_02330_),
    .DE(_00101_),
    .Q(\w[56][24] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][25]$_SDFFCE_PN0P_  (.D(_02331_),
    .DE(_00101_),
    .Q(\w[56][25] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][26]$_SDFFCE_PN0P_  (.D(_02332_),
    .DE(_00101_),
    .Q(\w[56][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][27]$_SDFFCE_PN0P_  (.D(_02333_),
    .DE(_00101_),
    .Q(\w[56][27] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][28]$_SDFFCE_PN0P_  (.D(_02334_),
    .DE(_00101_),
    .Q(\w[56][28] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][29]$_SDFFCE_PN0P_  (.D(_02335_),
    .DE(_00101_),
    .Q(\w[56][29] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][2]$_SDFFCE_PN0P_  (.D(_02336_),
    .DE(_00101_),
    .Q(\w[56][2] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][30]$_SDFFCE_PN0P_  (.D(_02337_),
    .DE(_00101_),
    .Q(\w[56][30] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][31]$_SDFFCE_PN0P_  (.D(_02338_),
    .DE(_00101_),
    .Q(\w[56][31] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][3]$_SDFFCE_PN0P_  (.D(_02339_),
    .DE(_00101_),
    .Q(\w[56][3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][4]$_SDFFCE_PN0P_  (.D(_02340_),
    .DE(_00101_),
    .Q(\w[56][4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][5]$_SDFFCE_PN0P_  (.D(_02341_),
    .DE(_00101_),
    .Q(\w[56][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][6]$_SDFFCE_PN0P_  (.D(_02342_),
    .DE(_00101_),
    .Q(\w[56][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][7]$_SDFFCE_PN0P_  (.D(_02343_),
    .DE(_00101_),
    .Q(\w[56][7] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][8]$_SDFFCE_PN0P_  (.D(_02344_),
    .DE(_00101_),
    .Q(\w[56][8] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][9]$_SDFFCE_PN0P_  (.D(_02345_),
    .DE(_00101_),
    .Q(\w[56][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][0]$_SDFFCE_PN0P_  (.D(_02346_),
    .DE(_00070_),
    .Q(\w[57][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][10]$_SDFFCE_PN0P_  (.D(_02347_),
    .DE(_00070_),
    .Q(\w[57][10] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][11]$_SDFFCE_PN0P_  (.D(_02348_),
    .DE(_00070_),
    .Q(\w[57][11] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][12]$_SDFFCE_PN0P_  (.D(_02349_),
    .DE(_00070_),
    .Q(\w[57][12] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][13]$_SDFFCE_PN0P_  (.D(_02350_),
    .DE(_00070_),
    .Q(\w[57][13] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][14]$_SDFFCE_PN0P_  (.D(_02351_),
    .DE(_00070_),
    .Q(\w[57][14] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][15]$_SDFFCE_PN0P_  (.D(_02352_),
    .DE(_00070_),
    .Q(\w[57][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][16]$_SDFFCE_PN0P_  (.D(_02353_),
    .DE(_00070_),
    .Q(\w[57][16] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][17]$_SDFFCE_PN0P_  (.D(_02354_),
    .DE(_00070_),
    .Q(\w[57][17] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][18]$_SDFFCE_PN0P_  (.D(_02355_),
    .DE(_00070_),
    .Q(\w[57][18] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][19]$_SDFFCE_PN0P_  (.D(_02356_),
    .DE(_00070_),
    .Q(\w[57][19] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][1]$_SDFFCE_PN0P_  (.D(_02357_),
    .DE(_00070_),
    .Q(\w[57][1] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][20]$_SDFFCE_PN0P_  (.D(_02358_),
    .DE(_00070_),
    .Q(\w[57][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][21]$_SDFFCE_PN0P_  (.D(_02359_),
    .DE(_00070_),
    .Q(\w[57][21] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][22]$_SDFFCE_PN0P_  (.D(_02360_),
    .DE(_00070_),
    .Q(\w[57][22] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][23]$_SDFFCE_PN0P_  (.D(_02361_),
    .DE(_00070_),
    .Q(\w[57][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][24]$_SDFFCE_PN0P_  (.D(_02362_),
    .DE(_00070_),
    .Q(\w[57][24] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][25]$_SDFFCE_PN0P_  (.D(_02363_),
    .DE(_00070_),
    .Q(\w[57][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][26]$_SDFFCE_PN0P_  (.D(_02364_),
    .DE(_00070_),
    .Q(\w[57][26] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][27]$_SDFFCE_PN0P_  (.D(_02365_),
    .DE(_00070_),
    .Q(\w[57][27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][28]$_SDFFCE_PN0P_  (.D(_02366_),
    .DE(_00070_),
    .Q(\w[57][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][29]$_SDFFCE_PN0P_  (.D(_02367_),
    .DE(_00070_),
    .Q(\w[57][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][2]$_SDFFCE_PN0P_  (.D(_02368_),
    .DE(_00070_),
    .Q(\w[57][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][30]$_SDFFCE_PN0P_  (.D(_02369_),
    .DE(_00070_),
    .Q(\w[57][30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][31]$_SDFFCE_PN0P_  (.D(_02370_),
    .DE(_00070_),
    .Q(\w[57][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][3]$_SDFFCE_PN0P_  (.D(_02371_),
    .DE(_00070_),
    .Q(\w[57][3] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][4]$_SDFFCE_PN0P_  (.D(_02372_),
    .DE(_00070_),
    .Q(\w[57][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][5]$_SDFFCE_PN0P_  (.D(_02373_),
    .DE(_00070_),
    .Q(\w[57][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][6]$_SDFFCE_PN0P_  (.D(_02374_),
    .DE(_00070_),
    .Q(\w[57][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][7]$_SDFFCE_PN0P_  (.D(_02375_),
    .DE(_00070_),
    .Q(\w[57][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][8]$_SDFFCE_PN0P_  (.D(_02376_),
    .DE(_00070_),
    .Q(\w[57][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][9]$_SDFFCE_PN0P_  (.D(_02377_),
    .DE(_00070_),
    .Q(\w[57][9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][0]$_SDFFCE_PN0P_  (.D(_02378_),
    .DE(_00100_),
    .Q(\w[58][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][10]$_SDFFCE_PN0P_  (.D(_02379_),
    .DE(_00100_),
    .Q(\w[58][10] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][11]$_SDFFCE_PN0P_  (.D(_02380_),
    .DE(_00100_),
    .Q(\w[58][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][12]$_SDFFCE_PN0P_  (.D(_02381_),
    .DE(_00100_),
    .Q(\w[58][12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][13]$_SDFFCE_PN0P_  (.D(_02382_),
    .DE(_00100_),
    .Q(\w[58][13] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][14]$_SDFFCE_PN0P_  (.D(_02383_),
    .DE(_00100_),
    .Q(\w[58][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][15]$_SDFFCE_PN0P_  (.D(_02384_),
    .DE(_00100_),
    .Q(\w[58][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][16]$_SDFFCE_PN0P_  (.D(_02385_),
    .DE(_00100_),
    .Q(\w[58][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][17]$_SDFFCE_PN0P_  (.D(_02386_),
    .DE(_00100_),
    .Q(\w[58][17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][18]$_SDFFCE_PN0P_  (.D(_02387_),
    .DE(_00100_),
    .Q(\w[58][18] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][19]$_SDFFCE_PN0P_  (.D(_02388_),
    .DE(_00100_),
    .Q(\w[58][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][1]$_SDFFCE_PN0P_  (.D(_02389_),
    .DE(_00100_),
    .Q(\w[58][1] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][20]$_SDFFCE_PN0P_  (.D(_02390_),
    .DE(_00100_),
    .Q(\w[58][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][21]$_SDFFCE_PN0P_  (.D(_02391_),
    .DE(_00100_),
    .Q(\w[58][21] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][22]$_SDFFCE_PN0P_  (.D(_02392_),
    .DE(_00100_),
    .Q(\w[58][22] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][23]$_SDFFCE_PN0P_  (.D(_02393_),
    .DE(_00100_),
    .Q(\w[58][23] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][24]$_SDFFCE_PN0P_  (.D(_02394_),
    .DE(_00100_),
    .Q(\w[58][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][25]$_SDFFCE_PN0P_  (.D(_02395_),
    .DE(_00100_),
    .Q(\w[58][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][26]$_SDFFCE_PN0P_  (.D(_02396_),
    .DE(_00100_),
    .Q(\w[58][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][27]$_SDFFCE_PN0P_  (.D(_02397_),
    .DE(_00100_),
    .Q(\w[58][27] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][28]$_SDFFCE_PN0P_  (.D(_02398_),
    .DE(_00100_),
    .Q(\w[58][28] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][29]$_SDFFCE_PN0P_  (.D(_02399_),
    .DE(_00100_),
    .Q(\w[58][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][2]$_SDFFCE_PN0P_  (.D(_02400_),
    .DE(_00100_),
    .Q(\w[58][2] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][30]$_SDFFCE_PN0P_  (.D(_02401_),
    .DE(_00100_),
    .Q(\w[58][30] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][31]$_SDFFCE_PN0P_  (.D(_02402_),
    .DE(_00100_),
    .Q(\w[58][31] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][3]$_SDFFCE_PN0P_  (.D(_02403_),
    .DE(_00100_),
    .Q(\w[58][3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][4]$_SDFFCE_PN0P_  (.D(_02404_),
    .DE(_00100_),
    .Q(\w[58][4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][5]$_SDFFCE_PN0P_  (.D(_02405_),
    .DE(_00100_),
    .Q(\w[58][5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][6]$_SDFFCE_PN0P_  (.D(_02406_),
    .DE(_00100_),
    .Q(\w[58][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][7]$_SDFFCE_PN0P_  (.D(_02407_),
    .DE(_00100_),
    .Q(\w[58][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][8]$_SDFFCE_PN0P_  (.D(_02408_),
    .DE(_00100_),
    .Q(\w[58][8] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][9]$_SDFFCE_PN0P_  (.D(_02409_),
    .DE(_00100_),
    .Q(\w[58][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][0]$_SDFFCE_PN0P_  (.D(_02410_),
    .DE(_00069_),
    .Q(\w[59][0] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][10]$_SDFFCE_PN0P_  (.D(_02411_),
    .DE(_00069_),
    .Q(\w[59][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][11]$_SDFFCE_PN0P_  (.D(_02412_),
    .DE(_00069_),
    .Q(\w[59][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][12]$_SDFFCE_PN0P_  (.D(_02413_),
    .DE(_00069_),
    .Q(\w[59][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][13]$_SDFFCE_PN0P_  (.D(_02414_),
    .DE(_00069_),
    .Q(\w[59][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][14]$_SDFFCE_PN0P_  (.D(_02415_),
    .DE(_00069_),
    .Q(\w[59][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][15]$_SDFFCE_PN0P_  (.D(_02416_),
    .DE(_00069_),
    .Q(\w[59][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][16]$_SDFFCE_PN0P_  (.D(_02417_),
    .DE(_00069_),
    .Q(\w[59][16] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][17]$_SDFFCE_PN0P_  (.D(_02418_),
    .DE(_00069_),
    .Q(\w[59][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][18]$_SDFFCE_PN0P_  (.D(_02419_),
    .DE(_00069_),
    .Q(\w[59][18] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][19]$_SDFFCE_PN0P_  (.D(_02420_),
    .DE(_00069_),
    .Q(\w[59][19] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][1]$_SDFFCE_PN0P_  (.D(_02421_),
    .DE(_00069_),
    .Q(\w[59][1] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][20]$_SDFFCE_PN0P_  (.D(_02422_),
    .DE(_00069_),
    .Q(\w[59][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][21]$_SDFFCE_PN0P_  (.D(_02423_),
    .DE(_00069_),
    .Q(\w[59][21] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][22]$_SDFFCE_PN0P_  (.D(_02424_),
    .DE(_00069_),
    .Q(\w[59][22] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][23]$_SDFFCE_PN0P_  (.D(_02425_),
    .DE(_00069_),
    .Q(\w[59][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][24]$_SDFFCE_PN0P_  (.D(_02426_),
    .DE(_00069_),
    .Q(\w[59][24] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][25]$_SDFFCE_PN0P_  (.D(_02427_),
    .DE(_00069_),
    .Q(\w[59][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][26]$_SDFFCE_PN0P_  (.D(_02428_),
    .DE(_00069_),
    .Q(\w[59][26] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][27]$_SDFFCE_PN0P_  (.D(_02429_),
    .DE(_00069_),
    .Q(\w[59][27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][28]$_SDFFCE_PN0P_  (.D(_02430_),
    .DE(_00069_),
    .Q(\w[59][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][29]$_SDFFCE_PN0P_  (.D(_02431_),
    .DE(_00069_),
    .Q(\w[59][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][2]$_SDFFCE_PN0P_  (.D(_02432_),
    .DE(_00069_),
    .Q(\w[59][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][30]$_SDFFCE_PN0P_  (.D(_02433_),
    .DE(_00069_),
    .Q(\w[59][30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][31]$_SDFFCE_PN0P_  (.D(_02434_),
    .DE(_00069_),
    .Q(\w[59][31] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][3]$_SDFFCE_PN0P_  (.D(_02435_),
    .DE(_00069_),
    .Q(\w[59][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][4]$_SDFFCE_PN0P_  (.D(_02436_),
    .DE(_00069_),
    .Q(\w[59][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][5]$_SDFFCE_PN0P_  (.D(_02437_),
    .DE(_00069_),
    .Q(\w[59][5] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][6]$_SDFFCE_PN0P_  (.D(_02438_),
    .DE(_00069_),
    .Q(\w[59][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][7]$_SDFFCE_PN0P_  (.D(_02439_),
    .DE(_00069_),
    .Q(\w[59][7] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][8]$_SDFFCE_PN0P_  (.D(_02440_),
    .DE(_00069_),
    .Q(\w[59][8] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][9]$_SDFFCE_PN0P_  (.D(_02441_),
    .DE(_00069_),
    .Q(\w[59][9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][0]$_DFFE_PP_  (.D(_00481_),
    .DE(_00068_),
    .Q(\w[5][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][10]$_DFFE_PP_  (.D(_00482_),
    .DE(_00068_),
    .Q(\w[5][10] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][11]$_DFFE_PP_  (.D(_00483_),
    .DE(_00068_),
    .Q(\w[5][11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][12]$_DFFE_PP_  (.D(_00484_),
    .DE(_00068_),
    .Q(\w[5][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][13]$_DFFE_PP_  (.D(_00485_),
    .DE(_00068_),
    .Q(\w[5][13] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][14]$_DFFE_PP_  (.D(_00486_),
    .DE(_00068_),
    .Q(\w[5][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][15]$_DFFE_PP_  (.D(_00487_),
    .DE(_00068_),
    .Q(\w[5][15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][16]$_DFFE_PP_  (.D(_00488_),
    .DE(_00068_),
    .Q(\w[5][16] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][17]$_DFFE_PP_  (.D(_00489_),
    .DE(_00068_),
    .Q(\w[5][17] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][18]$_DFFE_PP_  (.D(_00490_),
    .DE(_00068_),
    .Q(\w[5][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][19]$_DFFE_PP_  (.D(_00491_),
    .DE(_00068_),
    .Q(\w[5][19] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][1]$_DFFE_PP_  (.D(_00492_),
    .DE(_00068_),
    .Q(\w[5][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][20]$_DFFE_PP_  (.D(_00493_),
    .DE(_00068_),
    .Q(\w[5][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][21]$_DFFE_PP_  (.D(_00494_),
    .DE(_00068_),
    .Q(\w[5][21] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][22]$_DFFE_PP_  (.D(_00495_),
    .DE(_00068_),
    .Q(\w[5][22] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][23]$_DFFE_PP_  (.D(_00496_),
    .DE(_00068_),
    .Q(\w[5][23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][24]$_DFFE_PP_  (.D(_00497_),
    .DE(_00068_),
    .Q(\w[5][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][25]$_DFFE_PP_  (.D(_00498_),
    .DE(_00068_),
    .Q(\w[5][25] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][26]$_DFFE_PP_  (.D(_00499_),
    .DE(_00068_),
    .Q(\w[5][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][27]$_DFFE_PP_  (.D(_00500_),
    .DE(_00068_),
    .Q(\w[5][27] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][28]$_DFFE_PP_  (.D(_00501_),
    .DE(_00068_),
    .Q(\w[5][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][29]$_DFFE_PP_  (.D(_00502_),
    .DE(_00068_),
    .Q(\w[5][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][2]$_DFFE_PP_  (.D(_00503_),
    .DE(_00068_),
    .Q(\w[5][2] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][30]$_DFFE_PP_  (.D(_00504_),
    .DE(_00068_),
    .Q(\w[5][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][31]$_DFFE_PP_  (.D(_00505_),
    .DE(_00068_),
    .Q(\w[5][31] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][3]$_DFFE_PP_  (.D(_00506_),
    .DE(_00068_),
    .Q(\w[5][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][4]$_DFFE_PP_  (.D(_00507_),
    .DE(_00068_),
    .Q(\w[5][4] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][5]$_DFFE_PP_  (.D(_00508_),
    .DE(_00068_),
    .Q(\w[5][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][6]$_DFFE_PP_  (.D(_00509_),
    .DE(_00068_),
    .Q(\w[5][6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][7]$_DFFE_PP_  (.D(_00510_),
    .DE(_00068_),
    .Q(\w[5][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][8]$_DFFE_PP_  (.D(_00511_),
    .DE(_00068_),
    .Q(\w[5][8] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][9]$_DFFE_PP_  (.D(_00512_),
    .DE(_00068_),
    .Q(\w[5][9] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][0]$_SDFFCE_PN0P_  (.D(_02442_),
    .DE(_00099_),
    .Q(\w[60][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][10]$_SDFFCE_PN0P_  (.D(_02443_),
    .DE(_00099_),
    .Q(\w[60][10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][11]$_SDFFCE_PN0P_  (.D(_02444_),
    .DE(_00099_),
    .Q(\w[60][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][12]$_SDFFCE_PN0P_  (.D(_02445_),
    .DE(_00099_),
    .Q(\w[60][12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][13]$_SDFFCE_PN0P_  (.D(_02446_),
    .DE(_00099_),
    .Q(\w[60][13] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][14]$_SDFFCE_PN0P_  (.D(_02447_),
    .DE(_00099_),
    .Q(\w[60][14] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][15]$_SDFFCE_PN0P_  (.D(_02448_),
    .DE(_00099_),
    .Q(\w[60][15] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][16]$_SDFFCE_PN0P_  (.D(_02449_),
    .DE(_00099_),
    .Q(\w[60][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][17]$_SDFFCE_PN0P_  (.D(_02450_),
    .DE(_00099_),
    .Q(\w[60][17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][18]$_SDFFCE_PN0P_  (.D(_02451_),
    .DE(_00099_),
    .Q(\w[60][18] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][19]$_SDFFCE_PN0P_  (.D(_02452_),
    .DE(_00099_),
    .Q(\w[60][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][1]$_SDFFCE_PN0P_  (.D(_02453_),
    .DE(_00099_),
    .Q(\w[60][1] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][20]$_SDFFCE_PN0P_  (.D(_02454_),
    .DE(_00099_),
    .Q(\w[60][20] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][21]$_SDFFCE_PN0P_  (.D(_02455_),
    .DE(_00099_),
    .Q(\w[60][21] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][22]$_SDFFCE_PN0P_  (.D(_02456_),
    .DE(_00099_),
    .Q(\w[60][22] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][23]$_SDFFCE_PN0P_  (.D(_02457_),
    .DE(_00099_),
    .Q(\w[60][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][24]$_SDFFCE_PN0P_  (.D(_02458_),
    .DE(_00099_),
    .Q(\w[60][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][25]$_SDFFCE_PN0P_  (.D(_02459_),
    .DE(_00099_),
    .Q(\w[60][25] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][26]$_SDFFCE_PN0P_  (.D(_02460_),
    .DE(_00099_),
    .Q(\w[60][26] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][27]$_SDFFCE_PN0P_  (.D(_02461_),
    .DE(_00099_),
    .Q(\w[60][27] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][28]$_SDFFCE_PN0P_  (.D(_02462_),
    .DE(_00099_),
    .Q(\w[60][28] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][29]$_SDFFCE_PN0P_  (.D(_02463_),
    .DE(_00099_),
    .Q(\w[60][29] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][2]$_SDFFCE_PN0P_  (.D(_02464_),
    .DE(_00099_),
    .Q(\w[60][2] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][30]$_SDFFCE_PN0P_  (.D(_02465_),
    .DE(_00099_),
    .Q(\w[60][30] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][31]$_SDFFCE_PN0P_  (.D(_02466_),
    .DE(_00099_),
    .Q(\w[60][31] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][3]$_SDFFCE_PN0P_  (.D(_02467_),
    .DE(_00099_),
    .Q(\w[60][3] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][4]$_SDFFCE_PN0P_  (.D(_02468_),
    .DE(_00099_),
    .Q(\w[60][4] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][5]$_SDFFCE_PN0P_  (.D(_02469_),
    .DE(_00099_),
    .Q(\w[60][5] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][6]$_SDFFCE_PN0P_  (.D(_02470_),
    .DE(_00099_),
    .Q(\w[60][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][7]$_SDFFCE_PN0P_  (.D(_02471_),
    .DE(_00099_),
    .Q(\w[60][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][8]$_SDFFCE_PN0P_  (.D(_02472_),
    .DE(_00099_),
    .Q(\w[60][8] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][9]$_SDFFCE_PN0P_  (.D(_02473_),
    .DE(_00099_),
    .Q(\w[60][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][0]$_SDFFCE_PN0P_  (.D(_02474_),
    .DE(_00067_),
    .Q(\w[61][0] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][10]$_SDFFCE_PN0P_  (.D(_02475_),
    .DE(_00067_),
    .Q(\w[61][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][11]$_SDFFCE_PN0P_  (.D(_02476_),
    .DE(_00067_),
    .Q(\w[61][11] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][12]$_SDFFCE_PN0P_  (.D(_02477_),
    .DE(_00067_),
    .Q(\w[61][12] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][13]$_SDFFCE_PN0P_  (.D(_02478_),
    .DE(_00067_),
    .Q(\w[61][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][14]$_SDFFCE_PN0P_  (.D(_02479_),
    .DE(_00067_),
    .Q(\w[61][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][15]$_SDFFCE_PN0P_  (.D(_02480_),
    .DE(_00067_),
    .Q(\w[61][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][16]$_SDFFCE_PN0P_  (.D(_02481_),
    .DE(_00067_),
    .Q(\w[61][16] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][17]$_SDFFCE_PN0P_  (.D(_02482_),
    .DE(_00067_),
    .Q(\w[61][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][18]$_SDFFCE_PN0P_  (.D(_02483_),
    .DE(_00067_),
    .Q(\w[61][18] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][19]$_SDFFCE_PN0P_  (.D(_02484_),
    .DE(_00067_),
    .Q(\w[61][19] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][1]$_SDFFCE_PN0P_  (.D(_02485_),
    .DE(_00067_),
    .Q(\w[61][1] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][20]$_SDFFCE_PN0P_  (.D(_02486_),
    .DE(_00067_),
    .Q(\w[61][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][21]$_SDFFCE_PN0P_  (.D(_02487_),
    .DE(_00067_),
    .Q(\w[61][21] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][22]$_SDFFCE_PN0P_  (.D(_02488_),
    .DE(_00067_),
    .Q(\w[61][22] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][23]$_SDFFCE_PN0P_  (.D(_02489_),
    .DE(_00067_),
    .Q(\w[61][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][24]$_SDFFCE_PN0P_  (.D(_02490_),
    .DE(_00067_),
    .Q(\w[61][24] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][25]$_SDFFCE_PN0P_  (.D(_02491_),
    .DE(_00067_),
    .Q(\w[61][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][26]$_SDFFCE_PN0P_  (.D(_02492_),
    .DE(_00067_),
    .Q(\w[61][26] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][27]$_SDFFCE_PN0P_  (.D(_02493_),
    .DE(_00067_),
    .Q(\w[61][27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][28]$_SDFFCE_PN0P_  (.D(_02494_),
    .DE(_00067_),
    .Q(\w[61][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][29]$_SDFFCE_PN0P_  (.D(_02495_),
    .DE(_00067_),
    .Q(\w[61][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][2]$_SDFFCE_PN0P_  (.D(_02496_),
    .DE(_00067_),
    .Q(\w[61][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][30]$_SDFFCE_PN0P_  (.D(_02497_),
    .DE(_00067_),
    .Q(\w[61][30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][31]$_SDFFCE_PN0P_  (.D(_02498_),
    .DE(_00067_),
    .Q(\w[61][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][3]$_SDFFCE_PN0P_  (.D(_02499_),
    .DE(_00067_),
    .Q(\w[61][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][4]$_SDFFCE_PN0P_  (.D(_02500_),
    .DE(_00067_),
    .Q(\w[61][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][5]$_SDFFCE_PN0P_  (.D(_02501_),
    .DE(_00067_),
    .Q(\w[61][5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][6]$_SDFFCE_PN0P_  (.D(_02502_),
    .DE(_00067_),
    .Q(\w[61][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][7]$_SDFFCE_PN0P_  (.D(_02503_),
    .DE(_00067_),
    .Q(\w[61][7] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][8]$_SDFFCE_PN0P_  (.D(_02504_),
    .DE(_00067_),
    .Q(\w[61][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][9]$_SDFFCE_PN0P_  (.D(_02505_),
    .DE(_00067_),
    .Q(\w[61][9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][0]$_SDFFCE_PN0P_  (.D(_02506_),
    .DE(_00098_),
    .Q(\w[62][0] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][10]$_SDFFCE_PN0P_  (.D(_02507_),
    .DE(_00098_),
    .Q(\w[62][10] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][11]$_SDFFCE_PN0P_  (.D(_02508_),
    .DE(_00098_),
    .Q(\w[62][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][12]$_SDFFCE_PN0P_  (.D(_02509_),
    .DE(_00098_),
    .Q(\w[62][12] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][13]$_SDFFCE_PN0P_  (.D(_02510_),
    .DE(_00098_),
    .Q(\w[62][13] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][14]$_SDFFCE_PN0P_  (.D(_02511_),
    .DE(_00098_),
    .Q(\w[62][14] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][15]$_SDFFCE_PN0P_  (.D(_02512_),
    .DE(_00098_),
    .Q(\w[62][15] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][16]$_SDFFCE_PN0P_  (.D(_02513_),
    .DE(_00098_),
    .Q(\w[62][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][17]$_SDFFCE_PN0P_  (.D(_02514_),
    .DE(_00098_),
    .Q(\w[62][17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][18]$_SDFFCE_PN0P_  (.D(_02515_),
    .DE(_00098_),
    .Q(\w[62][18] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][19]$_SDFFCE_PN0P_  (.D(_02516_),
    .DE(_00098_),
    .Q(\w[62][19] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][1]$_SDFFCE_PN0P_  (.D(_02517_),
    .DE(_00098_),
    .Q(\w[62][1] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][20]$_SDFFCE_PN0P_  (.D(_02518_),
    .DE(_00098_),
    .Q(\w[62][20] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][21]$_SDFFCE_PN0P_  (.D(_02519_),
    .DE(_00098_),
    .Q(\w[62][21] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][22]$_SDFFCE_PN0P_  (.D(_02520_),
    .DE(_00098_),
    .Q(\w[62][22] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][23]$_SDFFCE_PN0P_  (.D(_02521_),
    .DE(_00098_),
    .Q(\w[62][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][24]$_SDFFCE_PN0P_  (.D(_02522_),
    .DE(_00098_),
    .Q(\w[62][24] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][25]$_SDFFCE_PN0P_  (.D(_02523_),
    .DE(_00098_),
    .Q(\w[62][25] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][26]$_SDFFCE_PN0P_  (.D(_02524_),
    .DE(_00098_),
    .Q(\w[62][26] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][27]$_SDFFCE_PN0P_  (.D(_02525_),
    .DE(_00098_),
    .Q(\w[62][27] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][28]$_SDFFCE_PN0P_  (.D(_02526_),
    .DE(_00098_),
    .Q(\w[62][28] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][29]$_SDFFCE_PN0P_  (.D(_02527_),
    .DE(_00098_),
    .Q(\w[62][29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][2]$_SDFFCE_PN0P_  (.D(_02528_),
    .DE(_00098_),
    .Q(\w[62][2] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][30]$_SDFFCE_PN0P_  (.D(_02529_),
    .DE(_00098_),
    .Q(\w[62][30] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][31]$_SDFFCE_PN0P_  (.D(_02530_),
    .DE(_00098_),
    .Q(\w[62][31] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][3]$_SDFFCE_PN0P_  (.D(_02531_),
    .DE(_00098_),
    .Q(\w[62][3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][4]$_SDFFCE_PN0P_  (.D(_02532_),
    .DE(_00098_),
    .Q(\w[62][4] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][5]$_SDFFCE_PN0P_  (.D(_02533_),
    .DE(_00098_),
    .Q(\w[62][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][6]$_SDFFCE_PN0P_  (.D(_02534_),
    .DE(_00098_),
    .Q(\w[62][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][7]$_SDFFCE_PN0P_  (.D(_02535_),
    .DE(_00098_),
    .Q(\w[62][7] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][8]$_SDFFCE_PN0P_  (.D(_02536_),
    .DE(_00098_),
    .Q(\w[62][8] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][9]$_SDFFCE_PN0P_  (.D(_02537_),
    .DE(_00098_),
    .Q(\w[62][9] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][0]$_SDFFCE_PN0P_  (.D(_02538_),
    .DE(_00066_),
    .Q(\w[63][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][10]$_SDFFCE_PN0P_  (.D(_02539_),
    .DE(_00066_),
    .Q(\w[63][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][11]$_SDFFCE_PN0P_  (.D(_02540_),
    .DE(_00066_),
    .Q(\w[63][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][12]$_SDFFCE_PN0P_  (.D(_02541_),
    .DE(_00066_),
    .Q(\w[63][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][13]$_SDFFCE_PN0P_  (.D(_02542_),
    .DE(_00066_),
    .Q(\w[63][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][14]$_SDFFCE_PN0P_  (.D(_02543_),
    .DE(_00066_),
    .Q(\w[63][14] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][15]$_SDFFCE_PN0P_  (.D(_02544_),
    .DE(_00066_),
    .Q(\w[63][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][16]$_SDFFCE_PN0P_  (.D(_02545_),
    .DE(_00066_),
    .Q(\w[63][16] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][17]$_SDFFCE_PN0P_  (.D(_02546_),
    .DE(_00066_),
    .Q(\w[63][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][18]$_SDFFCE_PN0P_  (.D(_02547_),
    .DE(_00066_),
    .Q(\w[63][18] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][19]$_SDFFCE_PN0P_  (.D(_02548_),
    .DE(_00066_),
    .Q(\w[63][19] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][1]$_SDFFCE_PN0P_  (.D(_02549_),
    .DE(_00066_),
    .Q(\w[63][1] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][20]$_SDFFCE_PN0P_  (.D(_02550_),
    .DE(_00066_),
    .Q(\w[63][20] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][21]$_SDFFCE_PN0P_  (.D(_02551_),
    .DE(_00066_),
    .Q(\w[63][21] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][22]$_SDFFCE_PN0P_  (.D(_02552_),
    .DE(_00066_),
    .Q(\w[63][22] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][23]$_SDFFCE_PN0P_  (.D(_02553_),
    .DE(_00066_),
    .Q(\w[63][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][24]$_SDFFCE_PN0P_  (.D(_02554_),
    .DE(_00066_),
    .Q(\w[63][24] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][25]$_SDFFCE_PN0P_  (.D(_02555_),
    .DE(_00066_),
    .Q(\w[63][25] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][26]$_SDFFCE_PN0P_  (.D(_02556_),
    .DE(_00066_),
    .Q(\w[63][26] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][27]$_SDFFCE_PN0P_  (.D(_02557_),
    .DE(_00066_),
    .Q(\w[63][27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][28]$_SDFFCE_PN0P_  (.D(_02558_),
    .DE(_00066_),
    .Q(\w[63][28] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][29]$_SDFFCE_PN0P_  (.D(_02559_),
    .DE(_00066_),
    .Q(\w[63][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][2]$_SDFFCE_PN0P_  (.D(_02560_),
    .DE(_00066_),
    .Q(\w[63][2] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][30]$_SDFFCE_PN0P_  (.D(_02561_),
    .DE(_00066_),
    .Q(\w[63][30] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][31]$_SDFFCE_PN0P_  (.D(_02562_),
    .DE(_00066_),
    .Q(\w[63][31] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][3]$_SDFFCE_PN0P_  (.D(_02563_),
    .DE(_00066_),
    .Q(\w[63][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][4]$_SDFFCE_PN0P_  (.D(_02564_),
    .DE(_00066_),
    .Q(\w[63][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][5]$_SDFFCE_PN0P_  (.D(_02565_),
    .DE(_00066_),
    .Q(\w[63][5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][6]$_SDFFCE_PN0P_  (.D(_02566_),
    .DE(_00066_),
    .Q(\w[63][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][7]$_SDFFCE_PN0P_  (.D(_02567_),
    .DE(_00066_),
    .Q(\w[63][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][8]$_SDFFCE_PN0P_  (.D(_02568_),
    .DE(_00066_),
    .Q(\w[63][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][9]$_SDFFCE_PN0P_  (.D(_02569_),
    .DE(_00066_),
    .Q(\w[63][9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][0]$_DFFE_PP_  (.D(_00513_),
    .DE(_00097_),
    .Q(\w[6][0] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][10]$_DFFE_PP_  (.D(_00514_),
    .DE(_00097_),
    .Q(\w[6][10] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][11]$_DFFE_PP_  (.D(_00515_),
    .DE(_00097_),
    .Q(\w[6][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][12]$_DFFE_PP_  (.D(_00516_),
    .DE(_00097_),
    .Q(\w[6][12] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][13]$_DFFE_PP_  (.D(_00517_),
    .DE(_00097_),
    .Q(\w[6][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][14]$_DFFE_PP_  (.D(_00518_),
    .DE(_00097_),
    .Q(\w[6][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][15]$_DFFE_PP_  (.D(_00519_),
    .DE(_00097_),
    .Q(\w[6][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][16]$_DFFE_PP_  (.D(_00520_),
    .DE(_00097_),
    .Q(\w[6][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][17]$_DFFE_PP_  (.D(_00521_),
    .DE(_00097_),
    .Q(\w[6][17] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][18]$_DFFE_PP_  (.D(_00522_),
    .DE(_00097_),
    .Q(\w[6][18] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][19]$_DFFE_PP_  (.D(_00523_),
    .DE(_00097_),
    .Q(\w[6][19] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][1]$_DFFE_PP_  (.D(_00524_),
    .DE(_00097_),
    .Q(\w[6][1] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][20]$_DFFE_PP_  (.D(_00525_),
    .DE(_00097_),
    .Q(\w[6][20] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][21]$_DFFE_PP_  (.D(_00526_),
    .DE(_00097_),
    .Q(\w[6][21] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][22]$_DFFE_PP_  (.D(_00527_),
    .DE(_00097_),
    .Q(\w[6][22] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][23]$_DFFE_PP_  (.D(_00528_),
    .DE(_00097_),
    .Q(\w[6][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][24]$_DFFE_PP_  (.D(_00529_),
    .DE(_00097_),
    .Q(\w[6][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][25]$_DFFE_PP_  (.D(_00530_),
    .DE(_00097_),
    .Q(\w[6][25] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][26]$_DFFE_PP_  (.D(_00531_),
    .DE(_00097_),
    .Q(\w[6][26] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][27]$_DFFE_PP_  (.D(_00532_),
    .DE(_00097_),
    .Q(\w[6][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][28]$_DFFE_PP_  (.D(_00533_),
    .DE(_00097_),
    .Q(\w[6][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][29]$_DFFE_PP_  (.D(_00534_),
    .DE(_00097_),
    .Q(\w[6][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][2]$_DFFE_PP_  (.D(_00535_),
    .DE(_00097_),
    .Q(\w[6][2] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][30]$_DFFE_PP_  (.D(_00536_),
    .DE(_00097_),
    .Q(\w[6][30] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][31]$_DFFE_PP_  (.D(_00537_),
    .DE(_00097_),
    .Q(\w[6][31] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][3]$_DFFE_PP_  (.D(_00538_),
    .DE(_00097_),
    .Q(\w[6][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][4]$_DFFE_PP_  (.D(_00539_),
    .DE(_00097_),
    .Q(\w[6][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][5]$_DFFE_PP_  (.D(_00540_),
    .DE(_00097_),
    .Q(\w[6][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][6]$_DFFE_PP_  (.D(_00541_),
    .DE(_00097_),
    .Q(\w[6][6] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][7]$_DFFE_PP_  (.D(_00542_),
    .DE(_00097_),
    .Q(\w[6][7] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][8]$_DFFE_PP_  (.D(_00543_),
    .DE(_00097_),
    .Q(\w[6][8] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][9]$_DFFE_PP_  (.D(_00544_),
    .DE(_00097_),
    .Q(\w[6][9] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][0]$_DFFE_PP_  (.D(_00545_),
    .DE(_00065_),
    .Q(\w[7][0] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][10]$_DFFE_PP_  (.D(_00546_),
    .DE(_00065_),
    .Q(\w[7][10] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][11]$_DFFE_PP_  (.D(_00547_),
    .DE(_00065_),
    .Q(\w[7][11] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][12]$_DFFE_PP_  (.D(_00548_),
    .DE(_00065_),
    .Q(\w[7][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][13]$_DFFE_PP_  (.D(_00549_),
    .DE(_00065_),
    .Q(\w[7][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][14]$_DFFE_PP_  (.D(_00550_),
    .DE(_00065_),
    .Q(\w[7][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][15]$_DFFE_PP_  (.D(_00551_),
    .DE(_00065_),
    .Q(\w[7][15] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][16]$_DFFE_PP_  (.D(_00552_),
    .DE(_00065_),
    .Q(\w[7][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][17]$_DFFE_PP_  (.D(_00553_),
    .DE(_00065_),
    .Q(\w[7][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][18]$_DFFE_PP_  (.D(_00554_),
    .DE(_00065_),
    .Q(\w[7][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][19]$_DFFE_PP_  (.D(_00555_),
    .DE(_00065_),
    .Q(\w[7][19] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][1]$_DFFE_PP_  (.D(_00556_),
    .DE(_00065_),
    .Q(\w[7][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][20]$_DFFE_PP_  (.D(_00557_),
    .DE(_00065_),
    .Q(\w[7][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][21]$_DFFE_PP_  (.D(_00558_),
    .DE(_00065_),
    .Q(\w[7][21] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][22]$_DFFE_PP_  (.D(_00559_),
    .DE(_00065_),
    .Q(\w[7][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][23]$_DFFE_PP_  (.D(_00560_),
    .DE(_00065_),
    .Q(\w[7][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][24]$_DFFE_PP_  (.D(_00561_),
    .DE(_00065_),
    .Q(\w[7][24] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][25]$_DFFE_PP_  (.D(_00562_),
    .DE(_00065_),
    .Q(\w[7][25] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][26]$_DFFE_PP_  (.D(_00563_),
    .DE(_00065_),
    .Q(\w[7][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][27]$_DFFE_PP_  (.D(_00564_),
    .DE(_00065_),
    .Q(\w[7][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][28]$_DFFE_PP_  (.D(_00565_),
    .DE(_00065_),
    .Q(\w[7][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][29]$_DFFE_PP_  (.D(_00566_),
    .DE(_00065_),
    .Q(\w[7][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][2]$_DFFE_PP_  (.D(_00567_),
    .DE(_00065_),
    .Q(\w[7][2] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][30]$_DFFE_PP_  (.D(_00568_),
    .DE(_00065_),
    .Q(\w[7][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][31]$_DFFE_PP_  (.D(_00569_),
    .DE(_00065_),
    .Q(\w[7][31] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][3]$_DFFE_PP_  (.D(_00570_),
    .DE(_00065_),
    .Q(\w[7][3] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][4]$_DFFE_PP_  (.D(_00571_),
    .DE(_00065_),
    .Q(\w[7][4] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][5]$_DFFE_PP_  (.D(_00572_),
    .DE(_00065_),
    .Q(\w[7][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][6]$_DFFE_PP_  (.D(_00573_),
    .DE(_00065_),
    .Q(\w[7][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][7]$_DFFE_PP_  (.D(_00574_),
    .DE(_00065_),
    .Q(\w[7][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][8]$_DFFE_PP_  (.D(_00575_),
    .DE(_00065_),
    .Q(\w[7][8] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][9]$_DFFE_PP_  (.D(_00576_),
    .DE(_00065_),
    .Q(\w[7][9] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][0]$_DFFE_PP_  (.D(_00577_),
    .DE(_00096_),
    .Q(\w[8][0] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][10]$_DFFE_PP_  (.D(_00578_),
    .DE(_00096_),
    .Q(\w[8][10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][11]$_DFFE_PP_  (.D(_00579_),
    .DE(_00096_),
    .Q(\w[8][11] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][12]$_DFFE_PP_  (.D(_00580_),
    .DE(_00096_),
    .Q(\w[8][12] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][13]$_DFFE_PP_  (.D(_00581_),
    .DE(_00096_),
    .Q(\w[8][13] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][14]$_DFFE_PP_  (.D(_00582_),
    .DE(_00096_),
    .Q(\w[8][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][15]$_DFFE_PP_  (.D(_00583_),
    .DE(_00096_),
    .Q(\w[8][15] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][16]$_DFFE_PP_  (.D(_00584_),
    .DE(_00096_),
    .Q(\w[8][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][17]$_DFFE_PP_  (.D(_00585_),
    .DE(_00096_),
    .Q(\w[8][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][18]$_DFFE_PP_  (.D(_00586_),
    .DE(_00096_),
    .Q(\w[8][18] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][19]$_DFFE_PP_  (.D(_00587_),
    .DE(_00096_),
    .Q(\w[8][19] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][1]$_DFFE_PP_  (.D(_00588_),
    .DE(_00096_),
    .Q(\w[8][1] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][20]$_DFFE_PP_  (.D(_00589_),
    .DE(_00096_),
    .Q(\w[8][20] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][21]$_DFFE_PP_  (.D(_00590_),
    .DE(_00096_),
    .Q(\w[8][21] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][22]$_DFFE_PP_  (.D(_00591_),
    .DE(_00096_),
    .Q(\w[8][22] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][23]$_DFFE_PP_  (.D(_00592_),
    .DE(_00096_),
    .Q(\w[8][23] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][24]$_DFFE_PP_  (.D(_00593_),
    .DE(_00096_),
    .Q(\w[8][24] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][25]$_DFFE_PP_  (.D(_00594_),
    .DE(_00096_),
    .Q(\w[8][25] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][26]$_DFFE_PP_  (.D(_00595_),
    .DE(_00096_),
    .Q(\w[8][26] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][27]$_DFFE_PP_  (.D(_00596_),
    .DE(_00096_),
    .Q(\w[8][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][28]$_DFFE_PP_  (.D(_00597_),
    .DE(_00096_),
    .Q(\w[8][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][29]$_DFFE_PP_  (.D(_00598_),
    .DE(_00096_),
    .Q(\w[8][29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][2]$_DFFE_PP_  (.D(_00599_),
    .DE(_00096_),
    .Q(\w[8][2] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][30]$_DFFE_PP_  (.D(_00600_),
    .DE(_00096_),
    .Q(\w[8][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][31]$_DFFE_PP_  (.D(_00601_),
    .DE(_00096_),
    .Q(\w[8][31] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][3]$_DFFE_PP_  (.D(_00602_),
    .DE(_00096_),
    .Q(\w[8][3] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][4]$_DFFE_PP_  (.D(_00603_),
    .DE(_00096_),
    .Q(\w[8][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][5]$_DFFE_PP_  (.D(_00604_),
    .DE(_00096_),
    .Q(\w[8][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][6]$_DFFE_PP_  (.D(_00605_),
    .DE(_00096_),
    .Q(\w[8][6] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][7]$_DFFE_PP_  (.D(_00606_),
    .DE(_00096_),
    .Q(\w[8][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][8]$_DFFE_PP_  (.D(_00607_),
    .DE(_00096_),
    .Q(\w[8][8] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][9]$_DFFE_PP_  (.D(_00608_),
    .DE(_00096_),
    .Q(\w[8][9] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][0]$_DFFE_PP_  (.D(_00609_),
    .DE(_00064_),
    .Q(\w[9][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][10]$_DFFE_PP_  (.D(_00610_),
    .DE(_00064_),
    .Q(\w[9][10] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][11]$_DFFE_PP_  (.D(_00611_),
    .DE(_00064_),
    .Q(\w[9][11] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][12]$_DFFE_PP_  (.D(_00612_),
    .DE(_00064_),
    .Q(\w[9][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][13]$_DFFE_PP_  (.D(_00613_),
    .DE(_00064_),
    .Q(\w[9][13] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][14]$_DFFE_PP_  (.D(_00614_),
    .DE(_00064_),
    .Q(\w[9][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][15]$_DFFE_PP_  (.D(_00615_),
    .DE(_00064_),
    .Q(\w[9][15] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][16]$_DFFE_PP_  (.D(_00616_),
    .DE(_00064_),
    .Q(\w[9][16] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][17]$_DFFE_PP_  (.D(_00617_),
    .DE(_00064_),
    .Q(\w[9][17] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][18]$_DFFE_PP_  (.D(_00618_),
    .DE(_00064_),
    .Q(\w[9][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][19]$_DFFE_PP_  (.D(_00619_),
    .DE(_00064_),
    .Q(\w[9][19] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][1]$_DFFE_PP_  (.D(_00620_),
    .DE(_00064_),
    .Q(\w[9][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][20]$_DFFE_PP_  (.D(_00621_),
    .DE(_00064_),
    .Q(\w[9][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][21]$_DFFE_PP_  (.D(_00622_),
    .DE(_00064_),
    .Q(\w[9][21] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][22]$_DFFE_PP_  (.D(_00623_),
    .DE(_00064_),
    .Q(\w[9][22] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][23]$_DFFE_PP_  (.D(_00624_),
    .DE(_00064_),
    .Q(\w[9][23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][24]$_DFFE_PP_  (.D(_00625_),
    .DE(_00064_),
    .Q(\w[9][24] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][25]$_DFFE_PP_  (.D(_00626_),
    .DE(_00064_),
    .Q(\w[9][25] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][26]$_DFFE_PP_  (.D(_00627_),
    .DE(_00064_),
    .Q(\w[9][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][27]$_DFFE_PP_  (.D(_00628_),
    .DE(_00064_),
    .Q(\w[9][27] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][28]$_DFFE_PP_  (.D(_00629_),
    .DE(_00064_),
    .Q(\w[9][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][29]$_DFFE_PP_  (.D(_00630_),
    .DE(_00064_),
    .Q(\w[9][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][2]$_DFFE_PP_  (.D(_00631_),
    .DE(_00064_),
    .Q(\w[9][2] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][30]$_DFFE_PP_  (.D(_00632_),
    .DE(_00064_),
    .Q(\w[9][30] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][31]$_DFFE_PP_  (.D(_00633_),
    .DE(_00064_),
    .Q(\w[9][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][3]$_DFFE_PP_  (.D(_00634_),
    .DE(_00064_),
    .Q(\w[9][3] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][4]$_DFFE_PP_  (.D(_00635_),
    .DE(_00064_),
    .Q(\w[9][4] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][5]$_DFFE_PP_  (.D(_00636_),
    .DE(_00064_),
    .Q(\w[9][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][6]$_DFFE_PP_  (.D(_00637_),
    .DE(_00064_),
    .Q(\w[9][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][7]$_DFFE_PP_  (.D(_00638_),
    .DE(_00064_),
    .Q(\w[9][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][8]$_DFFE_PP_  (.D(_00639_),
    .DE(_00064_),
    .Q(\w[9][8] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][9]$_DFFE_PP_  (.D(_00640_),
    .DE(_00064_),
    .Q(\w[9][9] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[0]$_DFF_P_  (.D(_00000_),
    .Q(\hash.CA1.w_i1[0] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[10]$_DFF_P_  (.D(_00001_),
    .Q(\hash.CA1.w_i1[10] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[11]$_DFF_P_  (.D(_00002_),
    .Q(\hash.CA1.w_i1[11] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[12]$_DFF_P_  (.D(_00003_),
    .Q(\hash.CA1.w_i1[12] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[13]$_DFF_P_  (.D(_00004_),
    .Q(\hash.CA1.w_i1[13] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[14]$_DFF_P_  (.D(_00005_),
    .Q(\hash.CA1.w_i1[14] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[15]$_DFF_P_  (.D(_00006_),
    .Q(\hash.CA1.w_i1[15] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[16]$_DFF_P_  (.D(_00007_),
    .Q(\hash.CA1.w_i1[16] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[17]$_DFF_P_  (.D(_00008_),
    .Q(\hash.CA1.w_i1[17] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[18]$_DFF_P_  (.D(_00009_),
    .Q(\hash.CA1.w_i1[18] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[19]$_DFF_P_  (.D(_00010_),
    .Q(\hash.CA1.w_i1[19] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[1]$_DFF_P_  (.D(_00011_),
    .Q(\hash.CA1.w_i1[1] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[20]$_DFF_P_  (.D(_00012_),
    .Q(\hash.CA1.w_i1[20] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[21]$_DFF_P_  (.D(_00013_),
    .Q(\hash.CA1.w_i1[21] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[22]$_DFF_P_  (.D(_00014_),
    .Q(\hash.CA1.w_i1[22] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[23]$_DFF_P_  (.D(_00015_),
    .Q(\hash.CA1.w_i1[23] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[24]$_DFF_P_  (.D(_00016_),
    .Q(\hash.CA1.w_i1[24] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[25]$_DFF_P_  (.D(_00017_),
    .Q(\hash.CA1.w_i1[25] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[26]$_DFF_P_  (.D(_00018_),
    .Q(\hash.CA1.w_i1[26] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[27]$_DFF_P_  (.D(_00019_),
    .Q(\hash.CA1.w_i1[27] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[28]$_DFF_P_  (.D(_00020_),
    .Q(\hash.CA1.w_i1[28] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[29]$_DFF_P_  (.D(_00021_),
    .Q(\hash.CA1.w_i1[29] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[2]$_DFF_P_  (.D(_00022_),
    .Q(\hash.CA1.w_i1[2] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[30]$_DFF_P_  (.D(_00023_),
    .Q(\hash.CA1.w_i1[30] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[31]$_DFF_P_  (.D(_00024_),
    .Q(\hash.CA1.w_i1[31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[3]$_DFF_P_  (.D(_00025_),
    .Q(\hash.CA1.w_i1[3] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[4]$_DFF_P_  (.D(_00026_),
    .Q(\hash.CA1.w_i1[4] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[5]$_DFF_P_  (.D(_00027_),
    .Q(\hash.CA1.w_i1[5] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[6]$_DFF_P_  (.D(_00028_),
    .Q(\hash.CA1.w_i1[6] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[7]$_DFF_P_  (.D(_00029_),
    .Q(\hash.CA1.w_i1[7] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[8]$_DFF_P_  (.D(_00030_),
    .Q(\hash.CA1.w_i1[8] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[9]$_DFF_P_  (.D(_00031_),
    .Q(\hash.CA1.w_i1[9] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[0]$_DFF_P_  (.D(_00032_),
    .Q(\hash.CA1.w_i2[0] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[10]$_DFF_P_  (.D(_00033_),
    .Q(\hash.CA1.w_i2[10] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[11]$_DFF_P_  (.D(_00034_),
    .Q(\hash.CA1.w_i2[11] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[12]$_DFF_P_  (.D(_00035_),
    .Q(\hash.CA1.w_i2[12] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[13]$_DFF_P_  (.D(_00036_),
    .Q(\hash.CA1.w_i2[13] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[14]$_DFF_P_  (.D(_00037_),
    .Q(\hash.CA1.w_i2[14] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[15]$_DFF_P_  (.D(_00038_),
    .Q(\hash.CA1.w_i2[15] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[16]$_DFF_P_  (.D(_00039_),
    .Q(\hash.CA1.w_i2[16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[17]$_DFF_P_  (.D(_00040_),
    .Q(\hash.CA1.w_i2[17] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[18]$_DFF_P_  (.D(_00041_),
    .Q(\hash.CA1.w_i2[18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[19]$_DFF_P_  (.D(_00042_),
    .Q(\hash.CA1.w_i2[19] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[1]$_DFF_P_  (.D(_00043_),
    .Q(\hash.CA1.w_i2[1] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[20]$_DFF_P_  (.D(_00044_),
    .Q(\hash.CA1.w_i2[20] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[21]$_DFF_P_  (.D(_00045_),
    .Q(\hash.CA1.w_i2[21] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[22]$_DFF_P_  (.D(_00046_),
    .Q(\hash.CA1.w_i2[22] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[23]$_DFF_P_  (.D(_00047_),
    .Q(\hash.CA1.w_i2[23] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[24]$_DFF_P_  (.D(_00048_),
    .Q(\hash.CA1.w_i2[24] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[25]$_DFF_P_  (.D(_00049_),
    .Q(\hash.CA1.w_i2[25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[26]$_DFF_P_  (.D(_00050_),
    .Q(\hash.CA1.w_i2[26] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[27]$_DFF_P_  (.D(_00051_),
    .Q(\hash.CA1.w_i2[27] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[28]$_DFF_P_  (.D(_00052_),
    .Q(\hash.CA1.w_i2[28] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[29]$_DFF_P_  (.D(_00053_),
    .Q(\hash.CA1.w_i2[29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[2]$_DFF_P_  (.D(_00054_),
    .Q(\hash.CA1.w_i2[2] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[30]$_DFF_P_  (.D(_00055_),
    .Q(\hash.CA1.w_i2[30] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[31]$_DFF_P_  (.D(_00056_),
    .Q(\hash.CA1.w_i2[31] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[3]$_DFF_P_  (.D(_00057_),
    .Q(\hash.CA1.w_i2[3] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[4]$_DFF_P_  (.D(_00058_),
    .Q(\hash.CA1.w_i2[4] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[5]$_DFF_P_  (.D(_00059_),
    .Q(\hash.CA1.w_i2[5] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[6]$_DFF_P_  (.D(_00060_),
    .Q(\hash.CA1.w_i2[6] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[7]$_DFF_P_  (.D(_00061_),
    .Q(\hash.CA1.w_i2[7] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[8]$_DFF_P_  (.D(_00062_),
    .Q(\hash.CA1.w_i2[8] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[9]$_DFF_P_  (.D(_00063_),
    .Q(\hash.CA1.w_i2[9] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5686 ();
 sky130_fd_sc_hd__buf_12 load_slew290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_12 load_slew291 (.A(_09875_),
    .X(net291));
 sky130_fd_sc_hd__buf_12 load_slew292 (.A(_09875_),
    .X(net292));
 sky130_fd_sc_hd__buf_12 max_cap293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_12 load_slew294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_12 load_slew295 (.A(_10373_),
    .X(net295));
 sky130_fd_sc_hd__buf_12 load_slew296 (.A(_10373_),
    .X(net296));
 sky130_fd_sc_hd__buf_12 load_slew297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_12 max_cap298 (.A(net300),
    .X(net298));
 sky130_fd_sc_hd__buf_12 load_slew299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 wire300 (.A(_09867_),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 wire301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__buf_12 load_slew302 (.A(_00071_),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_4 wire303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_12 load_slew304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__buf_12 load_slew305 (.A(_00080_),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_4 wire306 (.A(_00088_),
    .X(net306));
 sky130_fd_sc_hd__buf_12 load_slew307 (.A(_00088_),
    .X(net307));
 sky130_fd_sc_hd__buf_12 load_slew308 (.A(net310),
    .X(net308));
 sky130_fd_sc_hd__buf_12 load_slew309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_12 load_slew310 (.A(_00655_),
    .X(net310));
 sky130_fd_sc_hd__buf_12 load_slew311 (.A(_00655_),
    .X(net311));
 sky130_fd_sc_hd__buf_12 load_slew312 (.A(_00655_),
    .X(net312));
 sky130_fd_sc_hd__buf_12 load_slew313 (.A(net316),
    .X(net313));
 sky130_fd_sc_hd__buf_12 load_slew314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_12 load_slew315 (.A(net317),
    .X(net315));
 sky130_fd_sc_hd__buf_12 load_slew316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_12 load_slew317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__buf_12 load_slew318 (.A(_00657_),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_16 load_slew319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__buf_12 load_slew320 (.A(net324),
    .X(net320));
 sky130_fd_sc_hd__buf_12 load_slew321 (.A(net323),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_16 max_cap322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 wire323 (.A(net325),
    .X(net323));
 sky130_fd_sc_hd__buf_12 max_cap324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_12 load_slew325 (.A(_10352_),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_4 wire326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__buf_12 load_slew327 (.A(net332),
    .X(net327));
 sky130_fd_sc_hd__buf_12 load_slew328 (.A(net330),
    .X(net328));
 sky130_fd_sc_hd__buf_12 load_slew329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__buf_12 max_cap330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__buf_12 load_slew331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__buf_12 max_cap332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_12 load_slew333 (.A(_10348_),
    .X(net333));
 sky130_fd_sc_hd__buf_12 load_slew334 (.A(net335),
    .X(net334));
 sky130_fd_sc_hd__buf_12 load_slew335 (.A(net339),
    .X(net335));
 sky130_fd_sc_hd__buf_12 load_slew336 (.A(net338),
    .X(net336));
 sky130_fd_sc_hd__buf_12 load_slew337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_12 load_slew338 (.A(_09857_),
    .X(net338));
 sky130_fd_sc_hd__buf_12 load_slew339 (.A(_09857_),
    .X(net339));
 sky130_fd_sc_hd__buf_12 max_cap340 (.A(_09857_),
    .X(net340));
 sky130_fd_sc_hd__buf_12 max_cap341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 wire342 (.A(net346),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 wire343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__buf_12 load_slew344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_16 max_cap345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__buf_12 load_slew346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_12 load_slew347 (.A(_09854_),
    .X(net347));
 sky130_fd_sc_hd__buf_12 load_slew348 (.A(_04797_),
    .X(net348));
 sky130_fd_sc_hd__buf_12 load_slew349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__buf_12 load_slew350 (.A(\hash.reset ),
    .X(net350));
 sky130_fd_sc_hd__buf_12 load_slew351 (.A(net355),
    .X(net351));
 sky130_fd_sc_hd__buf_12 load_slew352 (.A(net354),
    .X(net352));
 sky130_fd_sc_hd__buf_12 load_slew353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 load_slew354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__buf_12 load_slew355 (.A(\hash.reset ),
    .X(net355));
 sky130_fd_sc_hd__buf_12 load_slew356 (.A(reset_hash),
    .X(net356));
 sky130_fd_sc_hd__buf_12 max_cap357 (.A(reset_hash),
    .X(net357));
 sky130_fd_sc_hd__buf_12 load_slew358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_12 load_slew359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__buf_12 load_slew360 (.A(net364),
    .X(net360));
 sky130_fd_sc_hd__buf_12 load_slew361 (.A(net363),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_16 max_cap362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 wire363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_12 load_slew364 (.A(done),
    .X(net364));
 sky130_fd_sc_hd__buf_12 load_slew365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_12 load_slew366 (.A(net372),
    .X(net366));
 sky130_fd_sc_hd__buf_12 load_slew367 (.A(net372),
    .X(net367));
 sky130_fd_sc_hd__buf_12 load_slew368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_12 load_slew369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_12 load_slew370 (.A(net372),
    .X(net370));
 sky130_fd_sc_hd__buf_12 load_slew371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_12 load_slew372 (.A(\count_hash2[1] ),
    .X(net372));
 sky130_fd_sc_hd__buf_12 load_slew373 (.A(net375),
    .X(net373));
 sky130_fd_sc_hd__buf_12 load_slew374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__buf_12 load_slew375 (.A(net379),
    .X(net375));
 sky130_fd_sc_hd__buf_12 load_slew376 (.A(net378),
    .X(net376));
 sky130_fd_sc_hd__buf_12 load_slew377 (.A(net541),
    .X(net377));
 sky130_fd_sc_hd__buf_12 load_slew378 (.A(net541),
    .X(net378));
 sky130_fd_sc_hd__buf_12 load_slew379 (.A(net541),
    .X(net379));
 sky130_fd_sc_hd__buf_12 load_slew380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__buf_12 load_slew381 (.A(\count7_2[5] ),
    .X(net381));
 sky130_fd_sc_hd__buf_12 load_slew382 (.A(\count7_2[4] ),
    .X(net382));
 sky130_fd_sc_hd__buf_12 load_slew383 (.A(net542),
    .X(net383));
 sky130_fd_sc_hd__buf_12 load_slew384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__buf_12 load_slew385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_12 load_slew386 (.A(\count7_2[3] ),
    .X(net386));
 sky130_fd_sc_hd__buf_12 load_slew387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_12 load_slew388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__buf_12 load_slew389 (.A(net393),
    .X(net389));
 sky130_fd_sc_hd__buf_12 load_slew390 (.A(net392),
    .X(net390));
 sky130_fd_sc_hd__buf_12 load_slew391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_12 load_slew392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_12 load_slew393 (.A(\count7_2[2] ),
    .X(net393));
 sky130_fd_sc_hd__buf_12 load_slew394 (.A(\count7_2[1] ),
    .X(net394));
 sky130_fd_sc_hd__buf_12 load_slew395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_12 load_slew396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_12 load_slew397 (.A(net544),
    .X(net397));
 sky130_fd_sc_hd__buf_12 load_slew398 (.A(net544),
    .X(net398));
 sky130_fd_sc_hd__buf_12 load_slew399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__buf_12 load_slew400 (.A(\count7_1[5] ),
    .X(net400));
 sky130_fd_sc_hd__buf_12 load_slew401 (.A(net545),
    .X(net401));
 sky130_fd_sc_hd__buf_12 load_slew402 (.A(\count7_1[4] ),
    .X(net402));
 sky130_fd_sc_hd__buf_12 load_slew403 (.A(\count7_1[3] ),
    .X(net403));
 sky130_fd_sc_hd__buf_12 load_slew404 (.A(net546),
    .X(net404));
 sky130_fd_sc_hd__buf_12 load_slew405 (.A(\count7_1[2] ),
    .X(net405));
 sky130_fd_sc_hd__buf_12 load_slew406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__buf_12 load_slew407 (.A(net409),
    .X(net407));
 sky130_fd_sc_hd__buf_12 max_cap408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__buf_12 load_slew409 (.A(net412),
    .X(net409));
 sky130_fd_sc_hd__buf_12 load_slew410 (.A(net412),
    .X(net410));
 sky130_fd_sc_hd__buf_12 load_slew411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_12 load_slew412 (.A(\count7_1[2] ),
    .X(net412));
 sky130_fd_sc_hd__buf_12 load_slew413 (.A(net416),
    .X(net413));
 sky130_fd_sc_hd__buf_12 load_slew414 (.A(net416),
    .X(net414));
 sky130_fd_sc_hd__buf_12 max_cap415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__buf_12 max_cap416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__buf_12 load_slew417 (.A(\count7_1[1] ),
    .X(net417));
 sky130_fd_sc_hd__buf_12 load_slew418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__buf_12 load_slew419 (.A(\count2_2[5] ),
    .X(net419));
 sky130_fd_sc_hd__buf_12 load_slew420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__buf_12 load_slew421 (.A(net548),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_4 wire422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_12 load_slew423 (.A(\count2_2[3] ),
    .X(net423));
 sky130_fd_sc_hd__buf_12 load_slew424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_12 load_slew425 (.A(\count2_2[2] ),
    .X(net425));
 sky130_fd_sc_hd__buf_12 load_slew426 (.A(net429),
    .X(net426));
 sky130_fd_sc_hd__buf_12 load_slew427 (.A(net429),
    .X(net427));
 sky130_fd_sc_hd__buf_12 load_slew428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_12 load_slew429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_12 load_slew430 (.A(\count2_2[2] ),
    .X(net430));
 sky130_fd_sc_hd__buf_12 load_slew431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_12 load_slew432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_12 load_slew433 (.A(net435),
    .X(net433));
 sky130_fd_sc_hd__buf_12 load_slew434 (.A(\count2_2[1] ),
    .X(net434));
 sky130_fd_sc_hd__buf_12 load_slew435 (.A(\count2_2[1] ),
    .X(net435));
 sky130_fd_sc_hd__buf_12 load_slew436 (.A(\count2_2[1] ),
    .X(net436));
 sky130_fd_sc_hd__buf_12 load_slew437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_12 load_slew438 (.A(\count2_1[5] ),
    .X(net438));
 sky130_fd_sc_hd__buf_12 load_slew439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_12 load_slew440 (.A(net550),
    .X(net440));
 sky130_fd_sc_hd__buf_12 load_slew441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_12 load_slew442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_12 load_slew443 (.A(\count2_1[3] ),
    .X(net443));
 sky130_fd_sc_hd__buf_12 load_slew444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_12 load_slew445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_12 load_slew446 (.A(\count2_1[2] ),
    .X(net446));
 sky130_fd_sc_hd__buf_12 load_slew447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_12 load_slew448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_12 load_slew449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_12 load_slew450 (.A(\count2_1[2] ),
    .X(net450));
 sky130_fd_sc_hd__buf_12 load_slew451 (.A(net552),
    .X(net451));
 sky130_fd_sc_hd__buf_12 load_slew452 (.A(\count2_1[1] ),
    .X(net452));
 sky130_fd_sc_hd__buf_12 load_slew453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_12 load_slew454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_12 load_slew455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_12 load_slew456 (.A(\count2_1[1] ),
    .X(net456));
 sky130_fd_sc_hd__buf_12 load_slew457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_12 load_slew458 (.A(\count16_2[5] ),
    .X(net458));
 sky130_fd_sc_hd__buf_12 load_slew459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_12 load_slew460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_12 load_slew461 (.A(\count16_2[4] ),
    .X(net461));
 sky130_fd_sc_hd__buf_12 load_slew462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_12 load_slew463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_12 load_slew464 (.A(\count16_2[3] ),
    .X(net464));
 sky130_fd_sc_hd__buf_12 load_slew465 (.A(net467),
    .X(net465));
 sky130_fd_sc_hd__buf_12 load_slew466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_12 load_slew467 (.A(net469),
    .X(net467));
 sky130_fd_sc_hd__buf_12 load_slew468 (.A(net471),
    .X(net468));
 sky130_fd_sc_hd__buf_12 load_slew469 (.A(net471),
    .X(net469));
 sky130_fd_sc_hd__buf_12 load_slew470 (.A(net472),
    .X(net470));
 sky130_fd_sc_hd__buf_12 load_slew471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_12 load_slew472 (.A(\count16_2[2] ),
    .X(net472));
 sky130_fd_sc_hd__buf_12 load_slew473 (.A(\count16_2[1] ),
    .X(net473));
 sky130_fd_sc_hd__buf_12 load_slew474 (.A(net476),
    .X(net474));
 sky130_fd_sc_hd__buf_12 load_slew475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_12 load_slew476 (.A(net553),
    .X(net476));
 sky130_fd_sc_hd__buf_12 load_slew477 (.A(\count16_2[1] ),
    .X(net477));
 sky130_fd_sc_hd__buf_12 load_slew478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__buf_12 load_slew479 (.A(\count16_1[5] ),
    .X(net479));
 sky130_fd_sc_hd__buf_12 load_slew480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_12 load_slew481 (.A(\count16_1[4] ),
    .X(net481));
 sky130_fd_sc_hd__buf_12 load_slew482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_12 load_slew483 (.A(\count16_1[3] ),
    .X(net483));
 sky130_fd_sc_hd__buf_12 load_slew484 (.A(\count16_1[3] ),
    .X(net484));
 sky130_fd_sc_hd__buf_12 load_slew485 (.A(net491),
    .X(net485));
 sky130_fd_sc_hd__buf_12 load_slew486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_12 load_slew487 (.A(net489),
    .X(net487));
 sky130_fd_sc_hd__buf_12 load_slew488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_12 load_slew489 (.A(net491),
    .X(net489));
 sky130_fd_sc_hd__buf_12 load_slew490 (.A(net555),
    .X(net490));
 sky130_fd_sc_hd__buf_12 load_slew491 (.A(\count16_1[2] ),
    .X(net491));
 sky130_fd_sc_hd__buf_12 load_slew492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_12 load_slew493 (.A(net556),
    .X(net493));
 sky130_fd_sc_hd__buf_12 load_slew494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__buf_12 load_slew495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_12 load_slew496 (.A(\count16_1[1] ),
    .X(net496));
 sky130_fd_sc_hd__buf_12 load_slew497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_12 load_slew498 (.A(\count15_2[5] ),
    .X(net498));
 sky130_fd_sc_hd__buf_12 load_slew499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_12 load_slew500 (.A(\count15_2[4] ),
    .X(net500));
 sky130_fd_sc_hd__buf_12 load_slew501 (.A(\count15_2[4] ),
    .X(net501));
 sky130_fd_sc_hd__buf_12 load_slew502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_12 load_slew503 (.A(\count15_2[3] ),
    .X(net503));
 sky130_fd_sc_hd__buf_12 load_slew504 (.A(\count15_2[3] ),
    .X(net504));
 sky130_fd_sc_hd__buf_12 load_slew505 (.A(net557),
    .X(net505));
 sky130_fd_sc_hd__buf_12 load_slew506 (.A(net511),
    .X(net506));
 sky130_fd_sc_hd__buf_12 load_slew507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_12 load_slew508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_12 load_slew509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_12 load_slew510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__buf_12 load_slew511 (.A(\count15_2[2] ),
    .X(net511));
 sky130_fd_sc_hd__buf_12 load_slew512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__buf_12 load_slew513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_12 load_slew514 (.A(net516),
    .X(net514));
 sky130_fd_sc_hd__buf_12 load_slew515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__buf_12 load_slew516 (.A(\count15_2[1] ),
    .X(net516));
 sky130_fd_sc_hd__buf_12 load_slew517 (.A(\count15_2[1] ),
    .X(net517));
 sky130_fd_sc_hd__buf_12 load_slew518 (.A(\count15_1[5] ),
    .X(net518));
 sky130_fd_sc_hd__buf_12 load_slew519 (.A(\count15_1[5] ),
    .X(net519));
 sky130_fd_sc_hd__buf_12 load_slew520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_12 load_slew521 (.A(\count15_1[4] ),
    .X(net521));
 sky130_fd_sc_hd__buf_12 load_slew522 (.A(\count15_1[3] ),
    .X(net522));
 sky130_fd_sc_hd__buf_12 load_slew523 (.A(\count15_1[3] ),
    .X(net523));
 sky130_fd_sc_hd__buf_12 load_slew524 (.A(\count15_1[3] ),
    .X(net524));
 sky130_fd_sc_hd__buf_12 load_slew525 (.A(net530),
    .X(net525));
 sky130_fd_sc_hd__buf_12 load_slew526 (.A(net528),
    .X(net526));
 sky130_fd_sc_hd__buf_12 load_slew527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__buf_12 load_slew528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__buf_12 load_slew529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__buf_12 load_slew530 (.A(\count15_1[2] ),
    .X(net530));
 sky130_fd_sc_hd__buf_12 load_slew531 (.A(net532),
    .X(net531));
 sky130_fd_sc_hd__buf_12 load_slew532 (.A(\count15_1[2] ),
    .X(net532));
 sky130_fd_sc_hd__buf_12 load_slew533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__buf_12 load_slew534 (.A(net536),
    .X(net534));
 sky130_fd_sc_hd__buf_12 load_slew535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_12 max_cap536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_12 load_slew537 (.A(\count15_1[1] ),
    .X(net537));
 sky130_fd_sc_hd__buf_12 load_slew538 (.A(_05358_),
    .X(net538));
 sky130_fd_sc_hd__buf_12 max_cap539 (.A(_08591_),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 wire540 (.A(reset_hash),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_4 wire541 (.A(\count_hash1[1] ),
    .X(net541));
 sky130_fd_sc_hd__buf_12 load_slew542 (.A(\count7_2[4] ),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_4 wire543 (.A(\count7_2[2] ),
    .X(net543));
 sky130_fd_sc_hd__buf_12 load_slew544 (.A(\count7_2[1] ),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_4 wire545 (.A(\count7_1[4] ),
    .X(net545));
 sky130_fd_sc_hd__buf_12 load_slew546 (.A(\count7_1[3] ),
    .X(net546));
 sky130_fd_sc_hd__buf_12 load_slew547 (.A(\count7_1[1] ),
    .X(net547));
 sky130_fd_sc_hd__buf_12 load_slew548 (.A(\count2_2[4] ),
    .X(net548));
 sky130_fd_sc_hd__buf_12 load_slew549 (.A(\count2_2[3] ),
    .X(net549));
 sky130_fd_sc_hd__buf_12 load_slew550 (.A(\count2_1[4] ),
    .X(net550));
 sky130_fd_sc_hd__buf_12 load_slew551 (.A(\count2_1[2] ),
    .X(net551));
 sky130_fd_sc_hd__buf_12 load_slew552 (.A(\count2_1[1] ),
    .X(net552));
 sky130_fd_sc_hd__buf_12 load_slew553 (.A(\count16_2[1] ),
    .X(net553));
 sky130_fd_sc_hd__buf_12 load_slew554 (.A(\count16_1[4] ),
    .X(net554));
 sky130_fd_sc_hd__buf_12 load_slew555 (.A(\count16_1[2] ),
    .X(net555));
 sky130_fd_sc_hd__buf_12 load_slew556 (.A(\count16_1[1] ),
    .X(net556));
 sky130_fd_sc_hd__buf_12 load_slew557 (.A(\count15_2[2] ),
    .X(net557));
 sky130_fd_sc_hd__buf_12 load_slew558 (.A(\count15_1[5] ),
    .X(net558));
 sky130_fd_sc_hd__buf_12 load_slew559 (.A(\count15_1[4] ),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_4 wire560 (.A(\count15_1[1] ),
    .X(net560));
 sky130_fd_sc_hd__buf_1 input1 (.A(message[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(message[100]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(message[101]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(message[102]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(message[103]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(message[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(message[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(message[106]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(message[107]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(message[108]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(message[109]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(message[10]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(message[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(message[111]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(message[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(message[113]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(message[114]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(message[115]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(message[116]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(message[117]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(message[118]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(message[119]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(message[11]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(message[120]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(message[121]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(message[122]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(message[123]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(message[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(message[125]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(message[126]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(message[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(message[128]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(message[129]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(message[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(message[130]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(message[131]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(message[132]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(message[133]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(message[134]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(message[135]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(message[136]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(message[137]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(message[138]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(message[139]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(message[13]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(message[140]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(message[141]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(message[142]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(message[143]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(message[144]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(message[145]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(message[146]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(message[147]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(message[148]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(message[149]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(message[14]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(message[150]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(message[151]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(message[152]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(message[153]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(message[154]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(message[155]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(message[156]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(message[157]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(message[158]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(message[159]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(message[15]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(message[160]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(message[161]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(message[162]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(message[163]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(message[164]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(message[165]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(message[166]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(message[167]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(message[168]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(message[169]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(message[16]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(message[170]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(message[171]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(message[172]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(message[173]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(message[174]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(message[175]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(message[176]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(message[177]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(message[178]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(message[179]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(message[17]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(message[180]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(message[181]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(message[182]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(message[183]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(message[184]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(message[185]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(message[186]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(message[187]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(message[188]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(message[189]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(message[18]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(message[190]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(message[191]),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input103 (.A(message[192]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(message[193]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input105 (.A(message[194]),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input106 (.A(message[195]),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(message[196]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(message[197]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(message[198]),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input110 (.A(message[199]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input111 (.A(message[19]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(message[1]),
    .X(net112));
 sky130_fd_sc_hd__buf_1 input113 (.A(message[200]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(message[201]),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(message[202]),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(message[203]),
    .X(net116));
 sky130_fd_sc_hd__buf_1 input117 (.A(message[204]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(message[205]),
    .X(net118));
 sky130_fd_sc_hd__buf_1 input119 (.A(message[206]),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input120 (.A(message[207]),
    .X(net120));
 sky130_fd_sc_hd__buf_1 input121 (.A(message[208]),
    .X(net121));
 sky130_fd_sc_hd__buf_1 input122 (.A(message[209]),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input123 (.A(message[20]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 input124 (.A(message[210]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(message[211]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(message[212]),
    .X(net126));
 sky130_fd_sc_hd__buf_1 input127 (.A(message[213]),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input128 (.A(message[214]),
    .X(net128));
 sky130_fd_sc_hd__buf_1 input129 (.A(message[215]),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input130 (.A(message[216]),
    .X(net130));
 sky130_fd_sc_hd__buf_1 input131 (.A(message[217]),
    .X(net131));
 sky130_fd_sc_hd__buf_1 input132 (.A(message[218]),
    .X(net132));
 sky130_fd_sc_hd__buf_1 input133 (.A(message[219]),
    .X(net133));
 sky130_fd_sc_hd__buf_1 input134 (.A(message[21]),
    .X(net134));
 sky130_fd_sc_hd__buf_1 input135 (.A(message[220]),
    .X(net135));
 sky130_fd_sc_hd__buf_1 input136 (.A(message[221]),
    .X(net136));
 sky130_fd_sc_hd__buf_1 input137 (.A(message[222]),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input138 (.A(message[223]),
    .X(net138));
 sky130_fd_sc_hd__buf_1 input139 (.A(message[224]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input140 (.A(message[225]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(message[226]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(message[227]),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input143 (.A(message[228]),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input144 (.A(message[229]),
    .X(net144));
 sky130_fd_sc_hd__buf_1 input145 (.A(message[22]),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(message[230]),
    .X(net146));
 sky130_fd_sc_hd__buf_1 input147 (.A(message[231]),
    .X(net147));
 sky130_fd_sc_hd__buf_1 input148 (.A(message[232]),
    .X(net148));
 sky130_fd_sc_hd__buf_1 input149 (.A(message[233]),
    .X(net149));
 sky130_fd_sc_hd__buf_1 input150 (.A(message[234]),
    .X(net150));
 sky130_fd_sc_hd__buf_1 input151 (.A(message[235]),
    .X(net151));
 sky130_fd_sc_hd__buf_1 input152 (.A(message[236]),
    .X(net152));
 sky130_fd_sc_hd__buf_1 input153 (.A(message[237]),
    .X(net153));
 sky130_fd_sc_hd__buf_1 input154 (.A(message[238]),
    .X(net154));
 sky130_fd_sc_hd__buf_1 input155 (.A(message[239]),
    .X(net155));
 sky130_fd_sc_hd__buf_1 input156 (.A(message[23]),
    .X(net156));
 sky130_fd_sc_hd__buf_1 input157 (.A(message[240]),
    .X(net157));
 sky130_fd_sc_hd__buf_1 input158 (.A(message[241]),
    .X(net158));
 sky130_fd_sc_hd__buf_1 input159 (.A(message[242]),
    .X(net159));
 sky130_fd_sc_hd__buf_1 input160 (.A(message[243]),
    .X(net160));
 sky130_fd_sc_hd__buf_1 input161 (.A(message[244]),
    .X(net161));
 sky130_fd_sc_hd__buf_1 input162 (.A(message[245]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 input163 (.A(message[246]),
    .X(net163));
 sky130_fd_sc_hd__buf_1 input164 (.A(message[247]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 input165 (.A(message[248]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input166 (.A(message[249]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 input167 (.A(message[24]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input168 (.A(message[250]),
    .X(net168));
 sky130_fd_sc_hd__buf_1 input169 (.A(message[251]),
    .X(net169));
 sky130_fd_sc_hd__buf_1 input170 (.A(message[252]),
    .X(net170));
 sky130_fd_sc_hd__buf_1 input171 (.A(message[253]),
    .X(net171));
 sky130_fd_sc_hd__buf_1 input172 (.A(message[254]),
    .X(net172));
 sky130_fd_sc_hd__buf_1 input173 (.A(message[255]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 input174 (.A(message[256]),
    .X(net174));
 sky130_fd_sc_hd__buf_1 input175 (.A(message[257]),
    .X(net175));
 sky130_fd_sc_hd__buf_1 input176 (.A(message[258]),
    .X(net176));
 sky130_fd_sc_hd__buf_1 input177 (.A(message[259]),
    .X(net177));
 sky130_fd_sc_hd__buf_1 input178 (.A(message[25]),
    .X(net178));
 sky130_fd_sc_hd__buf_1 input179 (.A(message[260]),
    .X(net179));
 sky130_fd_sc_hd__buf_1 input180 (.A(message[261]),
    .X(net180));
 sky130_fd_sc_hd__buf_1 input181 (.A(message[262]),
    .X(net181));
 sky130_fd_sc_hd__buf_1 input182 (.A(message[263]),
    .X(net182));
 sky130_fd_sc_hd__buf_1 input183 (.A(message[264]),
    .X(net183));
 sky130_fd_sc_hd__buf_1 input184 (.A(message[265]),
    .X(net184));
 sky130_fd_sc_hd__buf_1 input185 (.A(message[266]),
    .X(net185));
 sky130_fd_sc_hd__buf_1 input186 (.A(message[267]),
    .X(net186));
 sky130_fd_sc_hd__buf_1 input187 (.A(message[268]),
    .X(net187));
 sky130_fd_sc_hd__buf_1 input188 (.A(message[269]),
    .X(net188));
 sky130_fd_sc_hd__buf_1 input189 (.A(message[26]),
    .X(net189));
 sky130_fd_sc_hd__buf_1 input190 (.A(message[270]),
    .X(net190));
 sky130_fd_sc_hd__buf_1 input191 (.A(message[271]),
    .X(net191));
 sky130_fd_sc_hd__buf_1 input192 (.A(message[272]),
    .X(net192));
 sky130_fd_sc_hd__buf_1 input193 (.A(message[273]),
    .X(net193));
 sky130_fd_sc_hd__buf_1 input194 (.A(message[274]),
    .X(net194));
 sky130_fd_sc_hd__buf_1 input195 (.A(message[275]),
    .X(net195));
 sky130_fd_sc_hd__buf_1 input196 (.A(message[276]),
    .X(net196));
 sky130_fd_sc_hd__buf_1 input197 (.A(message[277]),
    .X(net197));
 sky130_fd_sc_hd__buf_1 input198 (.A(message[278]),
    .X(net198));
 sky130_fd_sc_hd__buf_1 input199 (.A(message[279]),
    .X(net199));
 sky130_fd_sc_hd__buf_1 input200 (.A(message[27]),
    .X(net200));
 sky130_fd_sc_hd__buf_1 input201 (.A(message[280]),
    .X(net201));
 sky130_fd_sc_hd__buf_1 input202 (.A(message[281]),
    .X(net202));
 sky130_fd_sc_hd__buf_1 input203 (.A(message[282]),
    .X(net203));
 sky130_fd_sc_hd__buf_1 input204 (.A(message[283]),
    .X(net204));
 sky130_fd_sc_hd__buf_1 input205 (.A(message[284]),
    .X(net205));
 sky130_fd_sc_hd__buf_1 input206 (.A(message[285]),
    .X(net206));
 sky130_fd_sc_hd__buf_1 input207 (.A(message[286]),
    .X(net207));
 sky130_fd_sc_hd__buf_1 input208 (.A(message[287]),
    .X(net208));
 sky130_fd_sc_hd__buf_1 input209 (.A(message[288]),
    .X(net209));
 sky130_fd_sc_hd__buf_1 input210 (.A(message[289]),
    .X(net210));
 sky130_fd_sc_hd__buf_1 input211 (.A(message[28]),
    .X(net211));
 sky130_fd_sc_hd__buf_1 input212 (.A(message[290]),
    .X(net212));
 sky130_fd_sc_hd__buf_1 input213 (.A(message[291]),
    .X(net213));
 sky130_fd_sc_hd__buf_1 input214 (.A(message[292]),
    .X(net214));
 sky130_fd_sc_hd__buf_1 input215 (.A(message[293]),
    .X(net215));
 sky130_fd_sc_hd__buf_1 input216 (.A(message[294]),
    .X(net216));
 sky130_fd_sc_hd__buf_1 input217 (.A(message[295]),
    .X(net217));
 sky130_fd_sc_hd__buf_1 input218 (.A(message[296]),
    .X(net218));
 sky130_fd_sc_hd__buf_1 input219 (.A(message[297]),
    .X(net219));
 sky130_fd_sc_hd__buf_1 input220 (.A(message[298]),
    .X(net220));
 sky130_fd_sc_hd__buf_1 input221 (.A(message[299]),
    .X(net221));
 sky130_fd_sc_hd__buf_1 input222 (.A(message[29]),
    .X(net222));
 sky130_fd_sc_hd__buf_1 input223 (.A(message[2]),
    .X(net223));
 sky130_fd_sc_hd__buf_1 input224 (.A(message[300]),
    .X(net224));
 sky130_fd_sc_hd__buf_1 input225 (.A(message[301]),
    .X(net225));
 sky130_fd_sc_hd__buf_1 input226 (.A(message[302]),
    .X(net226));
 sky130_fd_sc_hd__buf_1 input227 (.A(message[303]),
    .X(net227));
 sky130_fd_sc_hd__buf_1 input228 (.A(message[304]),
    .X(net228));
 sky130_fd_sc_hd__buf_1 input229 (.A(message[305]),
    .X(net229));
 sky130_fd_sc_hd__buf_1 input230 (.A(message[306]),
    .X(net230));
 sky130_fd_sc_hd__buf_1 input231 (.A(message[307]),
    .X(net231));
 sky130_fd_sc_hd__buf_1 input232 (.A(message[308]),
    .X(net232));
 sky130_fd_sc_hd__buf_1 input233 (.A(message[309]),
    .X(net233));
 sky130_fd_sc_hd__buf_1 input234 (.A(message[30]),
    .X(net234));
 sky130_fd_sc_hd__buf_1 input235 (.A(message[310]),
    .X(net235));
 sky130_fd_sc_hd__buf_1 input236 (.A(message[311]),
    .X(net236));
 sky130_fd_sc_hd__buf_1 input237 (.A(message[312]),
    .X(net237));
 sky130_fd_sc_hd__buf_1 input238 (.A(message[313]),
    .X(net238));
 sky130_fd_sc_hd__buf_1 input239 (.A(message[314]),
    .X(net239));
 sky130_fd_sc_hd__buf_1 input240 (.A(message[315]),
    .X(net240));
 sky130_fd_sc_hd__buf_1 input241 (.A(message[316]),
    .X(net241));
 sky130_fd_sc_hd__buf_1 input242 (.A(message[317]),
    .X(net242));
 sky130_fd_sc_hd__buf_1 input243 (.A(message[318]),
    .X(net243));
 sky130_fd_sc_hd__buf_1 input244 (.A(message[319]),
    .X(net244));
 sky130_fd_sc_hd__buf_1 input245 (.A(message[31]),
    .X(net245));
 sky130_fd_sc_hd__buf_1 input246 (.A(message[320]),
    .X(net246));
 sky130_fd_sc_hd__buf_1 input247 (.A(message[321]),
    .X(net247));
 sky130_fd_sc_hd__buf_1 input248 (.A(message[322]),
    .X(net248));
 sky130_fd_sc_hd__buf_1 input249 (.A(message[323]),
    .X(net249));
 sky130_fd_sc_hd__buf_1 input250 (.A(message[324]),
    .X(net250));
 sky130_fd_sc_hd__buf_1 input251 (.A(message[325]),
    .X(net251));
 sky130_fd_sc_hd__buf_1 input252 (.A(message[326]),
    .X(net252));
 sky130_fd_sc_hd__buf_1 input253 (.A(message[327]),
    .X(net253));
 sky130_fd_sc_hd__buf_1 input254 (.A(message[328]),
    .X(net254));
 sky130_fd_sc_hd__buf_1 input255 (.A(message[329]),
    .X(net255));
 sky130_fd_sc_hd__buf_1 input256 (.A(message[32]),
    .X(net256));
 sky130_fd_sc_hd__buf_1 input257 (.A(message[330]),
    .X(net257));
 sky130_fd_sc_hd__buf_1 input258 (.A(message[331]),
    .X(net258));
 sky130_fd_sc_hd__buf_1 input259 (.A(message[332]),
    .X(net259));
 sky130_fd_sc_hd__buf_1 input260 (.A(message[333]),
    .X(net260));
 sky130_fd_sc_hd__buf_1 input261 (.A(message[334]),
    .X(net261));
 sky130_fd_sc_hd__buf_1 input262 (.A(message[335]),
    .X(net262));
 sky130_fd_sc_hd__buf_1 input263 (.A(message[336]),
    .X(net263));
 sky130_fd_sc_hd__buf_1 input264 (.A(message[337]),
    .X(net264));
 sky130_fd_sc_hd__buf_1 input265 (.A(message[338]),
    .X(net265));
 sky130_fd_sc_hd__buf_1 input266 (.A(message[339]),
    .X(net266));
 sky130_fd_sc_hd__buf_1 input267 (.A(message[33]),
    .X(net267));
 sky130_fd_sc_hd__buf_1 input268 (.A(message[340]),
    .X(net268));
 sky130_fd_sc_hd__buf_1 input269 (.A(message[341]),
    .X(net269));
 sky130_fd_sc_hd__buf_1 input270 (.A(message[342]),
    .X(net270));
 sky130_fd_sc_hd__buf_1 input271 (.A(message[343]),
    .X(net271));
 sky130_fd_sc_hd__buf_1 input272 (.A(message[344]),
    .X(net272));
 sky130_fd_sc_hd__buf_1 input273 (.A(message[345]),
    .X(net273));
 sky130_fd_sc_hd__buf_1 input274 (.A(message[346]),
    .X(net274));
 sky130_fd_sc_hd__buf_1 input275 (.A(message[347]),
    .X(net275));
 sky130_fd_sc_hd__buf_1 input276 (.A(message[348]),
    .X(net276));
 sky130_fd_sc_hd__buf_1 input277 (.A(message[349]),
    .X(net277));
 sky130_fd_sc_hd__buf_1 input278 (.A(message[34]),
    .X(net278));
 sky130_fd_sc_hd__buf_1 input279 (.A(message[350]),
    .X(net279));
 sky130_fd_sc_hd__buf_1 input280 (.A(message[351]),
    .X(net280));
 sky130_fd_sc_hd__buf_1 input281 (.A(message[352]),
    .X(net281));
 sky130_fd_sc_hd__buf_1 input282 (.A(message[353]),
    .X(net282));
 sky130_fd_sc_hd__buf_1 input283 (.A(message[354]),
    .X(net283));
 sky130_fd_sc_hd__buf_1 input284 (.A(message[355]),
    .X(net284));
 sky130_fd_sc_hd__buf_1 input285 (.A(message[356]),
    .X(net285));
 sky130_fd_sc_hd__buf_1 input286 (.A(message[357]),
    .X(net286));
 sky130_fd_sc_hd__buf_1 input287 (.A(message[358]),
    .X(net287));
 sky130_fd_sc_hd__buf_1 input288 (.A(message[359]),
    .X(net288));
 sky130_fd_sc_hd__buf_1 input289 (.A(message[35]),
    .X(net289));
 sky130_fd_sc_hd__buf_1 input290 (.A(message[360]),
    .X(net561));
 sky130_fd_sc_hd__buf_1 input291 (.A(message[361]),
    .X(net562));
 sky130_fd_sc_hd__buf_1 input292 (.A(message[362]),
    .X(net563));
 sky130_fd_sc_hd__buf_1 input293 (.A(message[363]),
    .X(net564));
 sky130_fd_sc_hd__buf_1 input294 (.A(message[364]),
    .X(net565));
 sky130_fd_sc_hd__buf_1 input295 (.A(message[365]),
    .X(net566));
 sky130_fd_sc_hd__buf_1 input296 (.A(message[366]),
    .X(net567));
 sky130_fd_sc_hd__buf_1 input297 (.A(message[367]),
    .X(net568));
 sky130_fd_sc_hd__buf_1 input298 (.A(message[368]),
    .X(net569));
 sky130_fd_sc_hd__buf_1 input299 (.A(message[369]),
    .X(net570));
 sky130_fd_sc_hd__buf_1 input300 (.A(message[36]),
    .X(net571));
 sky130_fd_sc_hd__buf_1 input301 (.A(message[370]),
    .X(net572));
 sky130_fd_sc_hd__buf_1 input302 (.A(message[371]),
    .X(net573));
 sky130_fd_sc_hd__buf_1 input303 (.A(message[372]),
    .X(net574));
 sky130_fd_sc_hd__buf_1 input304 (.A(message[373]),
    .X(net575));
 sky130_fd_sc_hd__buf_1 input305 (.A(message[374]),
    .X(net576));
 sky130_fd_sc_hd__buf_1 input306 (.A(message[375]),
    .X(net577));
 sky130_fd_sc_hd__buf_1 input307 (.A(message[376]),
    .X(net578));
 sky130_fd_sc_hd__buf_1 input308 (.A(message[377]),
    .X(net579));
 sky130_fd_sc_hd__buf_1 input309 (.A(message[378]),
    .X(net580));
 sky130_fd_sc_hd__buf_1 input310 (.A(message[379]),
    .X(net581));
 sky130_fd_sc_hd__buf_1 input311 (.A(message[37]),
    .X(net582));
 sky130_fd_sc_hd__buf_1 input312 (.A(message[380]),
    .X(net583));
 sky130_fd_sc_hd__buf_1 input313 (.A(message[381]),
    .X(net584));
 sky130_fd_sc_hd__buf_1 input314 (.A(message[382]),
    .X(net585));
 sky130_fd_sc_hd__buf_1 input315 (.A(message[383]),
    .X(net586));
 sky130_fd_sc_hd__buf_1 input316 (.A(message[384]),
    .X(net587));
 sky130_fd_sc_hd__buf_1 input317 (.A(message[385]),
    .X(net588));
 sky130_fd_sc_hd__buf_1 input318 (.A(message[386]),
    .X(net589));
 sky130_fd_sc_hd__buf_1 input319 (.A(message[387]),
    .X(net590));
 sky130_fd_sc_hd__buf_1 input320 (.A(message[388]),
    .X(net591));
 sky130_fd_sc_hd__buf_1 input321 (.A(message[389]),
    .X(net592));
 sky130_fd_sc_hd__buf_1 input322 (.A(message[38]),
    .X(net593));
 sky130_fd_sc_hd__buf_1 input323 (.A(message[390]),
    .X(net594));
 sky130_fd_sc_hd__buf_1 input324 (.A(message[391]),
    .X(net595));
 sky130_fd_sc_hd__buf_1 input325 (.A(message[392]),
    .X(net596));
 sky130_fd_sc_hd__buf_1 input326 (.A(message[393]),
    .X(net597));
 sky130_fd_sc_hd__buf_1 input327 (.A(message[394]),
    .X(net598));
 sky130_fd_sc_hd__buf_1 input328 (.A(message[395]),
    .X(net599));
 sky130_fd_sc_hd__buf_1 input329 (.A(message[396]),
    .X(net600));
 sky130_fd_sc_hd__buf_1 input330 (.A(message[397]),
    .X(net601));
 sky130_fd_sc_hd__buf_1 input331 (.A(message[398]),
    .X(net602));
 sky130_fd_sc_hd__buf_1 input332 (.A(message[399]),
    .X(net603));
 sky130_fd_sc_hd__buf_1 input333 (.A(message[39]),
    .X(net604));
 sky130_fd_sc_hd__buf_1 input334 (.A(message[3]),
    .X(net605));
 sky130_fd_sc_hd__buf_1 input335 (.A(message[400]),
    .X(net606));
 sky130_fd_sc_hd__buf_1 input336 (.A(message[401]),
    .X(net607));
 sky130_fd_sc_hd__buf_1 input337 (.A(message[402]),
    .X(net608));
 sky130_fd_sc_hd__buf_1 input338 (.A(message[403]),
    .X(net609));
 sky130_fd_sc_hd__buf_1 input339 (.A(message[404]),
    .X(net610));
 sky130_fd_sc_hd__buf_1 input340 (.A(message[405]),
    .X(net611));
 sky130_fd_sc_hd__buf_1 input341 (.A(message[406]),
    .X(net612));
 sky130_fd_sc_hd__buf_1 input342 (.A(message[407]),
    .X(net613));
 sky130_fd_sc_hd__buf_1 input343 (.A(message[408]),
    .X(net614));
 sky130_fd_sc_hd__buf_1 input344 (.A(message[409]),
    .X(net615));
 sky130_fd_sc_hd__buf_1 input345 (.A(message[40]),
    .X(net616));
 sky130_fd_sc_hd__buf_1 input346 (.A(message[410]),
    .X(net617));
 sky130_fd_sc_hd__buf_1 input347 (.A(message[411]),
    .X(net618));
 sky130_fd_sc_hd__buf_1 input348 (.A(message[412]),
    .X(net619));
 sky130_fd_sc_hd__buf_1 input349 (.A(message[413]),
    .X(net620));
 sky130_fd_sc_hd__buf_1 input350 (.A(message[414]),
    .X(net621));
 sky130_fd_sc_hd__buf_1 input351 (.A(message[415]),
    .X(net622));
 sky130_fd_sc_hd__buf_1 input352 (.A(message[416]),
    .X(net623));
 sky130_fd_sc_hd__buf_1 input353 (.A(message[417]),
    .X(net624));
 sky130_fd_sc_hd__buf_1 input354 (.A(message[418]),
    .X(net625));
 sky130_fd_sc_hd__buf_1 input355 (.A(message[419]),
    .X(net626));
 sky130_fd_sc_hd__buf_1 input356 (.A(message[41]),
    .X(net627));
 sky130_fd_sc_hd__buf_1 input357 (.A(message[420]),
    .X(net628));
 sky130_fd_sc_hd__buf_1 input358 (.A(message[421]),
    .X(net629));
 sky130_fd_sc_hd__buf_1 input359 (.A(message[422]),
    .X(net630));
 sky130_fd_sc_hd__buf_1 input360 (.A(message[423]),
    .X(net631));
 sky130_fd_sc_hd__buf_1 input361 (.A(message[424]),
    .X(net632));
 sky130_fd_sc_hd__buf_1 input362 (.A(message[425]),
    .X(net633));
 sky130_fd_sc_hd__buf_1 input363 (.A(message[426]),
    .X(net634));
 sky130_fd_sc_hd__buf_1 input364 (.A(message[427]),
    .X(net635));
 sky130_fd_sc_hd__buf_1 input365 (.A(message[428]),
    .X(net636));
 sky130_fd_sc_hd__buf_1 input366 (.A(message[429]),
    .X(net637));
 sky130_fd_sc_hd__buf_1 input367 (.A(message[42]),
    .X(net638));
 sky130_fd_sc_hd__buf_1 input368 (.A(message[430]),
    .X(net639));
 sky130_fd_sc_hd__buf_1 input369 (.A(message[431]),
    .X(net640));
 sky130_fd_sc_hd__buf_1 input370 (.A(message[432]),
    .X(net641));
 sky130_fd_sc_hd__buf_1 input371 (.A(message[433]),
    .X(net642));
 sky130_fd_sc_hd__buf_1 input372 (.A(message[434]),
    .X(net643));
 sky130_fd_sc_hd__buf_1 input373 (.A(message[435]),
    .X(net644));
 sky130_fd_sc_hd__buf_1 input374 (.A(message[436]),
    .X(net645));
 sky130_fd_sc_hd__buf_1 input375 (.A(message[437]),
    .X(net646));
 sky130_fd_sc_hd__buf_1 input376 (.A(message[438]),
    .X(net647));
 sky130_fd_sc_hd__buf_1 input377 (.A(message[439]),
    .X(net648));
 sky130_fd_sc_hd__buf_1 input378 (.A(message[43]),
    .X(net649));
 sky130_fd_sc_hd__buf_1 input379 (.A(message[440]),
    .X(net650));
 sky130_fd_sc_hd__buf_1 input380 (.A(message[441]),
    .X(net651));
 sky130_fd_sc_hd__buf_1 input381 (.A(message[442]),
    .X(net652));
 sky130_fd_sc_hd__buf_1 input382 (.A(message[443]),
    .X(net653));
 sky130_fd_sc_hd__buf_1 input383 (.A(message[444]),
    .X(net654));
 sky130_fd_sc_hd__buf_1 input384 (.A(message[445]),
    .X(net655));
 sky130_fd_sc_hd__buf_1 input385 (.A(message[446]),
    .X(net656));
 sky130_fd_sc_hd__buf_1 input386 (.A(message[447]),
    .X(net657));
 sky130_fd_sc_hd__buf_1 input387 (.A(message[448]),
    .X(net658));
 sky130_fd_sc_hd__buf_1 input388 (.A(message[449]),
    .X(net659));
 sky130_fd_sc_hd__buf_1 input389 (.A(message[44]),
    .X(net660));
 sky130_fd_sc_hd__buf_1 input390 (.A(message[450]),
    .X(net661));
 sky130_fd_sc_hd__buf_1 input391 (.A(message[451]),
    .X(net662));
 sky130_fd_sc_hd__buf_1 input392 (.A(message[452]),
    .X(net663));
 sky130_fd_sc_hd__buf_1 input393 (.A(message[453]),
    .X(net664));
 sky130_fd_sc_hd__buf_1 input394 (.A(message[454]),
    .X(net665));
 sky130_fd_sc_hd__buf_1 input395 (.A(message[455]),
    .X(net666));
 sky130_fd_sc_hd__buf_1 input396 (.A(message[456]),
    .X(net667));
 sky130_fd_sc_hd__buf_1 input397 (.A(message[457]),
    .X(net668));
 sky130_fd_sc_hd__buf_1 input398 (.A(message[458]),
    .X(net669));
 sky130_fd_sc_hd__buf_1 input399 (.A(message[459]),
    .X(net670));
 sky130_fd_sc_hd__buf_1 input400 (.A(message[45]),
    .X(net671));
 sky130_fd_sc_hd__buf_1 input401 (.A(message[460]),
    .X(net672));
 sky130_fd_sc_hd__buf_1 input402 (.A(message[461]),
    .X(net673));
 sky130_fd_sc_hd__buf_1 input403 (.A(message[462]),
    .X(net674));
 sky130_fd_sc_hd__buf_1 input404 (.A(message[463]),
    .X(net675));
 sky130_fd_sc_hd__buf_1 input405 (.A(message[464]),
    .X(net676));
 sky130_fd_sc_hd__buf_1 input406 (.A(message[465]),
    .X(net677));
 sky130_fd_sc_hd__buf_1 input407 (.A(message[466]),
    .X(net678));
 sky130_fd_sc_hd__buf_1 input408 (.A(message[467]),
    .X(net679));
 sky130_fd_sc_hd__buf_1 input409 (.A(message[468]),
    .X(net680));
 sky130_fd_sc_hd__buf_1 input410 (.A(message[469]),
    .X(net681));
 sky130_fd_sc_hd__buf_1 input411 (.A(message[46]),
    .X(net682));
 sky130_fd_sc_hd__buf_1 input412 (.A(message[470]),
    .X(net683));
 sky130_fd_sc_hd__buf_1 input413 (.A(message[471]),
    .X(net684));
 sky130_fd_sc_hd__buf_1 input414 (.A(message[472]),
    .X(net685));
 sky130_fd_sc_hd__buf_1 input415 (.A(message[473]),
    .X(net686));
 sky130_fd_sc_hd__buf_1 input416 (.A(message[474]),
    .X(net687));
 sky130_fd_sc_hd__buf_1 input417 (.A(message[475]),
    .X(net688));
 sky130_fd_sc_hd__buf_1 input418 (.A(message[476]),
    .X(net689));
 sky130_fd_sc_hd__buf_1 input419 (.A(message[477]),
    .X(net690));
 sky130_fd_sc_hd__buf_1 input420 (.A(message[478]),
    .X(net691));
 sky130_fd_sc_hd__buf_1 input421 (.A(message[479]),
    .X(net692));
 sky130_fd_sc_hd__buf_1 input422 (.A(message[47]),
    .X(net693));
 sky130_fd_sc_hd__buf_1 input423 (.A(message[480]),
    .X(net694));
 sky130_fd_sc_hd__buf_1 input424 (.A(message[481]),
    .X(net695));
 sky130_fd_sc_hd__buf_1 input425 (.A(message[482]),
    .X(net696));
 sky130_fd_sc_hd__buf_1 input426 (.A(message[483]),
    .X(net697));
 sky130_fd_sc_hd__buf_1 input427 (.A(message[484]),
    .X(net698));
 sky130_fd_sc_hd__buf_1 input428 (.A(message[485]),
    .X(net699));
 sky130_fd_sc_hd__buf_1 input429 (.A(message[486]),
    .X(net700));
 sky130_fd_sc_hd__buf_1 input430 (.A(message[487]),
    .X(net701));
 sky130_fd_sc_hd__buf_1 input431 (.A(message[488]),
    .X(net702));
 sky130_fd_sc_hd__buf_1 input432 (.A(message[489]),
    .X(net703));
 sky130_fd_sc_hd__buf_1 input433 (.A(message[48]),
    .X(net704));
 sky130_fd_sc_hd__buf_1 input434 (.A(message[490]),
    .X(net705));
 sky130_fd_sc_hd__buf_1 input435 (.A(message[491]),
    .X(net706));
 sky130_fd_sc_hd__buf_1 input436 (.A(message[492]),
    .X(net707));
 sky130_fd_sc_hd__buf_1 input437 (.A(message[493]),
    .X(net708));
 sky130_fd_sc_hd__buf_1 input438 (.A(message[494]),
    .X(net709));
 sky130_fd_sc_hd__buf_1 input439 (.A(message[495]),
    .X(net710));
 sky130_fd_sc_hd__buf_1 input440 (.A(message[496]),
    .X(net711));
 sky130_fd_sc_hd__buf_1 input441 (.A(message[497]),
    .X(net712));
 sky130_fd_sc_hd__buf_1 input442 (.A(message[498]),
    .X(net713));
 sky130_fd_sc_hd__buf_1 input443 (.A(message[499]),
    .X(net714));
 sky130_fd_sc_hd__buf_1 input444 (.A(message[49]),
    .X(net715));
 sky130_fd_sc_hd__buf_1 input445 (.A(message[4]),
    .X(net716));
 sky130_fd_sc_hd__buf_1 input446 (.A(message[500]),
    .X(net717));
 sky130_fd_sc_hd__buf_1 input447 (.A(message[501]),
    .X(net718));
 sky130_fd_sc_hd__buf_1 input448 (.A(message[502]),
    .X(net719));
 sky130_fd_sc_hd__buf_1 input449 (.A(message[503]),
    .X(net720));
 sky130_fd_sc_hd__buf_1 input450 (.A(message[504]),
    .X(net721));
 sky130_fd_sc_hd__buf_1 input451 (.A(message[505]),
    .X(net722));
 sky130_fd_sc_hd__buf_1 input452 (.A(message[506]),
    .X(net723));
 sky130_fd_sc_hd__buf_1 input453 (.A(message[507]),
    .X(net724));
 sky130_fd_sc_hd__buf_1 input454 (.A(message[508]),
    .X(net725));
 sky130_fd_sc_hd__buf_1 input455 (.A(message[509]),
    .X(net726));
 sky130_fd_sc_hd__buf_1 input456 (.A(message[50]),
    .X(net727));
 sky130_fd_sc_hd__buf_1 input457 (.A(message[510]),
    .X(net728));
 sky130_fd_sc_hd__buf_1 input458 (.A(message[511]),
    .X(net729));
 sky130_fd_sc_hd__buf_1 input459 (.A(message[51]),
    .X(net730));
 sky130_fd_sc_hd__buf_1 input460 (.A(message[52]),
    .X(net731));
 sky130_fd_sc_hd__buf_1 input461 (.A(message[53]),
    .X(net732));
 sky130_fd_sc_hd__buf_1 input462 (.A(message[54]),
    .X(net733));
 sky130_fd_sc_hd__buf_1 input463 (.A(message[55]),
    .X(net734));
 sky130_fd_sc_hd__buf_1 input464 (.A(message[56]),
    .X(net735));
 sky130_fd_sc_hd__buf_1 input465 (.A(message[57]),
    .X(net736));
 sky130_fd_sc_hd__buf_1 input466 (.A(message[58]),
    .X(net737));
 sky130_fd_sc_hd__buf_1 input467 (.A(message[59]),
    .X(net738));
 sky130_fd_sc_hd__buf_1 input468 (.A(message[5]),
    .X(net739));
 sky130_fd_sc_hd__buf_1 input469 (.A(message[60]),
    .X(net740));
 sky130_fd_sc_hd__buf_1 input470 (.A(message[61]),
    .X(net741));
 sky130_fd_sc_hd__buf_1 input471 (.A(message[62]),
    .X(net742));
 sky130_fd_sc_hd__buf_1 input472 (.A(message[63]),
    .X(net743));
 sky130_fd_sc_hd__buf_1 input473 (.A(message[64]),
    .X(net744));
 sky130_fd_sc_hd__buf_1 input474 (.A(message[65]),
    .X(net745));
 sky130_fd_sc_hd__buf_1 input475 (.A(message[66]),
    .X(net746));
 sky130_fd_sc_hd__buf_1 input476 (.A(message[67]),
    .X(net747));
 sky130_fd_sc_hd__buf_1 input477 (.A(message[68]),
    .X(net748));
 sky130_fd_sc_hd__buf_1 input478 (.A(message[69]),
    .X(net749));
 sky130_fd_sc_hd__buf_1 input479 (.A(message[6]),
    .X(net750));
 sky130_fd_sc_hd__buf_1 input480 (.A(message[70]),
    .X(net751));
 sky130_fd_sc_hd__buf_1 input481 (.A(message[71]),
    .X(net752));
 sky130_fd_sc_hd__buf_1 input482 (.A(message[72]),
    .X(net753));
 sky130_fd_sc_hd__buf_1 input483 (.A(message[73]),
    .X(net754));
 sky130_fd_sc_hd__buf_1 input484 (.A(message[74]),
    .X(net755));
 sky130_fd_sc_hd__buf_1 input485 (.A(message[75]),
    .X(net756));
 sky130_fd_sc_hd__buf_1 input486 (.A(message[76]),
    .X(net757));
 sky130_fd_sc_hd__buf_1 input487 (.A(message[77]),
    .X(net758));
 sky130_fd_sc_hd__buf_1 input488 (.A(message[78]),
    .X(net759));
 sky130_fd_sc_hd__buf_1 input489 (.A(message[79]),
    .X(net760));
 sky130_fd_sc_hd__buf_1 input490 (.A(message[7]),
    .X(net761));
 sky130_fd_sc_hd__buf_1 input491 (.A(message[80]),
    .X(net762));
 sky130_fd_sc_hd__buf_1 input492 (.A(message[81]),
    .X(net763));
 sky130_fd_sc_hd__buf_1 input493 (.A(message[82]),
    .X(net764));
 sky130_fd_sc_hd__buf_1 input494 (.A(message[83]),
    .X(net765));
 sky130_fd_sc_hd__buf_1 input495 (.A(message[84]),
    .X(net766));
 sky130_fd_sc_hd__buf_1 input496 (.A(message[85]),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input497 (.A(message[86]),
    .X(net768));
 sky130_fd_sc_hd__buf_1 input498 (.A(message[87]),
    .X(net769));
 sky130_fd_sc_hd__buf_1 input499 (.A(message[88]),
    .X(net770));
 sky130_fd_sc_hd__buf_1 input500 (.A(message[89]),
    .X(net771));
 sky130_fd_sc_hd__buf_1 input501 (.A(message[8]),
    .X(net772));
 sky130_fd_sc_hd__buf_1 input502 (.A(message[90]),
    .X(net773));
 sky130_fd_sc_hd__buf_1 input503 (.A(message[91]),
    .X(net774));
 sky130_fd_sc_hd__buf_1 input504 (.A(message[92]),
    .X(net775));
 sky130_fd_sc_hd__buf_1 input505 (.A(message[93]),
    .X(net776));
 sky130_fd_sc_hd__buf_1 input506 (.A(message[94]),
    .X(net777));
 sky130_fd_sc_hd__buf_1 input507 (.A(message[95]),
    .X(net778));
 sky130_fd_sc_hd__buf_1 input508 (.A(message[96]),
    .X(net779));
 sky130_fd_sc_hd__buf_1 input509 (.A(message[97]),
    .X(net780));
 sky130_fd_sc_hd__buf_1 input510 (.A(message[98]),
    .X(net781));
 sky130_fd_sc_hd__buf_1 input511 (.A(message[99]),
    .X(net782));
 sky130_fd_sc_hd__buf_1 input512 (.A(message[9]),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_1 input513 (.A(reset),
    .X(net784));
 sky130_fd_sc_hd__buf_1 output514 (.A(net785),
    .X(hashvalue[0]));
 sky130_fd_sc_hd__buf_1 output515 (.A(net786),
    .X(hashvalue[100]));
 sky130_fd_sc_hd__buf_1 output516 (.A(net787),
    .X(hashvalue[101]));
 sky130_fd_sc_hd__buf_1 output517 (.A(net788),
    .X(hashvalue[102]));
 sky130_fd_sc_hd__buf_1 output518 (.A(net789),
    .X(hashvalue[103]));
 sky130_fd_sc_hd__buf_1 output519 (.A(net790),
    .X(hashvalue[104]));
 sky130_fd_sc_hd__buf_1 output520 (.A(net791),
    .X(hashvalue[105]));
 sky130_fd_sc_hd__buf_1 output521 (.A(net792),
    .X(hashvalue[106]));
 sky130_fd_sc_hd__buf_1 output522 (.A(net793),
    .X(hashvalue[107]));
 sky130_fd_sc_hd__buf_1 output523 (.A(net794),
    .X(hashvalue[108]));
 sky130_fd_sc_hd__buf_1 output524 (.A(net795),
    .X(hashvalue[109]));
 sky130_fd_sc_hd__buf_1 output525 (.A(net796),
    .X(hashvalue[10]));
 sky130_fd_sc_hd__buf_1 output526 (.A(net797),
    .X(hashvalue[110]));
 sky130_fd_sc_hd__buf_1 output527 (.A(net798),
    .X(hashvalue[111]));
 sky130_fd_sc_hd__buf_1 output528 (.A(net799),
    .X(hashvalue[112]));
 sky130_fd_sc_hd__buf_1 output529 (.A(net800),
    .X(hashvalue[113]));
 sky130_fd_sc_hd__buf_1 output530 (.A(net801),
    .X(hashvalue[114]));
 sky130_fd_sc_hd__buf_1 output531 (.A(net802),
    .X(hashvalue[115]));
 sky130_fd_sc_hd__buf_1 output532 (.A(net803),
    .X(hashvalue[116]));
 sky130_fd_sc_hd__buf_1 output533 (.A(net804),
    .X(hashvalue[117]));
 sky130_fd_sc_hd__buf_1 output534 (.A(net805),
    .X(hashvalue[118]));
 sky130_fd_sc_hd__buf_1 output535 (.A(net806),
    .X(hashvalue[119]));
 sky130_fd_sc_hd__buf_1 output536 (.A(net807),
    .X(hashvalue[11]));
 sky130_fd_sc_hd__buf_1 output537 (.A(net808),
    .X(hashvalue[120]));
 sky130_fd_sc_hd__buf_1 output538 (.A(net809),
    .X(hashvalue[121]));
 sky130_fd_sc_hd__buf_1 output539 (.A(net810),
    .X(hashvalue[122]));
 sky130_fd_sc_hd__buf_1 output540 (.A(net811),
    .X(hashvalue[123]));
 sky130_fd_sc_hd__buf_1 output541 (.A(net812),
    .X(hashvalue[124]));
 sky130_fd_sc_hd__buf_1 output542 (.A(net813),
    .X(hashvalue[125]));
 sky130_fd_sc_hd__buf_1 output543 (.A(net814),
    .X(hashvalue[126]));
 sky130_fd_sc_hd__buf_1 output544 (.A(net815),
    .X(hashvalue[127]));
 sky130_fd_sc_hd__buf_1 output545 (.A(net816),
    .X(hashvalue[128]));
 sky130_fd_sc_hd__buf_1 output546 (.A(net817),
    .X(hashvalue[129]));
 sky130_fd_sc_hd__buf_1 output547 (.A(net818),
    .X(hashvalue[12]));
 sky130_fd_sc_hd__buf_1 output548 (.A(net819),
    .X(hashvalue[130]));
 sky130_fd_sc_hd__buf_1 output549 (.A(net820),
    .X(hashvalue[131]));
 sky130_fd_sc_hd__buf_1 output550 (.A(net821),
    .X(hashvalue[132]));
 sky130_fd_sc_hd__buf_1 output551 (.A(net822),
    .X(hashvalue[133]));
 sky130_fd_sc_hd__buf_1 output552 (.A(net823),
    .X(hashvalue[134]));
 sky130_fd_sc_hd__buf_1 output553 (.A(net824),
    .X(hashvalue[135]));
 sky130_fd_sc_hd__buf_1 output554 (.A(net825),
    .X(hashvalue[136]));
 sky130_fd_sc_hd__buf_1 output555 (.A(net826),
    .X(hashvalue[137]));
 sky130_fd_sc_hd__buf_1 output556 (.A(net827),
    .X(hashvalue[138]));
 sky130_fd_sc_hd__buf_1 output557 (.A(net828),
    .X(hashvalue[139]));
 sky130_fd_sc_hd__buf_1 output558 (.A(net829),
    .X(hashvalue[13]));
 sky130_fd_sc_hd__buf_1 output559 (.A(net830),
    .X(hashvalue[140]));
 sky130_fd_sc_hd__buf_1 output560 (.A(net831),
    .X(hashvalue[141]));
 sky130_fd_sc_hd__buf_1 output561 (.A(net832),
    .X(hashvalue[142]));
 sky130_fd_sc_hd__buf_1 output562 (.A(net833),
    .X(hashvalue[143]));
 sky130_fd_sc_hd__buf_1 output563 (.A(net834),
    .X(hashvalue[144]));
 sky130_fd_sc_hd__buf_1 output564 (.A(net835),
    .X(hashvalue[145]));
 sky130_fd_sc_hd__buf_1 output565 (.A(net836),
    .X(hashvalue[146]));
 sky130_fd_sc_hd__buf_1 output566 (.A(net837),
    .X(hashvalue[147]));
 sky130_fd_sc_hd__buf_1 output567 (.A(net838),
    .X(hashvalue[148]));
 sky130_fd_sc_hd__buf_1 output568 (.A(net839),
    .X(hashvalue[149]));
 sky130_fd_sc_hd__buf_1 output569 (.A(net840),
    .X(hashvalue[14]));
 sky130_fd_sc_hd__buf_1 output570 (.A(net841),
    .X(hashvalue[150]));
 sky130_fd_sc_hd__buf_1 output571 (.A(net842),
    .X(hashvalue[151]));
 sky130_fd_sc_hd__buf_1 output572 (.A(net843),
    .X(hashvalue[152]));
 sky130_fd_sc_hd__buf_1 output573 (.A(net844),
    .X(hashvalue[153]));
 sky130_fd_sc_hd__buf_1 output574 (.A(net845),
    .X(hashvalue[154]));
 sky130_fd_sc_hd__buf_1 output575 (.A(net846),
    .X(hashvalue[155]));
 sky130_fd_sc_hd__buf_1 output576 (.A(net847),
    .X(hashvalue[156]));
 sky130_fd_sc_hd__buf_1 output577 (.A(net848),
    .X(hashvalue[157]));
 sky130_fd_sc_hd__buf_1 output578 (.A(net849),
    .X(hashvalue[158]));
 sky130_fd_sc_hd__buf_1 output579 (.A(net850),
    .X(hashvalue[159]));
 sky130_fd_sc_hd__buf_1 output580 (.A(net851),
    .X(hashvalue[15]));
 sky130_fd_sc_hd__buf_1 output581 (.A(net852),
    .X(hashvalue[160]));
 sky130_fd_sc_hd__buf_1 output582 (.A(net853),
    .X(hashvalue[161]));
 sky130_fd_sc_hd__buf_1 output583 (.A(net854),
    .X(hashvalue[162]));
 sky130_fd_sc_hd__buf_1 output584 (.A(net855),
    .X(hashvalue[163]));
 sky130_fd_sc_hd__buf_1 output585 (.A(net856),
    .X(hashvalue[164]));
 sky130_fd_sc_hd__buf_1 output586 (.A(net857),
    .X(hashvalue[165]));
 sky130_fd_sc_hd__buf_1 output587 (.A(net858),
    .X(hashvalue[166]));
 sky130_fd_sc_hd__buf_1 output588 (.A(net859),
    .X(hashvalue[167]));
 sky130_fd_sc_hd__buf_1 output589 (.A(net860),
    .X(hashvalue[168]));
 sky130_fd_sc_hd__buf_1 output590 (.A(net861),
    .X(hashvalue[169]));
 sky130_fd_sc_hd__buf_1 output591 (.A(net862),
    .X(hashvalue[16]));
 sky130_fd_sc_hd__buf_1 output592 (.A(net863),
    .X(hashvalue[170]));
 sky130_fd_sc_hd__buf_1 output593 (.A(net864),
    .X(hashvalue[171]));
 sky130_fd_sc_hd__buf_1 output594 (.A(net865),
    .X(hashvalue[172]));
 sky130_fd_sc_hd__buf_1 output595 (.A(net866),
    .X(hashvalue[173]));
 sky130_fd_sc_hd__buf_1 output596 (.A(net867),
    .X(hashvalue[174]));
 sky130_fd_sc_hd__buf_1 output597 (.A(net868),
    .X(hashvalue[175]));
 sky130_fd_sc_hd__buf_1 output598 (.A(net869),
    .X(hashvalue[176]));
 sky130_fd_sc_hd__buf_1 output599 (.A(net870),
    .X(hashvalue[177]));
 sky130_fd_sc_hd__buf_1 output600 (.A(net871),
    .X(hashvalue[178]));
 sky130_fd_sc_hd__buf_1 output601 (.A(net872),
    .X(hashvalue[179]));
 sky130_fd_sc_hd__buf_1 output602 (.A(net873),
    .X(hashvalue[17]));
 sky130_fd_sc_hd__buf_1 output603 (.A(net874),
    .X(hashvalue[180]));
 sky130_fd_sc_hd__buf_1 output604 (.A(net875),
    .X(hashvalue[181]));
 sky130_fd_sc_hd__buf_1 output605 (.A(net876),
    .X(hashvalue[182]));
 sky130_fd_sc_hd__buf_1 output606 (.A(net877),
    .X(hashvalue[183]));
 sky130_fd_sc_hd__buf_1 output607 (.A(net878),
    .X(hashvalue[184]));
 sky130_fd_sc_hd__buf_1 output608 (.A(net879),
    .X(hashvalue[185]));
 sky130_fd_sc_hd__buf_1 output609 (.A(net880),
    .X(hashvalue[186]));
 sky130_fd_sc_hd__buf_1 output610 (.A(net881),
    .X(hashvalue[187]));
 sky130_fd_sc_hd__buf_1 output611 (.A(net882),
    .X(hashvalue[188]));
 sky130_fd_sc_hd__buf_1 output612 (.A(net883),
    .X(hashvalue[189]));
 sky130_fd_sc_hd__buf_1 output613 (.A(net884),
    .X(hashvalue[18]));
 sky130_fd_sc_hd__buf_1 output614 (.A(net885),
    .X(hashvalue[190]));
 sky130_fd_sc_hd__buf_1 output615 (.A(net886),
    .X(hashvalue[191]));
 sky130_fd_sc_hd__buf_1 output616 (.A(net887),
    .X(hashvalue[192]));
 sky130_fd_sc_hd__buf_1 output617 (.A(net888),
    .X(hashvalue[193]));
 sky130_fd_sc_hd__buf_1 output618 (.A(net889),
    .X(hashvalue[194]));
 sky130_fd_sc_hd__buf_1 output619 (.A(net890),
    .X(hashvalue[195]));
 sky130_fd_sc_hd__buf_1 output620 (.A(net891),
    .X(hashvalue[196]));
 sky130_fd_sc_hd__buf_1 output621 (.A(net892),
    .X(hashvalue[197]));
 sky130_fd_sc_hd__buf_1 output622 (.A(net893),
    .X(hashvalue[198]));
 sky130_fd_sc_hd__buf_1 output623 (.A(net894),
    .X(hashvalue[199]));
 sky130_fd_sc_hd__buf_1 output624 (.A(net895),
    .X(hashvalue[19]));
 sky130_fd_sc_hd__buf_1 output625 (.A(net896),
    .X(hashvalue[1]));
 sky130_fd_sc_hd__buf_1 output626 (.A(net897),
    .X(hashvalue[200]));
 sky130_fd_sc_hd__buf_1 output627 (.A(net898),
    .X(hashvalue[201]));
 sky130_fd_sc_hd__buf_1 output628 (.A(net899),
    .X(hashvalue[202]));
 sky130_fd_sc_hd__buf_1 output629 (.A(net900),
    .X(hashvalue[203]));
 sky130_fd_sc_hd__buf_1 output630 (.A(net901),
    .X(hashvalue[204]));
 sky130_fd_sc_hd__buf_1 output631 (.A(net902),
    .X(hashvalue[205]));
 sky130_fd_sc_hd__buf_1 output632 (.A(net903),
    .X(hashvalue[206]));
 sky130_fd_sc_hd__buf_1 output633 (.A(net904),
    .X(hashvalue[207]));
 sky130_fd_sc_hd__buf_1 output634 (.A(net905),
    .X(hashvalue[208]));
 sky130_fd_sc_hd__buf_1 output635 (.A(net906),
    .X(hashvalue[209]));
 sky130_fd_sc_hd__buf_1 output636 (.A(net907),
    .X(hashvalue[20]));
 sky130_fd_sc_hd__buf_1 output637 (.A(net908),
    .X(hashvalue[210]));
 sky130_fd_sc_hd__buf_1 output638 (.A(net909),
    .X(hashvalue[211]));
 sky130_fd_sc_hd__buf_1 output639 (.A(net910),
    .X(hashvalue[212]));
 sky130_fd_sc_hd__buf_1 output640 (.A(net911),
    .X(hashvalue[213]));
 sky130_fd_sc_hd__buf_1 output641 (.A(net912),
    .X(hashvalue[214]));
 sky130_fd_sc_hd__buf_1 output642 (.A(net913),
    .X(hashvalue[215]));
 sky130_fd_sc_hd__buf_1 output643 (.A(net914),
    .X(hashvalue[216]));
 sky130_fd_sc_hd__buf_1 output644 (.A(net915),
    .X(hashvalue[217]));
 sky130_fd_sc_hd__buf_1 output645 (.A(net916),
    .X(hashvalue[218]));
 sky130_fd_sc_hd__buf_1 output646 (.A(net917),
    .X(hashvalue[219]));
 sky130_fd_sc_hd__buf_1 output647 (.A(net918),
    .X(hashvalue[21]));
 sky130_fd_sc_hd__buf_1 output648 (.A(net919),
    .X(hashvalue[220]));
 sky130_fd_sc_hd__buf_1 output649 (.A(net920),
    .X(hashvalue[221]));
 sky130_fd_sc_hd__buf_1 output650 (.A(net921),
    .X(hashvalue[222]));
 sky130_fd_sc_hd__buf_1 output651 (.A(net922),
    .X(hashvalue[223]));
 sky130_fd_sc_hd__buf_1 output652 (.A(net923),
    .X(hashvalue[224]));
 sky130_fd_sc_hd__buf_1 output653 (.A(net924),
    .X(hashvalue[225]));
 sky130_fd_sc_hd__buf_1 output654 (.A(net925),
    .X(hashvalue[226]));
 sky130_fd_sc_hd__buf_1 output655 (.A(net926),
    .X(hashvalue[227]));
 sky130_fd_sc_hd__buf_1 output656 (.A(net927),
    .X(hashvalue[228]));
 sky130_fd_sc_hd__buf_1 output657 (.A(net928),
    .X(hashvalue[229]));
 sky130_fd_sc_hd__buf_1 output658 (.A(net929),
    .X(hashvalue[22]));
 sky130_fd_sc_hd__buf_1 output659 (.A(net930),
    .X(hashvalue[230]));
 sky130_fd_sc_hd__buf_1 output660 (.A(net931),
    .X(hashvalue[231]));
 sky130_fd_sc_hd__buf_1 output661 (.A(net932),
    .X(hashvalue[232]));
 sky130_fd_sc_hd__buf_1 output662 (.A(net933),
    .X(hashvalue[233]));
 sky130_fd_sc_hd__buf_1 output663 (.A(net934),
    .X(hashvalue[234]));
 sky130_fd_sc_hd__buf_1 output664 (.A(net935),
    .X(hashvalue[235]));
 sky130_fd_sc_hd__buf_1 output665 (.A(net936),
    .X(hashvalue[236]));
 sky130_fd_sc_hd__buf_1 output666 (.A(net937),
    .X(hashvalue[237]));
 sky130_fd_sc_hd__buf_1 output667 (.A(net938),
    .X(hashvalue[238]));
 sky130_fd_sc_hd__buf_1 output668 (.A(net939),
    .X(hashvalue[239]));
 sky130_fd_sc_hd__buf_1 output669 (.A(net940),
    .X(hashvalue[23]));
 sky130_fd_sc_hd__buf_1 output670 (.A(net941),
    .X(hashvalue[240]));
 sky130_fd_sc_hd__buf_1 output671 (.A(net942),
    .X(hashvalue[241]));
 sky130_fd_sc_hd__buf_1 output672 (.A(net943),
    .X(hashvalue[242]));
 sky130_fd_sc_hd__buf_1 output673 (.A(net944),
    .X(hashvalue[243]));
 sky130_fd_sc_hd__buf_1 output674 (.A(net945),
    .X(hashvalue[244]));
 sky130_fd_sc_hd__buf_1 output675 (.A(net946),
    .X(hashvalue[245]));
 sky130_fd_sc_hd__buf_1 output676 (.A(net947),
    .X(hashvalue[246]));
 sky130_fd_sc_hd__buf_1 output677 (.A(net948),
    .X(hashvalue[247]));
 sky130_fd_sc_hd__buf_1 output678 (.A(net949),
    .X(hashvalue[248]));
 sky130_fd_sc_hd__buf_1 output679 (.A(net950),
    .X(hashvalue[249]));
 sky130_fd_sc_hd__buf_1 output680 (.A(net951),
    .X(hashvalue[24]));
 sky130_fd_sc_hd__buf_1 output681 (.A(net952),
    .X(hashvalue[250]));
 sky130_fd_sc_hd__buf_1 output682 (.A(net953),
    .X(hashvalue[251]));
 sky130_fd_sc_hd__buf_1 output683 (.A(net954),
    .X(hashvalue[252]));
 sky130_fd_sc_hd__buf_1 output684 (.A(net955),
    .X(hashvalue[253]));
 sky130_fd_sc_hd__buf_1 output685 (.A(net956),
    .X(hashvalue[254]));
 sky130_fd_sc_hd__buf_1 output686 (.A(net957),
    .X(hashvalue[255]));
 sky130_fd_sc_hd__buf_1 output687 (.A(net958),
    .X(hashvalue[25]));
 sky130_fd_sc_hd__buf_1 output688 (.A(net959),
    .X(hashvalue[26]));
 sky130_fd_sc_hd__buf_1 output689 (.A(net960),
    .X(hashvalue[27]));
 sky130_fd_sc_hd__buf_1 output690 (.A(net961),
    .X(hashvalue[28]));
 sky130_fd_sc_hd__buf_1 output691 (.A(net962),
    .X(hashvalue[29]));
 sky130_fd_sc_hd__buf_1 output692 (.A(net963),
    .X(hashvalue[2]));
 sky130_fd_sc_hd__buf_1 output693 (.A(net964),
    .X(hashvalue[30]));
 sky130_fd_sc_hd__buf_1 output694 (.A(net965),
    .X(hashvalue[31]));
 sky130_fd_sc_hd__buf_1 output695 (.A(net966),
    .X(hashvalue[32]));
 sky130_fd_sc_hd__buf_1 output696 (.A(net967),
    .X(hashvalue[33]));
 sky130_fd_sc_hd__buf_1 output697 (.A(net968),
    .X(hashvalue[34]));
 sky130_fd_sc_hd__buf_1 output698 (.A(net969),
    .X(hashvalue[35]));
 sky130_fd_sc_hd__buf_1 output699 (.A(net970),
    .X(hashvalue[36]));
 sky130_fd_sc_hd__buf_1 output700 (.A(net971),
    .X(hashvalue[37]));
 sky130_fd_sc_hd__buf_1 output701 (.A(net972),
    .X(hashvalue[38]));
 sky130_fd_sc_hd__buf_1 output702 (.A(net973),
    .X(hashvalue[39]));
 sky130_fd_sc_hd__buf_1 output703 (.A(net974),
    .X(hashvalue[3]));
 sky130_fd_sc_hd__buf_1 output704 (.A(net975),
    .X(hashvalue[40]));
 sky130_fd_sc_hd__buf_1 output705 (.A(net976),
    .X(hashvalue[41]));
 sky130_fd_sc_hd__buf_1 output706 (.A(net977),
    .X(hashvalue[42]));
 sky130_fd_sc_hd__buf_1 output707 (.A(net978),
    .X(hashvalue[43]));
 sky130_fd_sc_hd__buf_1 output708 (.A(net979),
    .X(hashvalue[44]));
 sky130_fd_sc_hd__buf_1 output709 (.A(net980),
    .X(hashvalue[45]));
 sky130_fd_sc_hd__buf_1 output710 (.A(net981),
    .X(hashvalue[46]));
 sky130_fd_sc_hd__buf_1 output711 (.A(net982),
    .X(hashvalue[47]));
 sky130_fd_sc_hd__buf_1 output712 (.A(net983),
    .X(hashvalue[48]));
 sky130_fd_sc_hd__buf_1 output713 (.A(net984),
    .X(hashvalue[49]));
 sky130_fd_sc_hd__buf_1 output714 (.A(net985),
    .X(hashvalue[4]));
 sky130_fd_sc_hd__buf_1 output715 (.A(net986),
    .X(hashvalue[50]));
 sky130_fd_sc_hd__buf_1 output716 (.A(net987),
    .X(hashvalue[51]));
 sky130_fd_sc_hd__buf_1 output717 (.A(net988),
    .X(hashvalue[52]));
 sky130_fd_sc_hd__buf_1 output718 (.A(net989),
    .X(hashvalue[53]));
 sky130_fd_sc_hd__buf_1 output719 (.A(net990),
    .X(hashvalue[54]));
 sky130_fd_sc_hd__buf_1 output720 (.A(net991),
    .X(hashvalue[55]));
 sky130_fd_sc_hd__buf_1 output721 (.A(net992),
    .X(hashvalue[56]));
 sky130_fd_sc_hd__buf_1 output722 (.A(net993),
    .X(hashvalue[57]));
 sky130_fd_sc_hd__buf_1 output723 (.A(net994),
    .X(hashvalue[58]));
 sky130_fd_sc_hd__buf_1 output724 (.A(net995),
    .X(hashvalue[59]));
 sky130_fd_sc_hd__buf_1 output725 (.A(net996),
    .X(hashvalue[5]));
 sky130_fd_sc_hd__buf_1 output726 (.A(net997),
    .X(hashvalue[60]));
 sky130_fd_sc_hd__buf_1 output727 (.A(net998),
    .X(hashvalue[61]));
 sky130_fd_sc_hd__buf_1 output728 (.A(net999),
    .X(hashvalue[62]));
 sky130_fd_sc_hd__buf_1 output729 (.A(net1000),
    .X(hashvalue[63]));
 sky130_fd_sc_hd__buf_1 output730 (.A(net1001),
    .X(hashvalue[64]));
 sky130_fd_sc_hd__buf_1 output731 (.A(net1002),
    .X(hashvalue[65]));
 sky130_fd_sc_hd__buf_1 output732 (.A(net1003),
    .X(hashvalue[66]));
 sky130_fd_sc_hd__buf_1 output733 (.A(net1004),
    .X(hashvalue[67]));
 sky130_fd_sc_hd__buf_1 output734 (.A(net1005),
    .X(hashvalue[68]));
 sky130_fd_sc_hd__buf_1 output735 (.A(net1006),
    .X(hashvalue[69]));
 sky130_fd_sc_hd__buf_1 output736 (.A(net1007),
    .X(hashvalue[6]));
 sky130_fd_sc_hd__buf_1 output737 (.A(net1008),
    .X(hashvalue[70]));
 sky130_fd_sc_hd__buf_1 output738 (.A(net1009),
    .X(hashvalue[71]));
 sky130_fd_sc_hd__buf_1 output739 (.A(net1010),
    .X(hashvalue[72]));
 sky130_fd_sc_hd__buf_1 output740 (.A(net1011),
    .X(hashvalue[73]));
 sky130_fd_sc_hd__buf_1 output741 (.A(net1012),
    .X(hashvalue[74]));
 sky130_fd_sc_hd__buf_1 output742 (.A(net1013),
    .X(hashvalue[75]));
 sky130_fd_sc_hd__buf_1 output743 (.A(net1014),
    .X(hashvalue[76]));
 sky130_fd_sc_hd__buf_1 output744 (.A(net1015),
    .X(hashvalue[77]));
 sky130_fd_sc_hd__buf_1 output745 (.A(net1016),
    .X(hashvalue[78]));
 sky130_fd_sc_hd__buf_1 output746 (.A(net1017),
    .X(hashvalue[79]));
 sky130_fd_sc_hd__buf_1 output747 (.A(net1018),
    .X(hashvalue[7]));
 sky130_fd_sc_hd__buf_1 output748 (.A(net1019),
    .X(hashvalue[80]));
 sky130_fd_sc_hd__buf_1 output749 (.A(net1020),
    .X(hashvalue[81]));
 sky130_fd_sc_hd__buf_1 output750 (.A(net1021),
    .X(hashvalue[82]));
 sky130_fd_sc_hd__buf_1 output751 (.A(net1022),
    .X(hashvalue[83]));
 sky130_fd_sc_hd__buf_1 output752 (.A(net1023),
    .X(hashvalue[84]));
 sky130_fd_sc_hd__buf_1 output753 (.A(net1024),
    .X(hashvalue[85]));
 sky130_fd_sc_hd__buf_1 output754 (.A(net1025),
    .X(hashvalue[86]));
 sky130_fd_sc_hd__buf_1 output755 (.A(net1026),
    .X(hashvalue[87]));
 sky130_fd_sc_hd__buf_1 output756 (.A(net1027),
    .X(hashvalue[88]));
 sky130_fd_sc_hd__buf_1 output757 (.A(net1028),
    .X(hashvalue[89]));
 sky130_fd_sc_hd__buf_1 output758 (.A(net1029),
    .X(hashvalue[8]));
 sky130_fd_sc_hd__buf_1 output759 (.A(net1030),
    .X(hashvalue[90]));
 sky130_fd_sc_hd__buf_1 output760 (.A(net1031),
    .X(hashvalue[91]));
 sky130_fd_sc_hd__buf_1 output761 (.A(net1032),
    .X(hashvalue[92]));
 sky130_fd_sc_hd__buf_1 output762 (.A(net1033),
    .X(hashvalue[93]));
 sky130_fd_sc_hd__buf_1 output763 (.A(net1034),
    .X(hashvalue[94]));
 sky130_fd_sc_hd__buf_1 output764 (.A(net1035),
    .X(hashvalue[95]));
 sky130_fd_sc_hd__buf_1 output765 (.A(net1036),
    .X(hashvalue[96]));
 sky130_fd_sc_hd__buf_1 output766 (.A(net1037),
    .X(hashvalue[97]));
 sky130_fd_sc_hd__buf_1 output767 (.A(net1038),
    .X(hashvalue[98]));
 sky130_fd_sc_hd__buf_1 output768 (.A(net1039),
    .X(hashvalue[99]));
 sky130_fd_sc_hd__buf_1 output769 (.A(net1040),
    .X(hashvalue[9]));
 sky130_fd_sc_hd__buf_1 output770 (.A(net1041),
    .X(ready));
 sky130_fd_sc_hd__buf_8 load_slew771 (.A(_05430_),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_1 load_slew772 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_1 load_slew773 (.A(net784),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_274_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_275_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_278_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_280_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_282_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_285_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_286_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_287_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_288_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload1 (.A(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload2 (.A(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload3 (.A(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload6 (.A(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload7 (.A(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload8 (.A(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload11 (.A(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload12 (.A(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload13 (.A(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload14 (.A(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload15 (.A(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload16 (.A(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload17 (.A(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload18 (.A(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload19 (.A(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload20 (.A(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload21 (.A(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload22 (.A(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload23 (.A(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload24 (.A(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload25 (.A(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload26 (.A(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload27 (.A(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__clkinv_1 clkload28 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload29 (.A(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload30 (.A(clknet_leaf_282_clk));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload32 (.A(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload33 (.A(clknet_leaf_285_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload34 (.A(clknet_leaf_287_clk));
 sky130_fd_sc_hd__clkinv_1 clkload35 (.A(clknet_leaf_288_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload36 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_4 clkload37 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__bufinv_16 clkload38 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__bufinv_16 clkload39 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_2 clkload40 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload41 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload42 (.A(clknet_leaf_279_clk));
 sky130_fd_sc_hd__bufinv_16 clkload43 (.A(clknet_leaf_280_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkinv_1 clkload45 (.A(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkinv_1 clkload46 (.A(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload47 (.A(clknet_leaf_270_clk));
 sky130_fd_sc_hd__bufinv_16 clkload48 (.A(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkinv_4 clkload49 (.A(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkinv_1 clkload50 (.A(clknet_leaf_274_clk));
 sky130_fd_sc_hd__clkinv_1 clkload51 (.A(clknet_leaf_275_clk));
 sky130_fd_sc_hd__clkinv_1 clkload52 (.A(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkinv_2 clkload53 (.A(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkinv_1 clkload54 (.A(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkinv_2 clkload55 (.A(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkinv_2 clkload56 (.A(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkinv_2 clkload57 (.A(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload58 (.A(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload59 (.A(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkinv_1 clkload60 (.A(clknet_leaf_265_clk));
 sky130_fd_sc_hd__bufinv_16 clkload61 (.A(clknet_leaf_277_clk));
 sky130_fd_sc_hd__bufinv_16 clkload62 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__bufinv_16 clkload63 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinv_2 clkload64 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload65 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__bufinv_16 clkload66 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkinv_1 clkload67 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_1 clkload68 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_1 clkload69 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload70 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkinv_2 clkload71 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload72 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinv_1 clkload73 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload74 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_1 clkload75 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__bufinv_16 clkload76 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload77 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload78 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__bufinv_16 clkload79 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__bufinv_16 clkload80 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload81 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload82 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_2 clkload83 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload84 (.A(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload85 (.A(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload86 (.A(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload87 (.A(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkinv_2 clkload88 (.A(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload89 (.A(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkinv_4 clkload90 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload91 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_4 clkload92 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__inv_8 clkload93 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload94 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload95 (.A(clknet_leaf_247_clk));
 sky130_fd_sc_hd__bufinv_16 clkload96 (.A(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload97 (.A(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload98 (.A(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload99 (.A(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkinv_2 clkload100 (.A(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload101 (.A(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload102 (.A(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload103 (.A(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkinv_2 clkload104 (.A(clknet_leaf_219_clk));
 sky130_fd_sc_hd__bufinv_16 clkload105 (.A(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload106 (.A(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload107 (.A(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkinv_4 clkload108 (.A(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkinv_1 clkload109 (.A(clknet_leaf_233_clk));
 sky130_fd_sc_hd__bufinv_16 clkload110 (.A(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload111 (.A(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload112 (.A(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload113 (.A(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload114 (.A(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkinv_1 clkload115 (.A(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload116 (.A(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkinv_1 clkload117 (.A(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload118 (.A(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload119 (.A(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkinv_2 clkload120 (.A(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload121 (.A(clknet_leaf_202_clk));
 sky130_fd_sc_hd__inv_6 clkload122 (.A(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkinv_2 clkload123 (.A(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload124 (.A(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload125 (.A(clknet_leaf_207_clk));
 sky130_fd_sc_hd__bufinv_16 clkload126 (.A(clknet_leaf_217_clk));
 sky130_fd_sc_hd__bufinv_16 clkload127 (.A(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkinv_4 clkload128 (.A(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload129 (.A(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkinv_4 clkload130 (.A(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkinv_1 clkload131 (.A(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkinv_2 clkload132 (.A(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkinv_1 clkload133 (.A(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload134 (.A(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload135 (.A(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload136 (.A(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload137 (.A(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload138 (.A(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload139 (.A(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload140 (.A(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload141 (.A(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkinv_4 clkload142 (.A(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload143 (.A(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload144 (.A(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkinv_1 clkload145 (.A(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkinv_1 clkload146 (.A(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkinv_1 clkload147 (.A(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload148 (.A(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkinv_2 clkload149 (.A(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkinv_2 clkload150 (.A(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload151 (.A(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload152 (.A(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload153 (.A(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload154 (.A(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkinv_2 clkload155 (.A(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload156 (.A(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkinv_4 clkload157 (.A(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload158 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload159 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload160 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload161 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload162 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload163 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinv_2 clkload164 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload165 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__bufinv_16 clkload166 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkinv_2 clkload167 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_2 clkload168 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_4 clkload169 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__bufinv_16 clkload170 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkinv_2 clkload171 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkinv_2 clkload172 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__bufinv_16 clkload173 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__bufinv_16 clkload174 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkinv_2 clkload175 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__inv_6 clkload176 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkinv_1 clkload177 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkinv_1 clkload178 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload179 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkinv_2 clkload180 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__bufinv_16 clkload181 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkinv_2 clkload182 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__bufinv_16 clkload183 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinv_2 clkload184 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload185 (.A(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkinv_1 clkload186 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkinv_1 clkload187 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__bufinv_16 clkload188 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinv_1 clkload189 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__bufinv_16 clkload190 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkinv_1 clkload191 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkinv_2 clkload192 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkinv_4 clkload193 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkinv_2 clkload194 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload195 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkinv_1 clkload196 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload197 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkinv_1 clkload198 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_1 clkload199 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkinv_1 clkload200 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload201 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__bufinv_16 clkload202 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkinv_2 clkload203 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__bufinv_16 clkload204 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkinv_1 clkload205 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__bufinv_16 clkload206 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkinv_1 clkload207 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__bufinv_16 clkload208 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload209 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_1 clkload210 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkinv_1 clkload211 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload212 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload213 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload214 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkinv_1 clkload215 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload216 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkinv_2 clkload217 (.A(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload218 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload219 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload220 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkinv_2 clkload221 (.A(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload222 (.A(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload223 (.A(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload224 (.A(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload225 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload226 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload227 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload228 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload229 (.A(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload230 (.A(clknet_leaf_158_clk));
 sky130_fd_sc_hd__bufinv_16 clkload231 (.A(clknet_leaf_159_clk));
 sky130_fd_sc_hd__bufinv_16 clkload232 (.A(clknet_leaf_161_clk));
 sky130_fd_sc_hd__bufinv_16 clkload233 (.A(clknet_leaf_162_clk));
 sky130_fd_sc_hd__inv_6 clkload234 (.A(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload235 (.A(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkinv_4 clkload236 (.A(clknet_leaf_165_clk));
 sky130_fd_sc_hd__bufinv_16 clkload237 (.A(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload238 (.A(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload239 (.A(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload240 (.A(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload241 (.A(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload242 (.A(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload243 (.A(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload244 (.A(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkinv_2 clkload245 (.A(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload246 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload247 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__bufinv_16 clkload248 (.A(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload249 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload250 (.A(clknet_leaf_123_clk));
 sky130_fd_sc_hd__bufinv_16 clkload251 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload252 (.A(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload253 (.A(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkinv_2 clkload254 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkinv_1 clkload255 (.A(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload256 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload257 (.A(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkinv_2 clkload258 (.A(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload259 (.A(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkinv_2 clkload260 (.A(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload261 (.A(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkinv_1 clkload262 (.A(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload263 (.A(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkinv_2 clkload264 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkinv_2 clkload265 (.A(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload266 (.A(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkinv_1 clkload267 (.A(clknet_leaf_144_clk));
 sky130_fd_sc_hd__bufinv_16 clkload268 (.A(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkinv_4 clkload269 (.A(clknet_leaf_149_clk));
 sky130_fd_sc_hd__bufinv_16 clkload270 (.A(clknet_leaf_150_clk));
 sky130_fd_sc_hd__bufinv_16 clkload271 (.A(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload272 (.A(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload273 (.A(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkinv_1 clkload274 (.A(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload275 (.A(clknet_leaf_147_clk));
 sky130_fd_sc_hd__inv_6 clkload276 (.A(clknet_leaf_148_clk));
 sky130_fd_sc_hd__buf_2 rebuffer1 (.A(\hash.CA1.S1.X[30] ),
    .X(net1045));
 sky130_fd_sc_hd__buf_2 rebuffer2 (.A(\hash.CA1.S1.X[30] ),
    .X(net1046));
 sky130_fd_sc_hd__buf_2 rebuffer3 (.A(net1046),
    .X(net1047));
 sky130_fd_sc_hd__buf_2 rebuffer4 (.A(net1081),
    .X(net1048));
 sky130_fd_sc_hd__buf_2 rebuffer5 (.A(_13237_),
    .X(net1049));
 sky130_fd_sc_hd__buf_2 rebuffer6 (.A(_06705_),
    .X(net1050));
 sky130_fd_sc_hd__buf_2 rebuffer7 (.A(_13288_),
    .X(net1051));
 sky130_fd_sc_hd__buf_2 rebuffer8 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__nor2_2 clone9 (.A(net1085),
    .B(net351),
    .Y(net1053));
 sky130_fd_sc_hd__nor2_2 clone10 (.A(_06688_),
    .B(net352),
    .Y(net1054));
 sky130_fd_sc_hd__buf_2 rebuffer11 (.A(_13231_),
    .X(net1055));
 sky130_fd_sc_hd__buf_4 rebuffer12 (.A(\hash.CA1.S0.X[25] ),
    .X(net1056));
 sky130_fd_sc_hd__buf_2 rebuffer13 (.A(_04509_),
    .X(net1057));
 sky130_fd_sc_hd__buf_2 rebuffer14 (.A(\hash.CA2.S1.X[7] ),
    .X(net1058));
 sky130_fd_sc_hd__buf_2 rebuffer15 (.A(net1106),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 rebuffer16 (.A(net1059),
    .X(net1060));
 sky130_fd_sc_hd__buf_2 rebuffer17 (.A(net1059),
    .X(net1061));
 sky130_fd_sc_hd__buf_2 rebuffer18 (.A(\hash.CA2.S1.X[7] ),
    .X(net1062));
 sky130_fd_sc_hd__buf_2 rebuffer19 (.A(\hash.CA2.S1.X[26] ),
    .X(net1063));
 sky130_fd_sc_hd__buf_2 rebuffer20 (.A(\hash.CA2.S1.X[26] ),
    .X(net1064));
 sky130_fd_sc_hd__buf_2 rebuffer21 (.A(\hash.CA2.S1.X[26] ),
    .X(net1065));
 sky130_fd_sc_hd__buf_2 rebuffer22 (.A(net1065),
    .X(net1066));
 sky130_fd_sc_hd__buf_2 rebuffer23 (.A(_13330_),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 rebuffer24 (.A(_04710_),
    .X(net1068));
 sky130_fd_sc_hd__buf_2 rebuffer25 (.A(_06727_),
    .X(net1069));
 sky130_fd_sc_hd__buf_2 rebuffer26 (.A(\hash.CA2.S1.X[25] ),
    .X(net1070));
 sky130_fd_sc_hd__buf_2 rebuffer27 (.A(\hash.CA2.S1.X[25] ),
    .X(net1071));
 sky130_fd_sc_hd__buf_2 rebuffer28 (.A(\hash.CA2.S1.X[25] ),
    .X(net1072));
 sky130_fd_sc_hd__buf_2 rebuffer34 (.A(_13379_),
    .X(net1078));
 sky130_fd_sc_hd__buf_2 rebuffer35 (.A(_13379_),
    .X(net1079));
 sky130_fd_sc_hd__buf_2 rebuffer63 (.A(_04402_),
    .X(net1112));
 sky130_fd_sc_hd__buf_1 rebuffer37 (.A(_06952_),
    .X(net1081));
 sky130_fd_sc_hd__buf_2 rebuffer38 (.A(_13414_),
    .X(net1082));
 sky130_fd_sc_hd__buf_2 rebuffer39 (.A(_12086_),
    .X(net1083));
 sky130_fd_sc_hd__buf_2 rebuffer40 (.A(_04710_),
    .X(net1084));
 sky130_fd_sc_hd__buf_2 rebuffer41 (.A(_06682_),
    .X(net1085));
 sky130_fd_sc_hd__buf_2 rebuffer45 (.A(net1112),
    .X(net1089));
 sky130_fd_sc_hd__buf_2 rebuffer46 (.A(_04549_),
    .X(net1090));
 sky130_fd_sc_hd__buf_4 rebuffer47 (.A(_04461_),
    .X(net1091));
 sky130_fd_sc_hd__buf_4 rebuffer48 (.A(_04475_),
    .X(net1092));
 sky130_fd_sc_hd__buf_2 rebuffer49 (.A(net1092),
    .X(net1093));
 sky130_fd_sc_hd__buf_8 rebuffer50 (.A(_06201_),
    .X(net1094));
 sky130_fd_sc_hd__buf_2 rebuffer51 (.A(net1094),
    .X(net1095));
 sky130_fd_sc_hd__buf_2 rebuffer52 (.A(net1095),
    .X(net1096));
 sky130_fd_sc_hd__buf_2 rebuffer53 (.A(_12081_),
    .X(net1097));
 sky130_fd_sc_hd__buf_4 rebuffer54 (.A(_06055_),
    .X(net1098));
 sky130_fd_sc_hd__buf_2 rebuffer55 (.A(_04427_),
    .X(net1099));
 sky130_fd_sc_hd__mux2i_4 clone56 (.A0(\w[63][24] ),
    .A1(_05325_),
    .S(_04797_),
    .Y(net1100));
 sky130_fd_sc_hd__a21oi_4 clone57 (.A1(\w[63][28] ),
    .A2(net360),
    .B1(_05371_),
    .Y(net1101));
 sky130_fd_sc_hd__a21oi_4 clone58 (.A1(\w[63][18] ),
    .A2(net358),
    .B1(_05266_),
    .Y(net1102));
 sky130_fd_sc_hd__clkbuf_4 wire1 (.A(_05639_),
    .X(net1073));
 sky130_fd_sc_hd__buf_6 rebuffer9 (.A(_04654_),
    .X(net1074));
 sky130_fd_sc_hd__buf_1 rebuffer10 (.A(_09560_),
    .X(net1075));
 sky130_fd_sc_hd__buf_1 rebuffer42 (.A(_04635_),
    .X(net1103));
 sky130_fd_sc_hd__buf_2 rebuffer43 (.A(_13316_),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 rebuffer44 (.A(_13461_),
    .X(net1105));
 sky130_fd_sc_hd__buf_2 rebuffer56 (.A(\hash.CA2.S1.X[7] ),
    .X(net1106));
 sky130_fd_sc_hd__buf_6 rebuffer64 (.A(_04588_),
    .X(net1113));
 sky130_fd_sc_hd__buf_2 rebuffer65 (.A(_04481_),
    .X(net1114));
 sky130_fd_sc_hd__buf_1 rebuffer74 (.A(_09265_),
    .X(net1123));
 sky130_fd_sc_hd__a21oi_4 clone80 (.A1(\w[63][30] ),
    .A2(net360),
    .B1(_05388_),
    .Y(net1129));
 sky130_fd_sc_hd__buf_12 rebuffer81 (.A(_03120_),
    .X(net1130));
 sky130_fd_sc_hd__buf_12 rebuffer82 (.A(_02994_),
    .X(net1131));
 sky130_fd_sc_hd__buf_2 rebuffer83 (.A(net1131),
    .X(net1132));
 sky130_fd_sc_hd__buf_2 rebuffer84 (.A(net1131),
    .X(net1133));
 sky130_fd_sc_hd__buf_12 rebuffer85 (.A(_05389_),
    .X(net1134));
 sky130_fd_sc_hd__a21oi_4 clone86 (.A1(\w[63][16] ),
    .A2(net359),
    .B1(_05246_),
    .Y(net1135));
 sky130_fd_sc_hd__a21oi_2 clone87 (.A1(\w[63][14] ),
    .A2(net358),
    .B1(_05227_),
    .Y(net1136));
 sky130_fd_sc_hd__mux2i_4 clone88 (.A0(\w[63][24] ),
    .A1(_05325_),
    .S(_04797_),
    .Y(net1137));
 sky130_fd_sc_hd__mux2i_4 clone89 (.A0(\w[62][28] ),
    .A1(_05034_),
    .S(net348),
    .Y(net1138));
 sky130_fd_sc_hd__a21oi_2 clone90 (.A1(\w[62][24] ),
    .A2(net361),
    .B1(_04999_),
    .Y(net1139));
 sky130_fd_sc_hd__buf_12 rebuffer91 (.A(_03005_),
    .X(net1140));
 sky130_fd_sc_hd__buf_2 rebuffer92 (.A(net1140),
    .X(net1141));
 sky130_fd_sc_hd__a21oi_2 clone93 (.A1(\w[63][28] ),
    .A2(net360),
    .B1(_05371_),
    .Y(net1142));
 sky130_fd_sc_hd__mux2i_2 clone94 (.A0(\w[62][29] ),
    .A1(_05043_),
    .S(net348),
    .Y(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_00026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_00027_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_11604_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_11645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_11661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_11676_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_11796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_12019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\hash.CA1.w_i1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\hash.CA1.w_i1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_00032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_00032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_00032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_00032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_00057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_00022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_00056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_00056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_11891_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(\hash.CA2.f_dash[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(_08973_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1328 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1220 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1292 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1300 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1164 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1077 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1137 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1372 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1241 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1396 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1150 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1144 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1320 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1304 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1343 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1352 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1304 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_983 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1386 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1394 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1402 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1050 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1150 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1232 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1340 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1410 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1271 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1326 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1377 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1402 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1268 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1282 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1326 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1374 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1263 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1294 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1384 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1238 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1243 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1285 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1341 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1257 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1316 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1387 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1400 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1172 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1292 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1300 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1316 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1410 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1414 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1314 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1244 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1298 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1324 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1387 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1395 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1402 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1293 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1396 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1202 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1244 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1328 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1172 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1308 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1361 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1296 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1363 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_998 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1312 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1344 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1328 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1271 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1322 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1368 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1341 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1390 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1326 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1404 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1107 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1338 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1398 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1406 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1370 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1362 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1177 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_687 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1232 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1394 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1262 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1341 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1377 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1350 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1274 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1295 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1309 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1371 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1375 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_994 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1177 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1223 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1263 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1396 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_902 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1013 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1270 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1340 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1354 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1050 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1398 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1414 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1191 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1317 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1372 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1126 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1341 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1385 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_846 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_954 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1295 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1408 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_927 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1243 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1284 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1347 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1191 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1326 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1374 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1290 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1341 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1352 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1376 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1191 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_948 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1304 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1352 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1361 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1036 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1326 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1384 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1044 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1052 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1208 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1362 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_930 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1363 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1375 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1387 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1392 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1408 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1418 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1296 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1344 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1022 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1194 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1220 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1370 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1290 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1298 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1312 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1396 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1396 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1184 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1357 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1150 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1146 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1160 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1309 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1360 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1387 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_846 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1140 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1243 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1363 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1414 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1193 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1290 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1343 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1394 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_654 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1317 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1332 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1374 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1298 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1390 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1006 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_923 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1140 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1017 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1300 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1372 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1384 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1328 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1406 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1421 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1194 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1256 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1326 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1271 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1413 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1268 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_5 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1418 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1361 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1372 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1368 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1384 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1100 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1184 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1302 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1347 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1282 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1384 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1300 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1334 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1103 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1317 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1334 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1120 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1230 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1363 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1366 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1275 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1292 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1190 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1251 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1309 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_872 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1232 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1303 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1405 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1082 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1131 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1384 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1385 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_930 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1287 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1407 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1200 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1382 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1396 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1144 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1384 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1414 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1293 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1266 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1280 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1360 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1107 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1164 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1172 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1232 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1256 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1274 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1300 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1414 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1266 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1308 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1339 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1047 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1293 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_654 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1212 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1361 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1128 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1267 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1372 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1412 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1126 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1303 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_954 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1316 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1052 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1208 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1190 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1316 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1401 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1369 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1163 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1372 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1326 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1350 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1064 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1308 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1414 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1340 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1369 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1403 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1031 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1264 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1221 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1275 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1298 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1328 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1311 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1362 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1374 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1294 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1339 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1286 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1283 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1360 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1250 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1310 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1391 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1044 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1251 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1312 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1382 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1293 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1372 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_687 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1276 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1311 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_908 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1350 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1358 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1320 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1373 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1406 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1026 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1347 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1383 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1421 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1047 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1295 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1363 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1406 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1418 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_906 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1275 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1328 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1403 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1410 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1044 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1274 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1310 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1414 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1287 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1312 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1358 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1420 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1107 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1163 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1410 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1414 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1375 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1395 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1404 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_902 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_687 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1401 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_964 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1177 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1202 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1405 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1031 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1403 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1410 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1418 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1421 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1013 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1202 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1232 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1254 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_927 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1212 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1190 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1421 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1022 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1421 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1421 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1164 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1077 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1142 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_930 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1022 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1013 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_946 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1421 ();
endmodule
