module sha256_unrolled_pipelined (clk,
    ready,
    reset,
    hashvalue,
    message);
 input clk;
 output ready;
 input reset;
 output [255:0] hashvalue;
 input [0:511] message;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02328_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02346_;
 wire _02351_;
 wire _02354_;
 wire _02357_;
 wire _02360_;
 wire _02363_;
 wire _02366_;
 wire _02369_;
 wire _02372_;
 wire _02375_;
 wire _02377_;
 wire _02378_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02407_;
 wire _02408_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02463_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02471_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02484_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02495_;
 wire _02496_;
 wire _02498_;
 wire _02499_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02528_;
 wire _02529_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02584_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02592_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02736_;
 wire _02742_;
 wire _02743_;
 wire _02745_;
 wire _02746_;
 wire _02753_;
 wire _02759_;
 wire _02760_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02781_;
 wire _02787_;
 wire _02788_;
 wire _02790_;
 wire _02791_;
 wire _02798_;
 wire _02804_;
 wire _02805_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02851_;
 wire _02853_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02879_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02910_;
 wire _02911_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02963_;
 wire _02965_;
 wire _02966_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03172_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03210_;
 wire _03212_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03223_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03241_;
 wire _03242_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03254_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03464_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03504_;
 wire _03539_;
 wire _03543_;
 wire _03547_;
 wire _03551_;
 wire _03555_;
 wire _03559_;
 wire _03564_;
 wire _03568_;
 wire _03572_;
 wire _03576_;
 wire _03580_;
 wire _03584_;
 wire _03588_;
 wire _03592_;
 wire _03596_;
 wire _03600_;
 wire _03604_;
 wire _03608_;
 wire _03613_;
 wire _03649_;
 wire _03684_;
 wire _03688_;
 wire _03692_;
 wire _03696_;
 wire _03700_;
 wire _03704_;
 wire _03708_;
 wire _03712_;
 wire _03716_;
 wire _03720_;
 wire _03724_;
 wire _03728_;
 wire _03732_;
 wire _03736_;
 wire _03740_;
 wire _03744_;
 wire _03748_;
 wire _03752_;
 wire _03757_;
 wire _03761_;
 wire _03765_;
 wire _03769_;
 wire _03773_;
 wire _03777_;
 wire _03781_;
 wire _03785_;
 wire _03793_;
 wire _03797_;
 wire _03801_;
 wire _03804_;
 wire _03808_;
 wire _03811_;
 wire _03814_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03871_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03894_;
 wire _03896_;
 wire _03897_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03926_;
 wire _03928_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03992_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04015_;
 wire _04017_;
 wire _04018_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04047_;
 wire _04049_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04178_;
 wire _04182_;
 wire _04186_;
 wire _04189_;
 wire _04193_;
 wire _04196_;
 wire _04199_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04256_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04279_;
 wire _04281_;
 wire _04282_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04311_;
 wire _04313_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04377_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04400_;
 wire _04402_;
 wire _04403_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04432_;
 wire _04434_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04563_;
 wire _04567_;
 wire _04571_;
 wire _04574_;
 wire _04578_;
 wire _04581_;
 wire _04584_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04641_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04664_;
 wire _04666_;
 wire _04667_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04696_;
 wire _04698_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04762_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04785_;
 wire _04787_;
 wire _04788_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04817_;
 wire _04819_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04948_;
 wire _04952_;
 wire _04956_;
 wire _04959_;
 wire _04963_;
 wire _04966_;
 wire _04969_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05026_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05049_;
 wire _05051_;
 wire _05052_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05081_;
 wire _05083_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05147_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05170_;
 wire _05172_;
 wire _05173_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05202_;
 wire _05204_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05330_;
 wire _05331_;
 wire _05334_;
 wire _05338_;
 wire _05340_;
 wire _05343_;
 wire _05345_;
 wire _05347_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05371_;
 wire _05372_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05385_;
 wire _05389_;
 wire _05391_;
 wire _05392_;
 wire _05395_;
 wire _05397_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05442_;
 wire _05448_;
 wire _05451_;
 wire _05452_;
 wire _05456_;
 wire _05458_;
 wire _05460_;
 wire _05461_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05475_;
 wire _05476_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05486_;
 wire _05491_;
 wire _05494_;
 wire _05497_;
 wire _05500_;
 wire _05504_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05512_;
 wire _05515_;
 wire _05518_;
 wire _05519_;
 wire _05521_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05581_;
 wire _05582_;
 wire _05584_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05594_;
 wire _05595_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05617_;
 wire _05618_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05630_;
 wire _05631_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05664_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05724_;
 wire _05725_;
 wire _05727_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05737_;
 wire _05738_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05760_;
 wire _05761_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05773_;
 wire _05774_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05807_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05937_;
 wire _05942_;
 wire _05945_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05961_;
 wire _05964_;
 wire _05967_;
 wire _05970_;
 wire _05973_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06064_;
 wire _06066_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06088_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06207_;
 wire _06209_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06231_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06344_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06414_;
 wire _06417_;
 wire _06422_;
 wire _06425_;
 wire _06431_;
 wire _06434_;
 wire _06437_;
 wire _06440_;
 wire _06444_;
 wire _06447_;
 wire _06450_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06468_;
 wire _06473_;
 wire _06476_;
 wire _06480_;
 wire _06487_;
 wire _06490_;
 wire _06493_;
 wire _06496_;
 wire _06499_;
 wire _06502_;
 wire _06505_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06599_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06620_;
 wire _06622_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06650_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06674_;
 wire _06675_;
 wire _06678_;
 wire _06680_;
 wire _06682_;
 wire _06684_;
 wire _06686_;
 wire _06688_;
 wire _06690_;
 wire _06692_;
 wire _06694_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06708_;
 wire _06710_;
 wire _06712_;
 wire _06714_;
 wire _06715_;
 wire _06717_;
 wire _06719_;
 wire _06721_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06747_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06841_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06862_;
 wire _06864_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06892_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06916_;
 wire _06917_;
 wire _06920_;
 wire _06922_;
 wire _06924_;
 wire _06926_;
 wire _06928_;
 wire _06930_;
 wire _06932_;
 wire _06934_;
 wire _06936_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06950_;
 wire _06952_;
 wire _06954_;
 wire _06956_;
 wire _06957_;
 wire _06959_;
 wire _06961_;
 wire _06963_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07177_;
 wire _07182_;
 wire _07185_;
 wire _07189_;
 wire _07195_;
 wire _07198_;
 wire _07201_;
 wire _07204_;
 wire _07207_;
 wire _07210_;
 wire _07213_;
 wire _07214_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07243_;
 wire _07244_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07299_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07307_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07320_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07331_;
 wire _07332_;
 wire _07334_;
 wire _07335_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07364_;
 wire _07365_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07420_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07428_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07530_;
 wire _07532_;
 wire _07533_;
 wire _07535_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07568_;
 wire _07572_;
 wire _07576_;
 wire _07577_;
 wire _07579_;
 wire _07581_;
 wire _07583_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07590_;
 wire _07591_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07600_;
 wire _07601_;
 wire _07603_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07619_;
 wire _07620_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07659_;
 wire _07660_;
 wire _07663_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07671_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07677_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07754_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07802_;
 wire _07803_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07930_;
 wire _07933_;
 wire _07934_;
 wire _07936_;
 wire _07937_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07983_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08084_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08116_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08144_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08186_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08256_;
 wire _08257_;
 wire _08259_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08275_;
 wire _08276_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08318_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08330_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08348_;
 wire _08351_;
 wire _08352_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08364_;
 wire _08365_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08404_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08416_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08433_;
 wire _08436_;
 wire _08437_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08449_;
 wire _08450_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08481_;
 wire _08482_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08493_;
 wire _08494_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08521_;
 wire _08522_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08534_;
 wire _08535_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08573_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08585_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08654_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08666_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08700_;
 wire _08701_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08735_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08747_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08764_;
 wire _08765_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08777_;
 wire _08778_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08817_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire \count15_1[1] ;
 wire \count15_1[2] ;
 wire \count15_1[3] ;
 wire \count15_1[4] ;
 wire \count15_1[5] ;
 wire \count15_2[1] ;
 wire \count15_2[2] ;
 wire \count15_2[3] ;
 wire \count15_2[4] ;
 wire \count15_2[5] ;
 wire \count16_1[1] ;
 wire \count16_1[2] ;
 wire \count16_1[3] ;
 wire \count16_1[4] ;
 wire \count16_1[5] ;
 wire \count16_2[1] ;
 wire \count16_2[2] ;
 wire \count16_2[3] ;
 wire \count16_2[4] ;
 wire \count16_2[5] ;
 wire \count2_1[1] ;
 wire \count2_1[2] ;
 wire \count2_1[3] ;
 wire \count2_1[4] ;
 wire \count2_1[5] ;
 wire \count2_2[1] ;
 wire \count2_2[2] ;
 wire \count2_2[3] ;
 wire \count2_2[4] ;
 wire \count2_2[5] ;
 wire \count7_1[1] ;
 wire \count7_1[2] ;
 wire \count7_1[3] ;
 wire \count7_1[4] ;
 wire \count7_1[5] ;
 wire \count7_2[1] ;
 wire \count7_2[2] ;
 wire \count7_2[3] ;
 wire \count7_2[4] ;
 wire \count7_2[5] ;
 wire \count_1[1] ;
 wire \count_1[2] ;
 wire \count_1[3] ;
 wire \count_1[4] ;
 wire \count_1[5] ;
 wire \count_2[1] ;
 wire \count_2[2] ;
 wire \count_2[3] ;
 wire \count_2[4] ;
 wire \count_2[5] ;
 wire \count_2[6] ;
 wire \count_hash1[1] ;
 wire \count_hash1[2] ;
 wire \count_hash1[3] ;
 wire \count_hash1[4] ;
 wire \count_hash1[5] ;
 wire \count_hash1[6] ;
 wire \count_hash2[1] ;
 wire \count_hash2[2] ;
 wire \count_hash2[3] ;
 wire \count_hash2[4] ;
 wire \count_hash2[5] ;
 wire done;
 wire \k_value1[0] ;
 wire \k_value1[10] ;
 wire \k_value1[11] ;
 wire \k_value1[12] ;
 wire \k_value1[13] ;
 wire \k_value1[14] ;
 wire \k_value1[15] ;
 wire \k_value1[16] ;
 wire \k_value1[17] ;
 wire \k_value1[18] ;
 wire \k_value1[19] ;
 wire \k_value1[1] ;
 wire \k_value1[20] ;
 wire \k_value1[21] ;
 wire \k_value1[22] ;
 wire \k_value1[23] ;
 wire \k_value1[24] ;
 wire \k_value1[25] ;
 wire \k_value1[26] ;
 wire \k_value1[27] ;
 wire \k_value1[28] ;
 wire \k_value1[29] ;
 wire \k_value1[2] ;
 wire \k_value1[30] ;
 wire \k_value1[31] ;
 wire \k_value1[3] ;
 wire \k_value1[4] ;
 wire \k_value1[5] ;
 wire \k_value1[6] ;
 wire \k_value1[7] ;
 wire \k_value1[8] ;
 wire \k_value1[9] ;
 wire \k_value2[0] ;
 wire \k_value2[10] ;
 wire \k_value2[11] ;
 wire \k_value2[12] ;
 wire \k_value2[13] ;
 wire \k_value2[14] ;
 wire \k_value2[15] ;
 wire \k_value2[16] ;
 wire \k_value2[17] ;
 wire \k_value2[18] ;
 wire \k_value2[19] ;
 wire \k_value2[1] ;
 wire \k_value2[20] ;
 wire \k_value2[21] ;
 wire \k_value2[22] ;
 wire \k_value2[23] ;
 wire \k_value2[24] ;
 wire \k_value2[25] ;
 wire \k_value2[26] ;
 wire \k_value2[27] ;
 wire \k_value2[28] ;
 wire \k_value2[29] ;
 wire \k_value2[2] ;
 wire \k_value2[30] ;
 wire \k_value2[31] ;
 wire \k_value2[3] ;
 wire \k_value2[4] ;
 wire \k_value2[5] ;
 wire \k_value2[6] ;
 wire \k_value2[7] ;
 wire \k_value2[8] ;
 wire \k_value2[9] ;
 wire ready_dash;
 wire reset_hash;
 wire reset_hash_dash;
 wire select;
 wire \w[0][0] ;
 wire \w[0][10] ;
 wire \w[0][11] ;
 wire \w[0][12] ;
 wire \w[0][13] ;
 wire \w[0][14] ;
 wire \w[0][15] ;
 wire \w[0][16] ;
 wire \w[0][17] ;
 wire \w[0][18] ;
 wire \w[0][19] ;
 wire \w[0][1] ;
 wire \w[0][20] ;
 wire \w[0][21] ;
 wire \w[0][22] ;
 wire \w[0][23] ;
 wire \w[0][24] ;
 wire \w[0][25] ;
 wire \w[0][26] ;
 wire \w[0][27] ;
 wire \w[0][28] ;
 wire \w[0][29] ;
 wire \w[0][2] ;
 wire \w[0][30] ;
 wire \w[0][31] ;
 wire \w[0][3] ;
 wire \w[0][4] ;
 wire \w[0][5] ;
 wire \w[0][6] ;
 wire \w[0][7] ;
 wire \w[0][8] ;
 wire \w[0][9] ;
 wire \w[10][0] ;
 wire \w[10][10] ;
 wire \w[10][11] ;
 wire \w[10][12] ;
 wire \w[10][13] ;
 wire \w[10][14] ;
 wire \w[10][15] ;
 wire \w[10][16] ;
 wire \w[10][17] ;
 wire \w[10][18] ;
 wire \w[10][19] ;
 wire \w[10][1] ;
 wire \w[10][20] ;
 wire \w[10][21] ;
 wire \w[10][22] ;
 wire \w[10][23] ;
 wire \w[10][24] ;
 wire \w[10][25] ;
 wire \w[10][26] ;
 wire \w[10][27] ;
 wire \w[10][28] ;
 wire \w[10][29] ;
 wire \w[10][2] ;
 wire \w[10][30] ;
 wire \w[10][31] ;
 wire \w[10][3] ;
 wire \w[10][4] ;
 wire \w[10][5] ;
 wire \w[10][6] ;
 wire \w[10][7] ;
 wire \w[10][8] ;
 wire \w[10][9] ;
 wire \w[11][0] ;
 wire \w[11][10] ;
 wire \w[11][11] ;
 wire \w[11][12] ;
 wire \w[11][13] ;
 wire \w[11][14] ;
 wire \w[11][15] ;
 wire \w[11][16] ;
 wire \w[11][17] ;
 wire \w[11][18] ;
 wire \w[11][19] ;
 wire \w[11][1] ;
 wire \w[11][20] ;
 wire \w[11][21] ;
 wire \w[11][22] ;
 wire \w[11][23] ;
 wire \w[11][24] ;
 wire \w[11][25] ;
 wire \w[11][26] ;
 wire \w[11][27] ;
 wire \w[11][28] ;
 wire \w[11][29] ;
 wire \w[11][2] ;
 wire \w[11][30] ;
 wire \w[11][31] ;
 wire \w[11][3] ;
 wire \w[11][4] ;
 wire \w[11][5] ;
 wire \w[11][6] ;
 wire \w[11][7] ;
 wire \w[11][8] ;
 wire \w[11][9] ;
 wire \w[12][0] ;
 wire \w[12][10] ;
 wire \w[12][11] ;
 wire \w[12][12] ;
 wire \w[12][13] ;
 wire \w[12][14] ;
 wire \w[12][15] ;
 wire \w[12][16] ;
 wire \w[12][17] ;
 wire \w[12][18] ;
 wire \w[12][19] ;
 wire \w[12][1] ;
 wire \w[12][20] ;
 wire \w[12][21] ;
 wire \w[12][22] ;
 wire \w[12][23] ;
 wire \w[12][24] ;
 wire \w[12][25] ;
 wire \w[12][26] ;
 wire \w[12][27] ;
 wire \w[12][28] ;
 wire \w[12][29] ;
 wire \w[12][2] ;
 wire \w[12][30] ;
 wire \w[12][31] ;
 wire \w[12][3] ;
 wire \w[12][4] ;
 wire \w[12][5] ;
 wire \w[12][6] ;
 wire \w[12][7] ;
 wire \w[12][8] ;
 wire \w[12][9] ;
 wire \w[13][0] ;
 wire \w[13][10] ;
 wire \w[13][11] ;
 wire \w[13][12] ;
 wire \w[13][13] ;
 wire \w[13][14] ;
 wire \w[13][15] ;
 wire \w[13][16] ;
 wire \w[13][17] ;
 wire \w[13][18] ;
 wire \w[13][19] ;
 wire \w[13][1] ;
 wire \w[13][20] ;
 wire \w[13][21] ;
 wire \w[13][22] ;
 wire \w[13][23] ;
 wire \w[13][24] ;
 wire \w[13][25] ;
 wire \w[13][26] ;
 wire \w[13][27] ;
 wire \w[13][28] ;
 wire \w[13][29] ;
 wire \w[13][2] ;
 wire \w[13][30] ;
 wire \w[13][31] ;
 wire \w[13][3] ;
 wire \w[13][4] ;
 wire \w[13][5] ;
 wire \w[13][6] ;
 wire \w[13][7] ;
 wire \w[13][8] ;
 wire \w[13][9] ;
 wire \w[14][0] ;
 wire \w[14][10] ;
 wire \w[14][11] ;
 wire \w[14][12] ;
 wire \w[14][13] ;
 wire \w[14][14] ;
 wire \w[14][15] ;
 wire \w[14][16] ;
 wire \w[14][17] ;
 wire \w[14][18] ;
 wire \w[14][19] ;
 wire \w[14][1] ;
 wire \w[14][20] ;
 wire \w[14][21] ;
 wire \w[14][22] ;
 wire \w[14][23] ;
 wire \w[14][24] ;
 wire \w[14][25] ;
 wire \w[14][26] ;
 wire \w[14][27] ;
 wire \w[14][28] ;
 wire \w[14][29] ;
 wire \w[14][2] ;
 wire \w[14][30] ;
 wire \w[14][31] ;
 wire \w[14][3] ;
 wire \w[14][4] ;
 wire \w[14][5] ;
 wire \w[14][6] ;
 wire \w[14][7] ;
 wire \w[14][8] ;
 wire \w[14][9] ;
 wire \w[15][0] ;
 wire \w[15][10] ;
 wire \w[15][11] ;
 wire \w[15][12] ;
 wire \w[15][13] ;
 wire \w[15][14] ;
 wire \w[15][15] ;
 wire \w[15][16] ;
 wire \w[15][17] ;
 wire \w[15][18] ;
 wire \w[15][19] ;
 wire \w[15][1] ;
 wire \w[15][20] ;
 wire \w[15][21] ;
 wire \w[15][22] ;
 wire \w[15][23] ;
 wire \w[15][24] ;
 wire \w[15][25] ;
 wire \w[15][26] ;
 wire \w[15][27] ;
 wire \w[15][28] ;
 wire \w[15][29] ;
 wire \w[15][2] ;
 wire \w[15][30] ;
 wire \w[15][31] ;
 wire \w[15][3] ;
 wire \w[15][4] ;
 wire \w[15][5] ;
 wire \w[15][6] ;
 wire \w[15][7] ;
 wire \w[15][8] ;
 wire \w[15][9] ;
 wire \w[16][0] ;
 wire \w[16][10] ;
 wire \w[16][11] ;
 wire \w[16][12] ;
 wire \w[16][13] ;
 wire \w[16][14] ;
 wire \w[16][15] ;
 wire \w[16][16] ;
 wire \w[16][17] ;
 wire \w[16][18] ;
 wire \w[16][19] ;
 wire \w[16][1] ;
 wire \w[16][20] ;
 wire \w[16][21] ;
 wire \w[16][22] ;
 wire \w[16][23] ;
 wire \w[16][24] ;
 wire \w[16][25] ;
 wire \w[16][26] ;
 wire \w[16][27] ;
 wire \w[16][28] ;
 wire \w[16][29] ;
 wire \w[16][2] ;
 wire \w[16][30] ;
 wire \w[16][31] ;
 wire \w[16][3] ;
 wire \w[16][4] ;
 wire \w[16][5] ;
 wire \w[16][6] ;
 wire \w[16][7] ;
 wire \w[16][8] ;
 wire \w[16][9] ;
 wire \w[17][0] ;
 wire \w[17][10] ;
 wire \w[17][11] ;
 wire \w[17][12] ;
 wire \w[17][13] ;
 wire \w[17][14] ;
 wire \w[17][15] ;
 wire \w[17][16] ;
 wire \w[17][17] ;
 wire \w[17][18] ;
 wire \w[17][19] ;
 wire \w[17][1] ;
 wire \w[17][20] ;
 wire \w[17][21] ;
 wire \w[17][22] ;
 wire \w[17][23] ;
 wire \w[17][24] ;
 wire \w[17][25] ;
 wire \w[17][26] ;
 wire \w[17][27] ;
 wire \w[17][28] ;
 wire \w[17][29] ;
 wire \w[17][2] ;
 wire \w[17][30] ;
 wire \w[17][31] ;
 wire \w[17][3] ;
 wire \w[17][4] ;
 wire \w[17][5] ;
 wire \w[17][6] ;
 wire \w[17][7] ;
 wire \w[17][8] ;
 wire \w[17][9] ;
 wire \w[18][0] ;
 wire \w[18][10] ;
 wire \w[18][11] ;
 wire \w[18][12] ;
 wire \w[18][13] ;
 wire \w[18][14] ;
 wire \w[18][15] ;
 wire \w[18][16] ;
 wire \w[18][17] ;
 wire \w[18][18] ;
 wire \w[18][19] ;
 wire \w[18][1] ;
 wire \w[18][20] ;
 wire \w[18][21] ;
 wire \w[18][22] ;
 wire \w[18][23] ;
 wire \w[18][24] ;
 wire \w[18][25] ;
 wire \w[18][26] ;
 wire \w[18][27] ;
 wire \w[18][28] ;
 wire \w[18][29] ;
 wire \w[18][2] ;
 wire \w[18][30] ;
 wire \w[18][31] ;
 wire \w[18][3] ;
 wire \w[18][4] ;
 wire \w[18][5] ;
 wire \w[18][6] ;
 wire \w[18][7] ;
 wire \w[18][8] ;
 wire \w[18][9] ;
 wire \w[19][0] ;
 wire \w[19][10] ;
 wire \w[19][11] ;
 wire \w[19][12] ;
 wire \w[19][13] ;
 wire \w[19][14] ;
 wire \w[19][15] ;
 wire \w[19][16] ;
 wire \w[19][17] ;
 wire \w[19][18] ;
 wire \w[19][19] ;
 wire \w[19][1] ;
 wire \w[19][20] ;
 wire \w[19][21] ;
 wire \w[19][22] ;
 wire \w[19][23] ;
 wire \w[19][24] ;
 wire \w[19][25] ;
 wire \w[19][26] ;
 wire \w[19][27] ;
 wire \w[19][28] ;
 wire \w[19][29] ;
 wire \w[19][2] ;
 wire \w[19][30] ;
 wire \w[19][31] ;
 wire \w[19][3] ;
 wire \w[19][4] ;
 wire \w[19][5] ;
 wire \w[19][6] ;
 wire \w[19][7] ;
 wire \w[19][8] ;
 wire \w[19][9] ;
 wire \w[1][0] ;
 wire \w[1][10] ;
 wire \w[1][11] ;
 wire \w[1][12] ;
 wire \w[1][13] ;
 wire \w[1][14] ;
 wire \w[1][15] ;
 wire \w[1][16] ;
 wire \w[1][17] ;
 wire \w[1][18] ;
 wire \w[1][19] ;
 wire \w[1][1] ;
 wire \w[1][20] ;
 wire \w[1][21] ;
 wire \w[1][22] ;
 wire \w[1][23] ;
 wire \w[1][24] ;
 wire \w[1][25] ;
 wire \w[1][26] ;
 wire \w[1][27] ;
 wire \w[1][28] ;
 wire \w[1][29] ;
 wire \w[1][2] ;
 wire \w[1][30] ;
 wire \w[1][31] ;
 wire \w[1][3] ;
 wire \w[1][4] ;
 wire \w[1][5] ;
 wire \w[1][6] ;
 wire \w[1][7] ;
 wire \w[1][8] ;
 wire \w[1][9] ;
 wire \w[20][0] ;
 wire \w[20][10] ;
 wire \w[20][11] ;
 wire \w[20][12] ;
 wire \w[20][13] ;
 wire \w[20][14] ;
 wire \w[20][15] ;
 wire \w[20][16] ;
 wire \w[20][17] ;
 wire \w[20][18] ;
 wire \w[20][19] ;
 wire \w[20][1] ;
 wire \w[20][20] ;
 wire \w[20][21] ;
 wire \w[20][22] ;
 wire \w[20][23] ;
 wire \w[20][24] ;
 wire \w[20][25] ;
 wire \w[20][26] ;
 wire \w[20][27] ;
 wire \w[20][28] ;
 wire \w[20][29] ;
 wire \w[20][2] ;
 wire \w[20][30] ;
 wire \w[20][31] ;
 wire \w[20][3] ;
 wire \w[20][4] ;
 wire \w[20][5] ;
 wire \w[20][6] ;
 wire \w[20][7] ;
 wire \w[20][8] ;
 wire \w[20][9] ;
 wire \w[21][0] ;
 wire \w[21][10] ;
 wire \w[21][11] ;
 wire \w[21][12] ;
 wire \w[21][13] ;
 wire \w[21][14] ;
 wire \w[21][15] ;
 wire \w[21][16] ;
 wire \w[21][17] ;
 wire \w[21][18] ;
 wire \w[21][19] ;
 wire \w[21][1] ;
 wire \w[21][20] ;
 wire \w[21][21] ;
 wire \w[21][22] ;
 wire \w[21][23] ;
 wire \w[21][24] ;
 wire \w[21][25] ;
 wire \w[21][26] ;
 wire \w[21][27] ;
 wire \w[21][28] ;
 wire \w[21][29] ;
 wire \w[21][2] ;
 wire \w[21][30] ;
 wire \w[21][31] ;
 wire \w[21][3] ;
 wire \w[21][4] ;
 wire \w[21][5] ;
 wire \w[21][6] ;
 wire \w[21][7] ;
 wire \w[21][8] ;
 wire \w[21][9] ;
 wire \w[22][0] ;
 wire \w[22][10] ;
 wire \w[22][11] ;
 wire \w[22][12] ;
 wire \w[22][13] ;
 wire \w[22][14] ;
 wire \w[22][15] ;
 wire \w[22][16] ;
 wire \w[22][17] ;
 wire \w[22][18] ;
 wire \w[22][19] ;
 wire \w[22][1] ;
 wire \w[22][20] ;
 wire \w[22][21] ;
 wire \w[22][22] ;
 wire \w[22][23] ;
 wire \w[22][24] ;
 wire \w[22][25] ;
 wire \w[22][26] ;
 wire \w[22][27] ;
 wire \w[22][28] ;
 wire \w[22][29] ;
 wire \w[22][2] ;
 wire \w[22][30] ;
 wire \w[22][31] ;
 wire \w[22][3] ;
 wire \w[22][4] ;
 wire \w[22][5] ;
 wire \w[22][6] ;
 wire \w[22][7] ;
 wire \w[22][8] ;
 wire \w[22][9] ;
 wire \w[23][0] ;
 wire \w[23][10] ;
 wire \w[23][11] ;
 wire \w[23][12] ;
 wire \w[23][13] ;
 wire \w[23][14] ;
 wire \w[23][15] ;
 wire \w[23][16] ;
 wire \w[23][17] ;
 wire \w[23][18] ;
 wire \w[23][19] ;
 wire \w[23][1] ;
 wire \w[23][20] ;
 wire \w[23][21] ;
 wire \w[23][22] ;
 wire \w[23][23] ;
 wire \w[23][24] ;
 wire \w[23][25] ;
 wire \w[23][26] ;
 wire \w[23][27] ;
 wire \w[23][28] ;
 wire \w[23][29] ;
 wire \w[23][2] ;
 wire \w[23][30] ;
 wire \w[23][31] ;
 wire \w[23][3] ;
 wire \w[23][4] ;
 wire \w[23][5] ;
 wire \w[23][6] ;
 wire \w[23][7] ;
 wire \w[23][8] ;
 wire \w[23][9] ;
 wire \w[24][0] ;
 wire \w[24][10] ;
 wire \w[24][11] ;
 wire \w[24][12] ;
 wire \w[24][13] ;
 wire \w[24][14] ;
 wire \w[24][15] ;
 wire \w[24][16] ;
 wire \w[24][17] ;
 wire \w[24][18] ;
 wire \w[24][19] ;
 wire \w[24][1] ;
 wire \w[24][20] ;
 wire \w[24][21] ;
 wire \w[24][22] ;
 wire \w[24][23] ;
 wire \w[24][24] ;
 wire \w[24][25] ;
 wire \w[24][26] ;
 wire \w[24][27] ;
 wire \w[24][28] ;
 wire \w[24][29] ;
 wire \w[24][2] ;
 wire \w[24][30] ;
 wire \w[24][31] ;
 wire \w[24][3] ;
 wire \w[24][4] ;
 wire \w[24][5] ;
 wire \w[24][6] ;
 wire \w[24][7] ;
 wire \w[24][8] ;
 wire \w[24][9] ;
 wire \w[25][0] ;
 wire \w[25][10] ;
 wire \w[25][11] ;
 wire \w[25][12] ;
 wire \w[25][13] ;
 wire \w[25][14] ;
 wire \w[25][15] ;
 wire \w[25][16] ;
 wire \w[25][17] ;
 wire \w[25][18] ;
 wire \w[25][19] ;
 wire \w[25][1] ;
 wire \w[25][20] ;
 wire \w[25][21] ;
 wire \w[25][22] ;
 wire \w[25][23] ;
 wire \w[25][24] ;
 wire \w[25][25] ;
 wire \w[25][26] ;
 wire \w[25][27] ;
 wire \w[25][28] ;
 wire \w[25][29] ;
 wire \w[25][2] ;
 wire \w[25][30] ;
 wire \w[25][31] ;
 wire \w[25][3] ;
 wire \w[25][4] ;
 wire \w[25][5] ;
 wire \w[25][6] ;
 wire \w[25][7] ;
 wire \w[25][8] ;
 wire \w[25][9] ;
 wire \w[26][0] ;
 wire \w[26][10] ;
 wire \w[26][11] ;
 wire \w[26][12] ;
 wire \w[26][13] ;
 wire \w[26][14] ;
 wire \w[26][15] ;
 wire \w[26][16] ;
 wire \w[26][17] ;
 wire \w[26][18] ;
 wire \w[26][19] ;
 wire \w[26][1] ;
 wire \w[26][20] ;
 wire \w[26][21] ;
 wire \w[26][22] ;
 wire \w[26][23] ;
 wire \w[26][24] ;
 wire \w[26][25] ;
 wire \w[26][26] ;
 wire \w[26][27] ;
 wire \w[26][28] ;
 wire \w[26][29] ;
 wire \w[26][2] ;
 wire \w[26][30] ;
 wire \w[26][31] ;
 wire \w[26][3] ;
 wire \w[26][4] ;
 wire \w[26][5] ;
 wire \w[26][6] ;
 wire \w[26][7] ;
 wire \w[26][8] ;
 wire \w[26][9] ;
 wire \w[27][0] ;
 wire \w[27][10] ;
 wire \w[27][11] ;
 wire \w[27][12] ;
 wire \w[27][13] ;
 wire \w[27][14] ;
 wire \w[27][15] ;
 wire \w[27][16] ;
 wire \w[27][17] ;
 wire \w[27][18] ;
 wire \w[27][19] ;
 wire \w[27][1] ;
 wire \w[27][20] ;
 wire \w[27][21] ;
 wire \w[27][22] ;
 wire \w[27][23] ;
 wire \w[27][24] ;
 wire \w[27][25] ;
 wire \w[27][26] ;
 wire \w[27][27] ;
 wire \w[27][28] ;
 wire \w[27][29] ;
 wire \w[27][2] ;
 wire \w[27][30] ;
 wire \w[27][31] ;
 wire \w[27][3] ;
 wire \w[27][4] ;
 wire \w[27][5] ;
 wire \w[27][6] ;
 wire \w[27][7] ;
 wire \w[27][8] ;
 wire \w[27][9] ;
 wire \w[28][0] ;
 wire \w[28][10] ;
 wire \w[28][11] ;
 wire \w[28][12] ;
 wire \w[28][13] ;
 wire \w[28][14] ;
 wire \w[28][15] ;
 wire \w[28][16] ;
 wire \w[28][17] ;
 wire \w[28][18] ;
 wire \w[28][19] ;
 wire \w[28][1] ;
 wire \w[28][20] ;
 wire \w[28][21] ;
 wire \w[28][22] ;
 wire \w[28][23] ;
 wire \w[28][24] ;
 wire \w[28][25] ;
 wire \w[28][26] ;
 wire \w[28][27] ;
 wire \w[28][28] ;
 wire \w[28][29] ;
 wire \w[28][2] ;
 wire \w[28][30] ;
 wire \w[28][31] ;
 wire \w[28][3] ;
 wire \w[28][4] ;
 wire \w[28][5] ;
 wire \w[28][6] ;
 wire \w[28][7] ;
 wire \w[28][8] ;
 wire \w[28][9] ;
 wire \w[29][0] ;
 wire \w[29][10] ;
 wire \w[29][11] ;
 wire \w[29][12] ;
 wire \w[29][13] ;
 wire \w[29][14] ;
 wire \w[29][15] ;
 wire \w[29][16] ;
 wire \w[29][17] ;
 wire \w[29][18] ;
 wire \w[29][19] ;
 wire \w[29][1] ;
 wire \w[29][20] ;
 wire \w[29][21] ;
 wire \w[29][22] ;
 wire \w[29][23] ;
 wire \w[29][24] ;
 wire \w[29][25] ;
 wire \w[29][26] ;
 wire \w[29][27] ;
 wire \w[29][28] ;
 wire \w[29][29] ;
 wire \w[29][2] ;
 wire \w[29][30] ;
 wire \w[29][31] ;
 wire \w[29][3] ;
 wire \w[29][4] ;
 wire \w[29][5] ;
 wire \w[29][6] ;
 wire \w[29][7] ;
 wire \w[29][8] ;
 wire \w[29][9] ;
 wire \w[2][0] ;
 wire \w[2][10] ;
 wire \w[2][11] ;
 wire \w[2][12] ;
 wire \w[2][13] ;
 wire \w[2][14] ;
 wire \w[2][15] ;
 wire \w[2][16] ;
 wire \w[2][17] ;
 wire \w[2][18] ;
 wire \w[2][19] ;
 wire \w[2][1] ;
 wire \w[2][20] ;
 wire \w[2][21] ;
 wire \w[2][22] ;
 wire \w[2][23] ;
 wire \w[2][24] ;
 wire \w[2][25] ;
 wire \w[2][26] ;
 wire \w[2][27] ;
 wire \w[2][28] ;
 wire \w[2][29] ;
 wire \w[2][2] ;
 wire \w[2][30] ;
 wire \w[2][31] ;
 wire \w[2][3] ;
 wire \w[2][4] ;
 wire \w[2][5] ;
 wire \w[2][6] ;
 wire \w[2][7] ;
 wire \w[2][8] ;
 wire \w[2][9] ;
 wire \w[30][0] ;
 wire \w[30][10] ;
 wire \w[30][11] ;
 wire \w[30][12] ;
 wire \w[30][13] ;
 wire \w[30][14] ;
 wire \w[30][15] ;
 wire \w[30][16] ;
 wire \w[30][17] ;
 wire \w[30][18] ;
 wire \w[30][19] ;
 wire \w[30][1] ;
 wire \w[30][20] ;
 wire \w[30][21] ;
 wire \w[30][22] ;
 wire \w[30][23] ;
 wire \w[30][24] ;
 wire \w[30][25] ;
 wire \w[30][26] ;
 wire \w[30][27] ;
 wire \w[30][28] ;
 wire \w[30][29] ;
 wire \w[30][2] ;
 wire \w[30][30] ;
 wire \w[30][31] ;
 wire \w[30][3] ;
 wire \w[30][4] ;
 wire \w[30][5] ;
 wire \w[30][6] ;
 wire \w[30][7] ;
 wire \w[30][8] ;
 wire \w[30][9] ;
 wire \w[31][0] ;
 wire \w[31][10] ;
 wire \w[31][11] ;
 wire \w[31][12] ;
 wire \w[31][13] ;
 wire \w[31][14] ;
 wire \w[31][15] ;
 wire \w[31][16] ;
 wire \w[31][17] ;
 wire \w[31][18] ;
 wire \w[31][19] ;
 wire \w[31][1] ;
 wire \w[31][20] ;
 wire \w[31][21] ;
 wire \w[31][22] ;
 wire \w[31][23] ;
 wire \w[31][24] ;
 wire \w[31][25] ;
 wire \w[31][26] ;
 wire \w[31][27] ;
 wire \w[31][28] ;
 wire \w[31][29] ;
 wire \w[31][2] ;
 wire \w[31][30] ;
 wire \w[31][31] ;
 wire \w[31][3] ;
 wire \w[31][4] ;
 wire \w[31][5] ;
 wire \w[31][6] ;
 wire \w[31][7] ;
 wire \w[31][8] ;
 wire \w[31][9] ;
 wire \w[32][0] ;
 wire \w[32][10] ;
 wire \w[32][11] ;
 wire \w[32][12] ;
 wire \w[32][13] ;
 wire \w[32][14] ;
 wire \w[32][15] ;
 wire \w[32][16] ;
 wire \w[32][17] ;
 wire \w[32][18] ;
 wire \w[32][19] ;
 wire \w[32][1] ;
 wire \w[32][20] ;
 wire \w[32][21] ;
 wire \w[32][22] ;
 wire \w[32][23] ;
 wire \w[32][24] ;
 wire \w[32][25] ;
 wire \w[32][26] ;
 wire \w[32][27] ;
 wire \w[32][28] ;
 wire \w[32][29] ;
 wire \w[32][2] ;
 wire \w[32][30] ;
 wire \w[32][31] ;
 wire \w[32][3] ;
 wire \w[32][4] ;
 wire \w[32][5] ;
 wire \w[32][6] ;
 wire \w[32][7] ;
 wire \w[32][8] ;
 wire \w[32][9] ;
 wire \w[33][0] ;
 wire \w[33][10] ;
 wire \w[33][11] ;
 wire \w[33][12] ;
 wire \w[33][13] ;
 wire \w[33][14] ;
 wire \w[33][15] ;
 wire \w[33][16] ;
 wire \w[33][17] ;
 wire \w[33][18] ;
 wire \w[33][19] ;
 wire \w[33][1] ;
 wire \w[33][20] ;
 wire \w[33][21] ;
 wire \w[33][22] ;
 wire \w[33][23] ;
 wire \w[33][24] ;
 wire \w[33][25] ;
 wire \w[33][26] ;
 wire \w[33][27] ;
 wire \w[33][28] ;
 wire \w[33][29] ;
 wire \w[33][2] ;
 wire \w[33][30] ;
 wire \w[33][31] ;
 wire \w[33][3] ;
 wire \w[33][4] ;
 wire \w[33][5] ;
 wire \w[33][6] ;
 wire \w[33][7] ;
 wire \w[33][8] ;
 wire \w[33][9] ;
 wire \w[34][0] ;
 wire \w[34][10] ;
 wire \w[34][11] ;
 wire \w[34][12] ;
 wire \w[34][13] ;
 wire \w[34][14] ;
 wire \w[34][15] ;
 wire \w[34][16] ;
 wire \w[34][17] ;
 wire \w[34][18] ;
 wire \w[34][19] ;
 wire \w[34][1] ;
 wire \w[34][20] ;
 wire \w[34][21] ;
 wire \w[34][22] ;
 wire \w[34][23] ;
 wire \w[34][24] ;
 wire \w[34][25] ;
 wire \w[34][26] ;
 wire \w[34][27] ;
 wire \w[34][28] ;
 wire \w[34][29] ;
 wire \w[34][2] ;
 wire \w[34][30] ;
 wire \w[34][31] ;
 wire \w[34][3] ;
 wire \w[34][4] ;
 wire \w[34][5] ;
 wire \w[34][6] ;
 wire \w[34][7] ;
 wire \w[34][8] ;
 wire \w[34][9] ;
 wire \w[35][0] ;
 wire \w[35][10] ;
 wire \w[35][11] ;
 wire \w[35][12] ;
 wire \w[35][13] ;
 wire \w[35][14] ;
 wire \w[35][15] ;
 wire \w[35][16] ;
 wire \w[35][17] ;
 wire \w[35][18] ;
 wire \w[35][19] ;
 wire \w[35][1] ;
 wire \w[35][20] ;
 wire \w[35][21] ;
 wire \w[35][22] ;
 wire \w[35][23] ;
 wire \w[35][24] ;
 wire \w[35][25] ;
 wire \w[35][26] ;
 wire \w[35][27] ;
 wire \w[35][28] ;
 wire \w[35][29] ;
 wire \w[35][2] ;
 wire \w[35][30] ;
 wire \w[35][31] ;
 wire \w[35][3] ;
 wire \w[35][4] ;
 wire \w[35][5] ;
 wire \w[35][6] ;
 wire \w[35][7] ;
 wire \w[35][8] ;
 wire \w[35][9] ;
 wire \w[36][0] ;
 wire \w[36][10] ;
 wire \w[36][11] ;
 wire \w[36][12] ;
 wire \w[36][13] ;
 wire \w[36][14] ;
 wire \w[36][15] ;
 wire \w[36][16] ;
 wire \w[36][17] ;
 wire \w[36][18] ;
 wire \w[36][19] ;
 wire \w[36][1] ;
 wire \w[36][20] ;
 wire \w[36][21] ;
 wire \w[36][22] ;
 wire \w[36][23] ;
 wire \w[36][24] ;
 wire \w[36][25] ;
 wire \w[36][26] ;
 wire \w[36][27] ;
 wire \w[36][28] ;
 wire \w[36][29] ;
 wire \w[36][2] ;
 wire \w[36][30] ;
 wire \w[36][31] ;
 wire \w[36][3] ;
 wire \w[36][4] ;
 wire \w[36][5] ;
 wire \w[36][6] ;
 wire \w[36][7] ;
 wire \w[36][8] ;
 wire \w[36][9] ;
 wire \w[37][0] ;
 wire \w[37][10] ;
 wire \w[37][11] ;
 wire \w[37][12] ;
 wire \w[37][13] ;
 wire \w[37][14] ;
 wire \w[37][15] ;
 wire \w[37][16] ;
 wire \w[37][17] ;
 wire \w[37][18] ;
 wire \w[37][19] ;
 wire \w[37][1] ;
 wire \w[37][20] ;
 wire \w[37][21] ;
 wire \w[37][22] ;
 wire \w[37][23] ;
 wire \w[37][24] ;
 wire \w[37][25] ;
 wire \w[37][26] ;
 wire \w[37][27] ;
 wire \w[37][28] ;
 wire \w[37][29] ;
 wire \w[37][2] ;
 wire \w[37][30] ;
 wire \w[37][31] ;
 wire \w[37][3] ;
 wire \w[37][4] ;
 wire \w[37][5] ;
 wire \w[37][6] ;
 wire \w[37][7] ;
 wire \w[37][8] ;
 wire \w[37][9] ;
 wire \w[38][0] ;
 wire \w[38][10] ;
 wire \w[38][11] ;
 wire \w[38][12] ;
 wire \w[38][13] ;
 wire \w[38][14] ;
 wire \w[38][15] ;
 wire \w[38][16] ;
 wire \w[38][17] ;
 wire \w[38][18] ;
 wire \w[38][19] ;
 wire \w[38][1] ;
 wire \w[38][20] ;
 wire \w[38][21] ;
 wire \w[38][22] ;
 wire \w[38][23] ;
 wire \w[38][24] ;
 wire \w[38][25] ;
 wire \w[38][26] ;
 wire \w[38][27] ;
 wire \w[38][28] ;
 wire \w[38][29] ;
 wire \w[38][2] ;
 wire \w[38][30] ;
 wire \w[38][31] ;
 wire \w[38][3] ;
 wire \w[38][4] ;
 wire \w[38][5] ;
 wire \w[38][6] ;
 wire \w[38][7] ;
 wire \w[38][8] ;
 wire \w[38][9] ;
 wire \w[39][0] ;
 wire \w[39][10] ;
 wire \w[39][11] ;
 wire \w[39][12] ;
 wire \w[39][13] ;
 wire \w[39][14] ;
 wire \w[39][15] ;
 wire \w[39][16] ;
 wire \w[39][17] ;
 wire \w[39][18] ;
 wire \w[39][19] ;
 wire \w[39][1] ;
 wire \w[39][20] ;
 wire \w[39][21] ;
 wire \w[39][22] ;
 wire \w[39][23] ;
 wire \w[39][24] ;
 wire \w[39][25] ;
 wire \w[39][26] ;
 wire \w[39][27] ;
 wire \w[39][28] ;
 wire \w[39][29] ;
 wire \w[39][2] ;
 wire \w[39][30] ;
 wire \w[39][31] ;
 wire \w[39][3] ;
 wire \w[39][4] ;
 wire \w[39][5] ;
 wire \w[39][6] ;
 wire \w[39][7] ;
 wire \w[39][8] ;
 wire \w[39][9] ;
 wire \w[3][0] ;
 wire \w[3][10] ;
 wire \w[3][11] ;
 wire \w[3][12] ;
 wire \w[3][13] ;
 wire \w[3][14] ;
 wire \w[3][15] ;
 wire \w[3][16] ;
 wire \w[3][17] ;
 wire \w[3][18] ;
 wire \w[3][19] ;
 wire \w[3][1] ;
 wire \w[3][20] ;
 wire \w[3][21] ;
 wire \w[3][22] ;
 wire \w[3][23] ;
 wire \w[3][24] ;
 wire \w[3][25] ;
 wire \w[3][26] ;
 wire \w[3][27] ;
 wire \w[3][28] ;
 wire \w[3][29] ;
 wire \w[3][2] ;
 wire \w[3][30] ;
 wire \w[3][31] ;
 wire \w[3][3] ;
 wire \w[3][4] ;
 wire \w[3][5] ;
 wire \w[3][6] ;
 wire \w[3][7] ;
 wire \w[3][8] ;
 wire \w[3][9] ;
 wire \w[40][0] ;
 wire \w[40][10] ;
 wire \w[40][11] ;
 wire \w[40][12] ;
 wire \w[40][13] ;
 wire \w[40][14] ;
 wire \w[40][15] ;
 wire \w[40][16] ;
 wire \w[40][17] ;
 wire \w[40][18] ;
 wire \w[40][19] ;
 wire \w[40][1] ;
 wire \w[40][20] ;
 wire \w[40][21] ;
 wire \w[40][22] ;
 wire \w[40][23] ;
 wire \w[40][24] ;
 wire \w[40][25] ;
 wire \w[40][26] ;
 wire \w[40][27] ;
 wire \w[40][28] ;
 wire \w[40][29] ;
 wire \w[40][2] ;
 wire \w[40][30] ;
 wire \w[40][31] ;
 wire \w[40][3] ;
 wire \w[40][4] ;
 wire \w[40][5] ;
 wire \w[40][6] ;
 wire \w[40][7] ;
 wire \w[40][8] ;
 wire \w[40][9] ;
 wire \w[41][0] ;
 wire \w[41][10] ;
 wire \w[41][11] ;
 wire \w[41][12] ;
 wire \w[41][13] ;
 wire \w[41][14] ;
 wire \w[41][15] ;
 wire \w[41][16] ;
 wire \w[41][17] ;
 wire \w[41][18] ;
 wire \w[41][19] ;
 wire \w[41][1] ;
 wire \w[41][20] ;
 wire \w[41][21] ;
 wire \w[41][22] ;
 wire \w[41][23] ;
 wire \w[41][24] ;
 wire \w[41][25] ;
 wire \w[41][26] ;
 wire \w[41][27] ;
 wire \w[41][28] ;
 wire \w[41][29] ;
 wire \w[41][2] ;
 wire \w[41][30] ;
 wire \w[41][31] ;
 wire \w[41][3] ;
 wire \w[41][4] ;
 wire \w[41][5] ;
 wire \w[41][6] ;
 wire \w[41][7] ;
 wire \w[41][8] ;
 wire \w[41][9] ;
 wire \w[42][0] ;
 wire \w[42][10] ;
 wire \w[42][11] ;
 wire \w[42][12] ;
 wire \w[42][13] ;
 wire \w[42][14] ;
 wire \w[42][15] ;
 wire \w[42][16] ;
 wire \w[42][17] ;
 wire \w[42][18] ;
 wire \w[42][19] ;
 wire \w[42][1] ;
 wire \w[42][20] ;
 wire \w[42][21] ;
 wire \w[42][22] ;
 wire \w[42][23] ;
 wire \w[42][24] ;
 wire \w[42][25] ;
 wire \w[42][26] ;
 wire \w[42][27] ;
 wire \w[42][28] ;
 wire \w[42][29] ;
 wire \w[42][2] ;
 wire \w[42][30] ;
 wire \w[42][31] ;
 wire \w[42][3] ;
 wire \w[42][4] ;
 wire \w[42][5] ;
 wire \w[42][6] ;
 wire \w[42][7] ;
 wire \w[42][8] ;
 wire \w[42][9] ;
 wire \w[43][0] ;
 wire \w[43][10] ;
 wire \w[43][11] ;
 wire \w[43][12] ;
 wire \w[43][13] ;
 wire \w[43][14] ;
 wire \w[43][15] ;
 wire \w[43][16] ;
 wire \w[43][17] ;
 wire \w[43][18] ;
 wire \w[43][19] ;
 wire \w[43][1] ;
 wire \w[43][20] ;
 wire \w[43][21] ;
 wire \w[43][22] ;
 wire \w[43][23] ;
 wire \w[43][24] ;
 wire \w[43][25] ;
 wire \w[43][26] ;
 wire \w[43][27] ;
 wire \w[43][28] ;
 wire \w[43][29] ;
 wire \w[43][2] ;
 wire \w[43][30] ;
 wire \w[43][31] ;
 wire \w[43][3] ;
 wire \w[43][4] ;
 wire \w[43][5] ;
 wire \w[43][6] ;
 wire \w[43][7] ;
 wire \w[43][8] ;
 wire \w[43][9] ;
 wire \w[44][0] ;
 wire \w[44][10] ;
 wire \w[44][11] ;
 wire \w[44][12] ;
 wire \w[44][13] ;
 wire \w[44][14] ;
 wire \w[44][15] ;
 wire \w[44][16] ;
 wire \w[44][17] ;
 wire \w[44][18] ;
 wire \w[44][19] ;
 wire \w[44][1] ;
 wire \w[44][20] ;
 wire \w[44][21] ;
 wire \w[44][22] ;
 wire \w[44][23] ;
 wire \w[44][24] ;
 wire \w[44][25] ;
 wire \w[44][26] ;
 wire \w[44][27] ;
 wire \w[44][28] ;
 wire \w[44][29] ;
 wire \w[44][2] ;
 wire \w[44][30] ;
 wire \w[44][31] ;
 wire \w[44][3] ;
 wire \w[44][4] ;
 wire \w[44][5] ;
 wire \w[44][6] ;
 wire \w[44][7] ;
 wire \w[44][8] ;
 wire \w[44][9] ;
 wire \w[45][0] ;
 wire \w[45][10] ;
 wire \w[45][11] ;
 wire \w[45][12] ;
 wire \w[45][13] ;
 wire \w[45][14] ;
 wire \w[45][15] ;
 wire \w[45][16] ;
 wire \w[45][17] ;
 wire \w[45][18] ;
 wire \w[45][19] ;
 wire \w[45][1] ;
 wire \w[45][20] ;
 wire \w[45][21] ;
 wire \w[45][22] ;
 wire \w[45][23] ;
 wire \w[45][24] ;
 wire \w[45][25] ;
 wire \w[45][26] ;
 wire \w[45][27] ;
 wire \w[45][28] ;
 wire \w[45][29] ;
 wire \w[45][2] ;
 wire \w[45][30] ;
 wire \w[45][31] ;
 wire \w[45][3] ;
 wire \w[45][4] ;
 wire \w[45][5] ;
 wire \w[45][6] ;
 wire \w[45][7] ;
 wire \w[45][8] ;
 wire \w[45][9] ;
 wire \w[46][0] ;
 wire \w[46][10] ;
 wire \w[46][11] ;
 wire \w[46][12] ;
 wire \w[46][13] ;
 wire \w[46][14] ;
 wire \w[46][15] ;
 wire \w[46][16] ;
 wire \w[46][17] ;
 wire \w[46][18] ;
 wire \w[46][19] ;
 wire \w[46][1] ;
 wire \w[46][20] ;
 wire \w[46][21] ;
 wire \w[46][22] ;
 wire \w[46][23] ;
 wire \w[46][24] ;
 wire \w[46][25] ;
 wire \w[46][26] ;
 wire \w[46][27] ;
 wire \w[46][28] ;
 wire \w[46][29] ;
 wire \w[46][2] ;
 wire \w[46][30] ;
 wire \w[46][31] ;
 wire \w[46][3] ;
 wire \w[46][4] ;
 wire \w[46][5] ;
 wire \w[46][6] ;
 wire \w[46][7] ;
 wire \w[46][8] ;
 wire \w[46][9] ;
 wire \w[47][0] ;
 wire \w[47][10] ;
 wire \w[47][11] ;
 wire \w[47][12] ;
 wire \w[47][13] ;
 wire \w[47][14] ;
 wire \w[47][15] ;
 wire \w[47][16] ;
 wire \w[47][17] ;
 wire \w[47][18] ;
 wire \w[47][19] ;
 wire \w[47][1] ;
 wire \w[47][20] ;
 wire \w[47][21] ;
 wire \w[47][22] ;
 wire \w[47][23] ;
 wire \w[47][24] ;
 wire \w[47][25] ;
 wire \w[47][26] ;
 wire \w[47][27] ;
 wire \w[47][28] ;
 wire \w[47][29] ;
 wire \w[47][2] ;
 wire \w[47][30] ;
 wire \w[47][31] ;
 wire \w[47][3] ;
 wire \w[47][4] ;
 wire \w[47][5] ;
 wire \w[47][6] ;
 wire \w[47][7] ;
 wire \w[47][8] ;
 wire \w[47][9] ;
 wire \w[48][0] ;
 wire \w[48][10] ;
 wire \w[48][11] ;
 wire \w[48][12] ;
 wire \w[48][13] ;
 wire \w[48][14] ;
 wire \w[48][15] ;
 wire \w[48][16] ;
 wire \w[48][17] ;
 wire \w[48][18] ;
 wire \w[48][19] ;
 wire \w[48][1] ;
 wire \w[48][20] ;
 wire \w[48][21] ;
 wire \w[48][22] ;
 wire \w[48][23] ;
 wire \w[48][24] ;
 wire \w[48][25] ;
 wire \w[48][26] ;
 wire \w[48][27] ;
 wire \w[48][28] ;
 wire \w[48][29] ;
 wire \w[48][2] ;
 wire \w[48][30] ;
 wire \w[48][31] ;
 wire \w[48][3] ;
 wire \w[48][4] ;
 wire \w[48][5] ;
 wire \w[48][6] ;
 wire \w[48][7] ;
 wire \w[48][8] ;
 wire \w[48][9] ;
 wire \w[49][0] ;
 wire \w[49][10] ;
 wire \w[49][11] ;
 wire \w[49][12] ;
 wire \w[49][13] ;
 wire \w[49][14] ;
 wire \w[49][15] ;
 wire \w[49][16] ;
 wire \w[49][17] ;
 wire \w[49][18] ;
 wire \w[49][19] ;
 wire \w[49][1] ;
 wire \w[49][20] ;
 wire \w[49][21] ;
 wire \w[49][22] ;
 wire \w[49][23] ;
 wire \w[49][24] ;
 wire \w[49][25] ;
 wire \w[49][26] ;
 wire \w[49][27] ;
 wire \w[49][28] ;
 wire \w[49][29] ;
 wire \w[49][2] ;
 wire \w[49][30] ;
 wire \w[49][31] ;
 wire \w[49][3] ;
 wire \w[49][4] ;
 wire \w[49][5] ;
 wire \w[49][6] ;
 wire \w[49][7] ;
 wire \w[49][8] ;
 wire \w[49][9] ;
 wire \w[4][0] ;
 wire \w[4][10] ;
 wire \w[4][11] ;
 wire \w[4][12] ;
 wire \w[4][13] ;
 wire \w[4][14] ;
 wire \w[4][15] ;
 wire \w[4][16] ;
 wire \w[4][17] ;
 wire \w[4][18] ;
 wire \w[4][19] ;
 wire \w[4][1] ;
 wire \w[4][20] ;
 wire \w[4][21] ;
 wire \w[4][22] ;
 wire \w[4][23] ;
 wire \w[4][24] ;
 wire \w[4][25] ;
 wire \w[4][26] ;
 wire \w[4][27] ;
 wire \w[4][28] ;
 wire \w[4][29] ;
 wire \w[4][2] ;
 wire \w[4][30] ;
 wire \w[4][31] ;
 wire \w[4][3] ;
 wire \w[4][4] ;
 wire \w[4][5] ;
 wire \w[4][6] ;
 wire \w[4][7] ;
 wire \w[4][8] ;
 wire \w[4][9] ;
 wire \w[50][0] ;
 wire \w[50][10] ;
 wire \w[50][11] ;
 wire \w[50][12] ;
 wire \w[50][13] ;
 wire \w[50][14] ;
 wire \w[50][15] ;
 wire \w[50][16] ;
 wire \w[50][17] ;
 wire \w[50][18] ;
 wire \w[50][19] ;
 wire \w[50][1] ;
 wire \w[50][20] ;
 wire \w[50][21] ;
 wire \w[50][22] ;
 wire \w[50][23] ;
 wire \w[50][24] ;
 wire \w[50][25] ;
 wire \w[50][26] ;
 wire \w[50][27] ;
 wire \w[50][28] ;
 wire \w[50][29] ;
 wire \w[50][2] ;
 wire \w[50][30] ;
 wire \w[50][31] ;
 wire \w[50][3] ;
 wire \w[50][4] ;
 wire \w[50][5] ;
 wire \w[50][6] ;
 wire \w[50][7] ;
 wire \w[50][8] ;
 wire \w[50][9] ;
 wire \w[51][0] ;
 wire \w[51][10] ;
 wire \w[51][11] ;
 wire \w[51][12] ;
 wire \w[51][13] ;
 wire \w[51][14] ;
 wire \w[51][15] ;
 wire \w[51][16] ;
 wire \w[51][17] ;
 wire \w[51][18] ;
 wire \w[51][19] ;
 wire \w[51][1] ;
 wire \w[51][20] ;
 wire \w[51][21] ;
 wire \w[51][22] ;
 wire \w[51][23] ;
 wire \w[51][24] ;
 wire \w[51][25] ;
 wire \w[51][26] ;
 wire \w[51][27] ;
 wire \w[51][28] ;
 wire \w[51][29] ;
 wire \w[51][2] ;
 wire \w[51][30] ;
 wire \w[51][31] ;
 wire \w[51][3] ;
 wire \w[51][4] ;
 wire \w[51][5] ;
 wire \w[51][6] ;
 wire \w[51][7] ;
 wire \w[51][8] ;
 wire \w[51][9] ;
 wire \w[52][0] ;
 wire \w[52][10] ;
 wire \w[52][11] ;
 wire \w[52][12] ;
 wire \w[52][13] ;
 wire \w[52][14] ;
 wire \w[52][15] ;
 wire \w[52][16] ;
 wire \w[52][17] ;
 wire \w[52][18] ;
 wire \w[52][19] ;
 wire \w[52][1] ;
 wire \w[52][20] ;
 wire \w[52][21] ;
 wire \w[52][22] ;
 wire \w[52][23] ;
 wire \w[52][24] ;
 wire \w[52][25] ;
 wire \w[52][26] ;
 wire \w[52][27] ;
 wire \w[52][28] ;
 wire \w[52][29] ;
 wire \w[52][2] ;
 wire \w[52][30] ;
 wire \w[52][31] ;
 wire \w[52][3] ;
 wire \w[52][4] ;
 wire \w[52][5] ;
 wire \w[52][6] ;
 wire \w[52][7] ;
 wire \w[52][8] ;
 wire \w[52][9] ;
 wire \w[53][0] ;
 wire \w[53][10] ;
 wire \w[53][11] ;
 wire \w[53][12] ;
 wire \w[53][13] ;
 wire \w[53][14] ;
 wire \w[53][15] ;
 wire \w[53][16] ;
 wire \w[53][17] ;
 wire \w[53][18] ;
 wire \w[53][19] ;
 wire \w[53][1] ;
 wire \w[53][20] ;
 wire \w[53][21] ;
 wire \w[53][22] ;
 wire \w[53][23] ;
 wire \w[53][24] ;
 wire \w[53][25] ;
 wire \w[53][26] ;
 wire \w[53][27] ;
 wire \w[53][28] ;
 wire \w[53][29] ;
 wire \w[53][2] ;
 wire \w[53][30] ;
 wire \w[53][31] ;
 wire \w[53][3] ;
 wire \w[53][4] ;
 wire \w[53][5] ;
 wire \w[53][6] ;
 wire \w[53][7] ;
 wire \w[53][8] ;
 wire \w[53][9] ;
 wire \w[54][0] ;
 wire \w[54][10] ;
 wire \w[54][11] ;
 wire \w[54][12] ;
 wire \w[54][13] ;
 wire \w[54][14] ;
 wire \w[54][15] ;
 wire \w[54][16] ;
 wire \w[54][17] ;
 wire \w[54][18] ;
 wire \w[54][19] ;
 wire \w[54][1] ;
 wire \w[54][20] ;
 wire \w[54][21] ;
 wire \w[54][22] ;
 wire \w[54][23] ;
 wire \w[54][24] ;
 wire \w[54][25] ;
 wire \w[54][26] ;
 wire \w[54][27] ;
 wire \w[54][28] ;
 wire \w[54][29] ;
 wire \w[54][2] ;
 wire \w[54][30] ;
 wire \w[54][31] ;
 wire \w[54][3] ;
 wire \w[54][4] ;
 wire \w[54][5] ;
 wire \w[54][6] ;
 wire \w[54][7] ;
 wire \w[54][8] ;
 wire \w[54][9] ;
 wire \w[55][0] ;
 wire \w[55][10] ;
 wire \w[55][11] ;
 wire \w[55][12] ;
 wire \w[55][13] ;
 wire \w[55][14] ;
 wire \w[55][15] ;
 wire \w[55][16] ;
 wire \w[55][17] ;
 wire \w[55][18] ;
 wire \w[55][19] ;
 wire \w[55][1] ;
 wire \w[55][20] ;
 wire \w[55][21] ;
 wire \w[55][22] ;
 wire \w[55][23] ;
 wire \w[55][24] ;
 wire \w[55][25] ;
 wire \w[55][26] ;
 wire \w[55][27] ;
 wire \w[55][28] ;
 wire \w[55][29] ;
 wire \w[55][2] ;
 wire \w[55][30] ;
 wire \w[55][31] ;
 wire \w[55][3] ;
 wire \w[55][4] ;
 wire \w[55][5] ;
 wire \w[55][6] ;
 wire \w[55][7] ;
 wire \w[55][8] ;
 wire \w[55][9] ;
 wire \w[56][0] ;
 wire \w[56][10] ;
 wire \w[56][11] ;
 wire \w[56][12] ;
 wire \w[56][13] ;
 wire \w[56][14] ;
 wire \w[56][15] ;
 wire \w[56][16] ;
 wire \w[56][17] ;
 wire \w[56][18] ;
 wire \w[56][19] ;
 wire \w[56][1] ;
 wire \w[56][20] ;
 wire \w[56][21] ;
 wire \w[56][22] ;
 wire \w[56][23] ;
 wire \w[56][24] ;
 wire \w[56][25] ;
 wire \w[56][26] ;
 wire \w[56][27] ;
 wire \w[56][28] ;
 wire \w[56][29] ;
 wire \w[56][2] ;
 wire \w[56][30] ;
 wire \w[56][31] ;
 wire \w[56][3] ;
 wire \w[56][4] ;
 wire \w[56][5] ;
 wire \w[56][6] ;
 wire \w[56][7] ;
 wire \w[56][8] ;
 wire \w[56][9] ;
 wire \w[57][0] ;
 wire \w[57][10] ;
 wire \w[57][11] ;
 wire \w[57][12] ;
 wire \w[57][13] ;
 wire \w[57][14] ;
 wire \w[57][15] ;
 wire \w[57][16] ;
 wire \w[57][17] ;
 wire \w[57][18] ;
 wire \w[57][19] ;
 wire \w[57][1] ;
 wire \w[57][20] ;
 wire \w[57][21] ;
 wire \w[57][22] ;
 wire \w[57][23] ;
 wire \w[57][24] ;
 wire \w[57][25] ;
 wire \w[57][26] ;
 wire \w[57][27] ;
 wire \w[57][28] ;
 wire \w[57][29] ;
 wire \w[57][2] ;
 wire \w[57][30] ;
 wire \w[57][31] ;
 wire \w[57][3] ;
 wire \w[57][4] ;
 wire \w[57][5] ;
 wire \w[57][6] ;
 wire \w[57][7] ;
 wire \w[57][8] ;
 wire \w[57][9] ;
 wire \w[58][0] ;
 wire \w[58][10] ;
 wire \w[58][11] ;
 wire \w[58][12] ;
 wire \w[58][13] ;
 wire \w[58][14] ;
 wire \w[58][15] ;
 wire \w[58][16] ;
 wire \w[58][17] ;
 wire \w[58][18] ;
 wire \w[58][19] ;
 wire \w[58][1] ;
 wire \w[58][20] ;
 wire \w[58][21] ;
 wire \w[58][22] ;
 wire \w[58][23] ;
 wire \w[58][24] ;
 wire \w[58][25] ;
 wire \w[58][26] ;
 wire \w[58][27] ;
 wire \w[58][28] ;
 wire \w[58][29] ;
 wire \w[58][2] ;
 wire \w[58][30] ;
 wire \w[58][31] ;
 wire \w[58][3] ;
 wire \w[58][4] ;
 wire \w[58][5] ;
 wire \w[58][6] ;
 wire \w[58][7] ;
 wire \w[58][8] ;
 wire \w[58][9] ;
 wire \w[59][0] ;
 wire \w[59][10] ;
 wire \w[59][11] ;
 wire \w[59][12] ;
 wire \w[59][13] ;
 wire \w[59][14] ;
 wire \w[59][15] ;
 wire \w[59][16] ;
 wire \w[59][17] ;
 wire \w[59][18] ;
 wire \w[59][19] ;
 wire \w[59][1] ;
 wire \w[59][20] ;
 wire \w[59][21] ;
 wire \w[59][22] ;
 wire \w[59][23] ;
 wire \w[59][24] ;
 wire \w[59][25] ;
 wire \w[59][26] ;
 wire \w[59][27] ;
 wire \w[59][28] ;
 wire \w[59][29] ;
 wire \w[59][2] ;
 wire \w[59][30] ;
 wire \w[59][31] ;
 wire \w[59][3] ;
 wire \w[59][4] ;
 wire \w[59][5] ;
 wire \w[59][6] ;
 wire \w[59][7] ;
 wire \w[59][8] ;
 wire \w[59][9] ;
 wire \w[5][0] ;
 wire \w[5][10] ;
 wire \w[5][11] ;
 wire \w[5][12] ;
 wire \w[5][13] ;
 wire \w[5][14] ;
 wire \w[5][15] ;
 wire \w[5][16] ;
 wire \w[5][17] ;
 wire \w[5][18] ;
 wire \w[5][19] ;
 wire \w[5][1] ;
 wire \w[5][20] ;
 wire \w[5][21] ;
 wire \w[5][22] ;
 wire \w[5][23] ;
 wire \w[5][24] ;
 wire \w[5][25] ;
 wire \w[5][26] ;
 wire \w[5][27] ;
 wire \w[5][28] ;
 wire \w[5][29] ;
 wire \w[5][2] ;
 wire \w[5][30] ;
 wire \w[5][31] ;
 wire \w[5][3] ;
 wire \w[5][4] ;
 wire \w[5][5] ;
 wire \w[5][6] ;
 wire \w[5][7] ;
 wire \w[5][8] ;
 wire \w[5][9] ;
 wire \w[60][0] ;
 wire \w[60][10] ;
 wire \w[60][11] ;
 wire \w[60][12] ;
 wire \w[60][13] ;
 wire \w[60][14] ;
 wire \w[60][15] ;
 wire \w[60][16] ;
 wire \w[60][17] ;
 wire \w[60][18] ;
 wire \w[60][19] ;
 wire \w[60][1] ;
 wire \w[60][20] ;
 wire \w[60][21] ;
 wire \w[60][22] ;
 wire \w[60][23] ;
 wire \w[60][24] ;
 wire \w[60][25] ;
 wire \w[60][26] ;
 wire \w[60][27] ;
 wire \w[60][28] ;
 wire \w[60][29] ;
 wire \w[60][2] ;
 wire \w[60][30] ;
 wire \w[60][31] ;
 wire \w[60][3] ;
 wire \w[60][4] ;
 wire \w[60][5] ;
 wire \w[60][6] ;
 wire \w[60][7] ;
 wire \w[60][8] ;
 wire \w[60][9] ;
 wire \w[61][0] ;
 wire \w[61][10] ;
 wire \w[61][11] ;
 wire \w[61][12] ;
 wire \w[61][13] ;
 wire \w[61][14] ;
 wire \w[61][15] ;
 wire \w[61][16] ;
 wire \w[61][17] ;
 wire \w[61][18] ;
 wire \w[61][19] ;
 wire \w[61][1] ;
 wire \w[61][20] ;
 wire \w[61][21] ;
 wire \w[61][22] ;
 wire \w[61][23] ;
 wire \w[61][24] ;
 wire \w[61][25] ;
 wire \w[61][26] ;
 wire \w[61][27] ;
 wire \w[61][28] ;
 wire \w[61][29] ;
 wire \w[61][2] ;
 wire \w[61][30] ;
 wire \w[61][31] ;
 wire \w[61][3] ;
 wire \w[61][4] ;
 wire \w[61][5] ;
 wire \w[61][6] ;
 wire \w[61][7] ;
 wire \w[61][8] ;
 wire \w[61][9] ;
 wire \w[62][0] ;
 wire \w[62][10] ;
 wire \w[62][11] ;
 wire \w[62][12] ;
 wire \w[62][13] ;
 wire \w[62][14] ;
 wire \w[62][15] ;
 wire \w[62][16] ;
 wire \w[62][17] ;
 wire \w[62][18] ;
 wire \w[62][19] ;
 wire \w[62][1] ;
 wire \w[62][20] ;
 wire \w[62][21] ;
 wire \w[62][22] ;
 wire \w[62][23] ;
 wire \w[62][24] ;
 wire \w[62][25] ;
 wire \w[62][26] ;
 wire \w[62][27] ;
 wire \w[62][28] ;
 wire \w[62][29] ;
 wire \w[62][2] ;
 wire \w[62][30] ;
 wire \w[62][31] ;
 wire \w[62][3] ;
 wire \w[62][4] ;
 wire \w[62][5] ;
 wire \w[62][6] ;
 wire \w[62][7] ;
 wire \w[62][8] ;
 wire \w[62][9] ;
 wire \w[63][0] ;
 wire \w[63][10] ;
 wire \w[63][11] ;
 wire \w[63][12] ;
 wire \w[63][13] ;
 wire \w[63][14] ;
 wire \w[63][15] ;
 wire \w[63][16] ;
 wire \w[63][17] ;
 wire \w[63][18] ;
 wire \w[63][19] ;
 wire \w[63][1] ;
 wire \w[63][20] ;
 wire \w[63][21] ;
 wire \w[63][22] ;
 wire \w[63][23] ;
 wire \w[63][24] ;
 wire \w[63][25] ;
 wire \w[63][26] ;
 wire \w[63][27] ;
 wire \w[63][28] ;
 wire \w[63][29] ;
 wire \w[63][2] ;
 wire \w[63][30] ;
 wire \w[63][31] ;
 wire \w[63][3] ;
 wire \w[63][4] ;
 wire \w[63][5] ;
 wire \w[63][6] ;
 wire \w[63][7] ;
 wire \w[63][8] ;
 wire \w[63][9] ;
 wire \w[6][0] ;
 wire \w[6][10] ;
 wire \w[6][11] ;
 wire \w[6][12] ;
 wire \w[6][13] ;
 wire \w[6][14] ;
 wire \w[6][15] ;
 wire \w[6][16] ;
 wire \w[6][17] ;
 wire \w[6][18] ;
 wire \w[6][19] ;
 wire \w[6][1] ;
 wire \w[6][20] ;
 wire \w[6][21] ;
 wire \w[6][22] ;
 wire \w[6][23] ;
 wire \w[6][24] ;
 wire \w[6][25] ;
 wire \w[6][26] ;
 wire \w[6][27] ;
 wire \w[6][28] ;
 wire \w[6][29] ;
 wire \w[6][2] ;
 wire \w[6][30] ;
 wire \w[6][31] ;
 wire \w[6][3] ;
 wire \w[6][4] ;
 wire \w[6][5] ;
 wire \w[6][6] ;
 wire \w[6][7] ;
 wire \w[6][8] ;
 wire \w[6][9] ;
 wire \w[7][0] ;
 wire \w[7][10] ;
 wire \w[7][11] ;
 wire \w[7][12] ;
 wire \w[7][13] ;
 wire \w[7][14] ;
 wire \w[7][15] ;
 wire \w[7][16] ;
 wire \w[7][17] ;
 wire \w[7][18] ;
 wire \w[7][19] ;
 wire \w[7][1] ;
 wire \w[7][20] ;
 wire \w[7][21] ;
 wire \w[7][22] ;
 wire \w[7][23] ;
 wire \w[7][24] ;
 wire \w[7][25] ;
 wire \w[7][26] ;
 wire \w[7][27] ;
 wire \w[7][28] ;
 wire \w[7][29] ;
 wire \w[7][2] ;
 wire \w[7][30] ;
 wire \w[7][31] ;
 wire \w[7][3] ;
 wire \w[7][4] ;
 wire \w[7][5] ;
 wire \w[7][6] ;
 wire \w[7][7] ;
 wire \w[7][8] ;
 wire \w[7][9] ;
 wire \w[8][0] ;
 wire \w[8][10] ;
 wire \w[8][11] ;
 wire \w[8][12] ;
 wire \w[8][13] ;
 wire \w[8][14] ;
 wire \w[8][15] ;
 wire \w[8][16] ;
 wire \w[8][17] ;
 wire \w[8][18] ;
 wire \w[8][19] ;
 wire \w[8][1] ;
 wire \w[8][20] ;
 wire \w[8][21] ;
 wire \w[8][22] ;
 wire \w[8][23] ;
 wire \w[8][24] ;
 wire \w[8][25] ;
 wire \w[8][26] ;
 wire \w[8][27] ;
 wire \w[8][28] ;
 wire \w[8][29] ;
 wire \w[8][2] ;
 wire \w[8][30] ;
 wire \w[8][31] ;
 wire \w[8][3] ;
 wire \w[8][4] ;
 wire \w[8][5] ;
 wire \w[8][6] ;
 wire \w[8][7] ;
 wire \w[8][8] ;
 wire \w[8][9] ;
 wire \w[9][0] ;
 wire \w[9][10] ;
 wire \w[9][11] ;
 wire \w[9][12] ;
 wire \w[9][13] ;
 wire \w[9][14] ;
 wire \w[9][15] ;
 wire \w[9][16] ;
 wire \w[9][17] ;
 wire \w[9][18] ;
 wire \w[9][19] ;
 wire \w[9][1] ;
 wire \w[9][20] ;
 wire \w[9][21] ;
 wire \w[9][22] ;
 wire \w[9][23] ;
 wire \w[9][24] ;
 wire \w[9][25] ;
 wire \w[9][26] ;
 wire \w[9][27] ;
 wire \w[9][28] ;
 wire \w[9][29] ;
 wire \w[9][2] ;
 wire \w[9][30] ;
 wire \w[9][31] ;
 wire \w[9][3] ;
 wire \w[9][4] ;
 wire \w[9][5] ;
 wire \w[9][6] ;
 wire \w[9][7] ;
 wire \w[9][8] ;
 wire \w[9][9] ;
 wire \w_new_calc1.temp1[0] ;
 wire \w_new_calc1.temp1[10] ;
 wire \w_new_calc1.temp1[11] ;
 wire \w_new_calc1.temp1[12] ;
 wire \w_new_calc1.temp1[13] ;
 wire \w_new_calc1.temp1[14] ;
 wire \w_new_calc1.temp1[15] ;
 wire \w_new_calc1.temp1[16] ;
 wire \w_new_calc1.temp1[17] ;
 wire \w_new_calc1.temp1[18] ;
 wire \w_new_calc1.temp1[19] ;
 wire \w_new_calc1.temp1[1] ;
 wire \w_new_calc1.temp1[20] ;
 wire \w_new_calc1.temp1[21] ;
 wire \w_new_calc1.temp1[22] ;
 wire \w_new_calc1.temp1[23] ;
 wire \w_new_calc1.temp1[24] ;
 wire \w_new_calc1.temp1[25] ;
 wire \w_new_calc1.temp1[26] ;
 wire \w_new_calc1.temp1[27] ;
 wire \w_new_calc1.temp1[28] ;
 wire \w_new_calc1.temp1[29] ;
 wire \w_new_calc1.temp1[2] ;
 wire \w_new_calc1.temp1[30] ;
 wire \w_new_calc1.temp1[31] ;
 wire \w_new_calc1.temp1[3] ;
 wire \w_new_calc1.temp1[4] ;
 wire \w_new_calc1.temp1[5] ;
 wire \w_new_calc1.temp1[6] ;
 wire \w_new_calc1.temp1[7] ;
 wire \w_new_calc1.temp1[8] ;
 wire \w_new_calc1.temp1[9] ;
 wire \w_new_calc1.temp2[0] ;
 wire \w_new_calc1.temp2[10] ;
 wire \w_new_calc1.temp2[11] ;
 wire \w_new_calc1.temp2[12] ;
 wire \w_new_calc1.temp2[13] ;
 wire \w_new_calc1.temp2[14] ;
 wire \w_new_calc1.temp2[15] ;
 wire \w_new_calc1.temp2[16] ;
 wire \w_new_calc1.temp2[17] ;
 wire \w_new_calc1.temp2[18] ;
 wire \w_new_calc1.temp2[19] ;
 wire \w_new_calc1.temp2[1] ;
 wire \w_new_calc1.temp2[20] ;
 wire \w_new_calc1.temp2[21] ;
 wire \w_new_calc1.temp2[22] ;
 wire \w_new_calc1.temp2[23] ;
 wire \w_new_calc1.temp2[24] ;
 wire \w_new_calc1.temp2[25] ;
 wire \w_new_calc1.temp2[26] ;
 wire \w_new_calc1.temp2[27] ;
 wire \w_new_calc1.temp2[28] ;
 wire \w_new_calc1.temp2[29] ;
 wire \w_new_calc1.temp2[2] ;
 wire \w_new_calc1.temp2[30] ;
 wire \w_new_calc1.temp2[31] ;
 wire \w_new_calc1.temp2[3] ;
 wire \w_new_calc1.temp2[4] ;
 wire \w_new_calc1.temp2[5] ;
 wire \w_new_calc1.temp2[6] ;
 wire \w_new_calc1.temp2[7] ;
 wire \w_new_calc1.temp2[8] ;
 wire \w_new_calc1.temp2[9] ;
 wire \w_new_calc1.w_15[0] ;
 wire \w_new_calc1.w_15[10] ;
 wire \w_new_calc1.w_15[11] ;
 wire \w_new_calc1.w_15[12] ;
 wire \w_new_calc1.w_15[13] ;
 wire \w_new_calc1.w_15[14] ;
 wire \w_new_calc1.w_15[15] ;
 wire \w_new_calc1.w_15[16] ;
 wire \w_new_calc1.w_15[17] ;
 wire \w_new_calc1.w_15[18] ;
 wire \w_new_calc1.w_15[19] ;
 wire \w_new_calc1.w_15[1] ;
 wire \w_new_calc1.w_15[20] ;
 wire \w_new_calc1.w_15[21] ;
 wire \w_new_calc1.w_15[22] ;
 wire \w_new_calc1.w_15[23] ;
 wire \w_new_calc1.w_15[24] ;
 wire \w_new_calc1.w_15[25] ;
 wire \w_new_calc1.w_15[26] ;
 wire \w_new_calc1.w_15[27] ;
 wire \w_new_calc1.w_15[28] ;
 wire \w_new_calc1.w_15[29] ;
 wire \w_new_calc1.w_15[2] ;
 wire \w_new_calc1.w_15[30] ;
 wire \w_new_calc1.w_15[31] ;
 wire \w_new_calc1.w_15[3] ;
 wire \w_new_calc1.w_15[4] ;
 wire \w_new_calc1.w_15[5] ;
 wire \w_new_calc1.w_15[6] ;
 wire \w_new_calc1.w_15[7] ;
 wire \w_new_calc1.w_15[8] ;
 wire \w_new_calc1.w_15[9] ;
 wire \w_new_calc1.w_2[0] ;
 wire \w_new_calc1.w_2[10] ;
 wire \w_new_calc1.w_2[11] ;
 wire \w_new_calc1.w_2[12] ;
 wire \w_new_calc1.w_2[13] ;
 wire \w_new_calc1.w_2[14] ;
 wire \w_new_calc1.w_2[15] ;
 wire \w_new_calc1.w_2[16] ;
 wire \w_new_calc1.w_2[17] ;
 wire \w_new_calc1.w_2[18] ;
 wire \w_new_calc1.w_2[19] ;
 wire \w_new_calc1.w_2[1] ;
 wire \w_new_calc1.w_2[20] ;
 wire \w_new_calc1.w_2[21] ;
 wire \w_new_calc1.w_2[22] ;
 wire \w_new_calc1.w_2[23] ;
 wire \w_new_calc1.w_2[24] ;
 wire \w_new_calc1.w_2[25] ;
 wire \w_new_calc1.w_2[26] ;
 wire \w_new_calc1.w_2[27] ;
 wire \w_new_calc1.w_2[28] ;
 wire \w_new_calc1.w_2[29] ;
 wire \w_new_calc1.w_2[2] ;
 wire \w_new_calc1.w_2[30] ;
 wire \w_new_calc1.w_2[31] ;
 wire \w_new_calc1.w_2[3] ;
 wire \w_new_calc1.w_2[4] ;
 wire \w_new_calc1.w_2[5] ;
 wire \w_new_calc1.w_2[6] ;
 wire \w_new_calc1.w_2[7] ;
 wire \w_new_calc1.w_2[8] ;
 wire \w_new_calc1.w_2[9] ;
 wire \w_new_calc2.temp1[0] ;
 wire \w_new_calc2.temp1[10] ;
 wire \w_new_calc2.temp1[11] ;
 wire \w_new_calc2.temp1[12] ;
 wire \w_new_calc2.temp1[13] ;
 wire \w_new_calc2.temp1[14] ;
 wire \w_new_calc2.temp1[15] ;
 wire \w_new_calc2.temp1[16] ;
 wire \w_new_calc2.temp1[17] ;
 wire \w_new_calc2.temp1[18] ;
 wire \w_new_calc2.temp1[19] ;
 wire \w_new_calc2.temp1[1] ;
 wire \w_new_calc2.temp1[20] ;
 wire \w_new_calc2.temp1[21] ;
 wire \w_new_calc2.temp1[22] ;
 wire \w_new_calc2.temp1[23] ;
 wire \w_new_calc2.temp1[24] ;
 wire \w_new_calc2.temp1[25] ;
 wire \w_new_calc2.temp1[26] ;
 wire \w_new_calc2.temp1[27] ;
 wire \w_new_calc2.temp1[28] ;
 wire \w_new_calc2.temp1[29] ;
 wire \w_new_calc2.temp1[2] ;
 wire \w_new_calc2.temp1[30] ;
 wire \w_new_calc2.temp1[31] ;
 wire \w_new_calc2.temp1[3] ;
 wire \w_new_calc2.temp1[4] ;
 wire \w_new_calc2.temp1[5] ;
 wire \w_new_calc2.temp1[6] ;
 wire \w_new_calc2.temp1[7] ;
 wire \w_new_calc2.temp1[8] ;
 wire \w_new_calc2.temp1[9] ;
 wire \w_new_calc2.temp2[0] ;
 wire \w_new_calc2.temp2[10] ;
 wire \w_new_calc2.temp2[11] ;
 wire \w_new_calc2.temp2[12] ;
 wire \w_new_calc2.temp2[13] ;
 wire \w_new_calc2.temp2[14] ;
 wire \w_new_calc2.temp2[15] ;
 wire \w_new_calc2.temp2[16] ;
 wire \w_new_calc2.temp2[17] ;
 wire \w_new_calc2.temp2[18] ;
 wire \w_new_calc2.temp2[19] ;
 wire \w_new_calc2.temp2[1] ;
 wire \w_new_calc2.temp2[20] ;
 wire \w_new_calc2.temp2[21] ;
 wire \w_new_calc2.temp2[22] ;
 wire \w_new_calc2.temp2[23] ;
 wire \w_new_calc2.temp2[24] ;
 wire \w_new_calc2.temp2[25] ;
 wire \w_new_calc2.temp2[26] ;
 wire \w_new_calc2.temp2[27] ;
 wire \w_new_calc2.temp2[28] ;
 wire \w_new_calc2.temp2[29] ;
 wire \w_new_calc2.temp2[2] ;
 wire \w_new_calc2.temp2[30] ;
 wire \w_new_calc2.temp2[31] ;
 wire \w_new_calc2.temp2[3] ;
 wire \w_new_calc2.temp2[4] ;
 wire \w_new_calc2.temp2[5] ;
 wire \w_new_calc2.temp2[6] ;
 wire \w_new_calc2.temp2[7] ;
 wire \w_new_calc2.temp2[8] ;
 wire \w_new_calc2.temp2[9] ;
 wire \w_new_calc2.w_15[0] ;
 wire \w_new_calc2.w_15[10] ;
 wire \w_new_calc2.w_15[11] ;
 wire \w_new_calc2.w_15[12] ;
 wire \w_new_calc2.w_15[13] ;
 wire \w_new_calc2.w_15[14] ;
 wire \w_new_calc2.w_15[15] ;
 wire \w_new_calc2.w_15[16] ;
 wire \w_new_calc2.w_15[17] ;
 wire \w_new_calc2.w_15[18] ;
 wire \w_new_calc2.w_15[19] ;
 wire \w_new_calc2.w_15[1] ;
 wire \w_new_calc2.w_15[20] ;
 wire \w_new_calc2.w_15[21] ;
 wire \w_new_calc2.w_15[22] ;
 wire \w_new_calc2.w_15[23] ;
 wire \w_new_calc2.w_15[24] ;
 wire \w_new_calc2.w_15[25] ;
 wire \w_new_calc2.w_15[26] ;
 wire \w_new_calc2.w_15[27] ;
 wire \w_new_calc2.w_15[28] ;
 wire \w_new_calc2.w_15[29] ;
 wire \w_new_calc2.w_15[2] ;
 wire \w_new_calc2.w_15[30] ;
 wire \w_new_calc2.w_15[31] ;
 wire \w_new_calc2.w_15[3] ;
 wire \w_new_calc2.w_15[4] ;
 wire \w_new_calc2.w_15[5] ;
 wire \w_new_calc2.w_15[6] ;
 wire \w_new_calc2.w_15[7] ;
 wire \w_new_calc2.w_15[8] ;
 wire \w_new_calc2.w_15[9] ;
 wire \w_new_calc2.w_2[0] ;
 wire \w_new_calc2.w_2[10] ;
 wire \w_new_calc2.w_2[11] ;
 wire \w_new_calc2.w_2[12] ;
 wire \w_new_calc2.w_2[13] ;
 wire \w_new_calc2.w_2[14] ;
 wire \w_new_calc2.w_2[15] ;
 wire \w_new_calc2.w_2[16] ;
 wire \w_new_calc2.w_2[17] ;
 wire \w_new_calc2.w_2[18] ;
 wire \w_new_calc2.w_2[19] ;
 wire \w_new_calc2.w_2[1] ;
 wire \w_new_calc2.w_2[20] ;
 wire \w_new_calc2.w_2[21] ;
 wire \w_new_calc2.w_2[22] ;
 wire \w_new_calc2.w_2[23] ;
 wire \w_new_calc2.w_2[24] ;
 wire \w_new_calc2.w_2[25] ;
 wire \w_new_calc2.w_2[26] ;
 wire \w_new_calc2.w_2[27] ;
 wire \w_new_calc2.w_2[28] ;
 wire \w_new_calc2.w_2[29] ;
 wire \w_new_calc2.w_2[2] ;
 wire \w_new_calc2.w_2[30] ;
 wire \w_new_calc2.w_2[31] ;
 wire \w_new_calc2.w_2[3] ;
 wire \w_new_calc2.w_2[4] ;
 wire \w_new_calc2.w_2[5] ;
 wire \w_new_calc2.w_2[6] ;
 wire \w_new_calc2.w_2[7] ;
 wire \w_new_calc2.w_2[8] ;
 wire \w_new_calc2.w_2[9] ;
 wire \w_value1[0] ;
 wire \w_value1[10] ;
 wire \w_value1[11] ;
 wire \w_value1[12] ;
 wire \w_value1[13] ;
 wire \w_value1[14] ;
 wire \w_value1[15] ;
 wire \w_value1[16] ;
 wire \w_value1[17] ;
 wire \w_value1[18] ;
 wire \w_value1[19] ;
 wire \w_value1[1] ;
 wire \w_value1[20] ;
 wire \w_value1[21] ;
 wire \w_value1[22] ;
 wire \w_value1[23] ;
 wire \w_value1[24] ;
 wire \w_value1[25] ;
 wire \w_value1[26] ;
 wire \w_value1[27] ;
 wire \w_value1[28] ;
 wire \w_value1[29] ;
 wire \w_value1[2] ;
 wire \w_value1[30] ;
 wire \w_value1[31] ;
 wire \w_value1[3] ;
 wire \w_value1[4] ;
 wire \w_value1[5] ;
 wire \w_value1[6] ;
 wire \w_value1[7] ;
 wire \w_value1[8] ;
 wire \w_value1[9] ;
 wire \w_value2[0] ;
 wire \w_value2[10] ;
 wire \w_value2[11] ;
 wire \w_value2[12] ;
 wire \w_value2[13] ;
 wire \w_value2[14] ;
 wire \w_value2[15] ;
 wire \w_value2[16] ;
 wire \w_value2[17] ;
 wire \w_value2[18] ;
 wire \w_value2[19] ;
 wire \w_value2[1] ;
 wire \w_value2[20] ;
 wire \w_value2[21] ;
 wire \w_value2[22] ;
 wire \w_value2[23] ;
 wire \w_value2[24] ;
 wire \w_value2[25] ;
 wire \w_value2[26] ;
 wire \w_value2[27] ;
 wire \w_value2[28] ;
 wire \w_value2[29] ;
 wire \w_value2[2] ;
 wire \w_value2[30] ;
 wire \w_value2[31] ;
 wire \w_value2[3] ;
 wire \w_value2[4] ;
 wire \w_value2[5] ;
 wire \w_value2[6] ;
 wire \w_value2[7] ;
 wire \w_value2[8] ;
 wire \w_value2[9] ;
 wire \hash/_0000_ ;
 wire \hash/_0001_ ;
 wire \hash/_0002_ ;
 wire \hash/_0003_ ;
 wire \hash/_0004_ ;
 wire \hash/_0005_ ;
 wire \hash/_0006_ ;
 wire \hash/_0007_ ;
 wire \hash/_0008_ ;
 wire \hash/_0009_ ;
 wire \hash/_0010_ ;
 wire \hash/_0011_ ;
 wire \hash/_0012_ ;
 wire \hash/_0013_ ;
 wire \hash/_0014_ ;
 wire \hash/_0015_ ;
 wire \hash/_0016_ ;
 wire \hash/_0017_ ;
 wire \hash/_0018_ ;
 wire \hash/_0019_ ;
 wire \hash/_0020_ ;
 wire \hash/_0021_ ;
 wire \hash/_0022_ ;
 wire \hash/_0023_ ;
 wire \hash/_0024_ ;
 wire \hash/_0025_ ;
 wire \hash/_0026_ ;
 wire \hash/_0027_ ;
 wire \hash/_0028_ ;
 wire \hash/_0029_ ;
 wire \hash/_0030_ ;
 wire \hash/_0031_ ;
 wire \hash/_0032_ ;
 wire \hash/_0033_ ;
 wire \hash/_0034_ ;
 wire \hash/_0035_ ;
 wire \hash/_0036_ ;
 wire \hash/_0037_ ;
 wire \hash/_0038_ ;
 wire \hash/_0039_ ;
 wire \hash/_0040_ ;
 wire \hash/_0041_ ;
 wire \hash/_0042_ ;
 wire \hash/_0043_ ;
 wire \hash/_0044_ ;
 wire \hash/_0045_ ;
 wire \hash/_0046_ ;
 wire \hash/_0047_ ;
 wire \hash/_0048_ ;
 wire \hash/_0049_ ;
 wire \hash/_0050_ ;
 wire \hash/_0051_ ;
 wire \hash/_0052_ ;
 wire \hash/_0053_ ;
 wire \hash/_0054_ ;
 wire \hash/_0055_ ;
 wire \hash/_0056_ ;
 wire \hash/_0057_ ;
 wire \hash/_0058_ ;
 wire \hash/_0059_ ;
 wire \hash/_0060_ ;
 wire \hash/_0061_ ;
 wire \hash/_0062_ ;
 wire \hash/_0063_ ;
 wire \hash/_0064_ ;
 wire \hash/_0065_ ;
 wire \hash/_0066_ ;
 wire \hash/_0067_ ;
 wire \hash/_0068_ ;
 wire \hash/_0069_ ;
 wire \hash/_0070_ ;
 wire \hash/_0071_ ;
 wire \hash/_0072_ ;
 wire \hash/_0073_ ;
 wire \hash/_0074_ ;
 wire \hash/_0075_ ;
 wire \hash/_0076_ ;
 wire \hash/_0077_ ;
 wire \hash/_0078_ ;
 wire \hash/_0079_ ;
 wire \hash/_0080_ ;
 wire \hash/_0081_ ;
 wire \hash/_0082_ ;
 wire \hash/_0083_ ;
 wire \hash/_0084_ ;
 wire \hash/_0085_ ;
 wire \hash/_0086_ ;
 wire \hash/_0087_ ;
 wire \hash/_0088_ ;
 wire \hash/_0089_ ;
 wire \hash/_0090_ ;
 wire \hash/_0091_ ;
 wire \hash/_0092_ ;
 wire \hash/_0093_ ;
 wire \hash/_0094_ ;
 wire \hash/_0095_ ;
 wire \hash/_0096_ ;
 wire \hash/_0097_ ;
 wire \hash/_0098_ ;
 wire \hash/_0099_ ;
 wire \hash/_0100_ ;
 wire \hash/_0101_ ;
 wire \hash/_0102_ ;
 wire \hash/_0103_ ;
 wire \hash/_0104_ ;
 wire \hash/_0105_ ;
 wire \hash/_0106_ ;
 wire \hash/_0107_ ;
 wire \hash/_0108_ ;
 wire \hash/_0109_ ;
 wire \hash/_0110_ ;
 wire \hash/_0111_ ;
 wire \hash/_0112_ ;
 wire \hash/_0113_ ;
 wire \hash/_0114_ ;
 wire \hash/_0115_ ;
 wire \hash/_0116_ ;
 wire \hash/_0117_ ;
 wire \hash/_0118_ ;
 wire \hash/_0119_ ;
 wire \hash/_0120_ ;
 wire \hash/_0121_ ;
 wire \hash/_0122_ ;
 wire \hash/_0123_ ;
 wire \hash/_0124_ ;
 wire \hash/_0125_ ;
 wire \hash/_0126_ ;
 wire \hash/_0127_ ;
 wire \hash/_0128_ ;
 wire \hash/_0129_ ;
 wire \hash/_0130_ ;
 wire \hash/_0131_ ;
 wire \hash/_0132_ ;
 wire \hash/_0133_ ;
 wire \hash/_0134_ ;
 wire \hash/_0135_ ;
 wire \hash/_0136_ ;
 wire \hash/_0137_ ;
 wire \hash/_0138_ ;
 wire \hash/_0139_ ;
 wire \hash/_0140_ ;
 wire \hash/_0141_ ;
 wire \hash/_0142_ ;
 wire \hash/_0143_ ;
 wire \hash/_0144_ ;
 wire \hash/_0145_ ;
 wire \hash/_0146_ ;
 wire \hash/_0147_ ;
 wire \hash/_0148_ ;
 wire \hash/_0149_ ;
 wire \hash/_0150_ ;
 wire \hash/_0151_ ;
 wire \hash/_0152_ ;
 wire \hash/_0153_ ;
 wire \hash/_0154_ ;
 wire \hash/_0155_ ;
 wire \hash/_0156_ ;
 wire \hash/_0157_ ;
 wire \hash/_0158_ ;
 wire \hash/_0159_ ;
 wire \hash/_0160_ ;
 wire \hash/_0161_ ;
 wire \hash/_0162_ ;
 wire \hash/_0163_ ;
 wire \hash/_0164_ ;
 wire \hash/_0165_ ;
 wire \hash/_0166_ ;
 wire \hash/_0167_ ;
 wire \hash/_0168_ ;
 wire \hash/_0169_ ;
 wire \hash/_0170_ ;
 wire \hash/_0171_ ;
 wire \hash/_0172_ ;
 wire \hash/_0173_ ;
 wire \hash/_0174_ ;
 wire \hash/_0175_ ;
 wire \hash/_0176_ ;
 wire \hash/_0177_ ;
 wire \hash/_0178_ ;
 wire \hash/_0179_ ;
 wire \hash/_0180_ ;
 wire \hash/_0181_ ;
 wire \hash/_0182_ ;
 wire \hash/_0183_ ;
 wire \hash/_0184_ ;
 wire \hash/_0185_ ;
 wire \hash/_0186_ ;
 wire \hash/_0187_ ;
 wire \hash/_0188_ ;
 wire \hash/_0189_ ;
 wire \hash/_0190_ ;
 wire \hash/_0191_ ;
 wire \hash/_0192_ ;
 wire \hash/_0193_ ;
 wire \hash/_0194_ ;
 wire \hash/_0195_ ;
 wire \hash/_0196_ ;
 wire \hash/_0197_ ;
 wire \hash/_0198_ ;
 wire \hash/_0199_ ;
 wire \hash/_0200_ ;
 wire \hash/_0201_ ;
 wire \hash/_0202_ ;
 wire \hash/_0203_ ;
 wire \hash/_0204_ ;
 wire \hash/_0205_ ;
 wire \hash/_0206_ ;
 wire \hash/_0207_ ;
 wire \hash/_0208_ ;
 wire \hash/_0209_ ;
 wire \hash/_0210_ ;
 wire \hash/_0211_ ;
 wire \hash/_0212_ ;
 wire \hash/_0213_ ;
 wire \hash/_0214_ ;
 wire \hash/_0215_ ;
 wire \hash/_0216_ ;
 wire \hash/_0217_ ;
 wire \hash/_0218_ ;
 wire \hash/_0219_ ;
 wire \hash/_0220_ ;
 wire \hash/_0221_ ;
 wire \hash/_0222_ ;
 wire \hash/_0223_ ;
 wire \hash/_0224_ ;
 wire \hash/_0225_ ;
 wire \hash/_0226_ ;
 wire \hash/_0227_ ;
 wire \hash/_0228_ ;
 wire \hash/_0229_ ;
 wire \hash/_0230_ ;
 wire \hash/_0231_ ;
 wire \hash/_0232_ ;
 wire \hash/_0233_ ;
 wire \hash/_0234_ ;
 wire \hash/_0235_ ;
 wire \hash/_0236_ ;
 wire \hash/_0237_ ;
 wire \hash/_0238_ ;
 wire \hash/_0239_ ;
 wire \hash/_0240_ ;
 wire \hash/_0241_ ;
 wire \hash/_0242_ ;
 wire \hash/_0243_ ;
 wire \hash/_0244_ ;
 wire \hash/_0245_ ;
 wire \hash/_0246_ ;
 wire \hash/_0247_ ;
 wire \hash/_0248_ ;
 wire \hash/_0249_ ;
 wire \hash/_0250_ ;
 wire \hash/_0251_ ;
 wire \hash/_0252_ ;
 wire \hash/_0253_ ;
 wire \hash/_0254_ ;
 wire \hash/_0255_ ;
 wire \hash/_0256_ ;
 wire \hash/_0257_ ;
 wire \hash/_0258_ ;
 wire \hash/_0259_ ;
 wire \hash/_0260_ ;
 wire \hash/_0261_ ;
 wire \hash/_0262_ ;
 wire \hash/_0263_ ;
 wire \hash/_0264_ ;
 wire \hash/_0265_ ;
 wire \hash/_0266_ ;
 wire \hash/_0267_ ;
 wire \hash/_0268_ ;
 wire \hash/_0269_ ;
 wire \hash/_0270_ ;
 wire \hash/_0271_ ;
 wire \hash/_0272_ ;
 wire \hash/_0273_ ;
 wire \hash/_0274_ ;
 wire \hash/_0275_ ;
 wire \hash/_0276_ ;
 wire \hash/_0278_ ;
 wire \hash/_0279_ ;
 wire \hash/_0281_ ;
 wire \hash/_0282_ ;
 wire \hash/_0283_ ;
 wire \hash/_0285_ ;
 wire \hash/_0286_ ;
 wire \hash/_0287_ ;
 wire \hash/_0288_ ;
 wire \hash/_0290_ ;
 wire \hash/_0291_ ;
 wire \hash/_0292_ ;
 wire \hash/_0293_ ;
 wire \hash/_0294_ ;
 wire \hash/_0295_ ;
 wire \hash/_0296_ ;
 wire \hash/_0297_ ;
 wire \hash/_0298_ ;
 wire \hash/_0299_ ;
 wire \hash/_0300_ ;
 wire \hash/_0301_ ;
 wire \hash/_0302_ ;
 wire \hash/_0303_ ;
 wire \hash/_0304_ ;
 wire \hash/_0305_ ;
 wire \hash/_0306_ ;
 wire \hash/_0307_ ;
 wire \hash/_0308_ ;
 wire \hash/_0309_ ;
 wire \hash/_0310_ ;
 wire \hash/_0311_ ;
 wire \hash/_0312_ ;
 wire \hash/_0313_ ;
 wire \hash/_0314_ ;
 wire \hash/_0315_ ;
 wire \hash/_0316_ ;
 wire \hash/_0317_ ;
 wire \hash/_0318_ ;
 wire \hash/_0319_ ;
 wire \hash/_0320_ ;
 wire \hash/_0321_ ;
 wire \hash/_0322_ ;
 wire \hash/_0323_ ;
 wire \hash/_0324_ ;
 wire \hash/_0325_ ;
 wire \hash/_0326_ ;
 wire \hash/_0327_ ;
 wire \hash/_0328_ ;
 wire \hash/_0329_ ;
 wire \hash/_0330_ ;
 wire \hash/_0331_ ;
 wire \hash/_0332_ ;
 wire \hash/_0333_ ;
 wire \hash/_0334_ ;
 wire \hash/_0335_ ;
 wire \hash/_0336_ ;
 wire \hash/_0337_ ;
 wire \hash/_0338_ ;
 wire \hash/_0339_ ;
 wire \hash/_0340_ ;
 wire \hash/_0341_ ;
 wire \hash/_0342_ ;
 wire \hash/_0343_ ;
 wire \hash/_0344_ ;
 wire \hash/_0345_ ;
 wire \hash/_0347_ ;
 wire \hash/_0348_ ;
 wire \hash/_0349_ ;
 wire \hash/_0350_ ;
 wire \hash/_0351_ ;
 wire \hash/_0352_ ;
 wire \hash/_0353_ ;
 wire \hash/_0354_ ;
 wire \hash/_0355_ ;
 wire \hash/_0356_ ;
 wire \hash/_0357_ ;
 wire \hash/_0358_ ;
 wire \hash/_0360_ ;
 wire \hash/_0361_ ;
 wire \hash/_0362_ ;
 wire \hash/_0363_ ;
 wire \hash/_0364_ ;
 wire \hash/_0365_ ;
 wire \hash/_0366_ ;
 wire \hash/_0367_ ;
 wire \hash/_0368_ ;
 wire \hash/_0369_ ;
 wire \hash/_0370_ ;
 wire \hash/_0371_ ;
 wire \hash/_0372_ ;
 wire \hash/_0373_ ;
 wire \hash/_0376_ ;
 wire \hash/_0377_ ;
 wire \hash/_0378_ ;
 wire \hash/_0379_ ;
 wire \hash/_0380_ ;
 wire \hash/_0381_ ;
 wire \hash/_0382_ ;
 wire \hash/_0383_ ;
 wire \hash/_0384_ ;
 wire \hash/_0385_ ;
 wire \hash/_0386_ ;
 wire \hash/_0387_ ;
 wire \hash/_0388_ ;
 wire \hash/_0389_ ;
 wire \hash/_0390_ ;
 wire \hash/_0391_ ;
 wire \hash/_0392_ ;
 wire \hash/_0393_ ;
 wire \hash/_0394_ ;
 wire \hash/_0395_ ;
 wire \hash/_0396_ ;
 wire \hash/_0397_ ;
 wire \hash/_0398_ ;
 wire \hash/_0399_ ;
 wire \hash/_0400_ ;
 wire \hash/_0401_ ;
 wire \hash/_0402_ ;
 wire \hash/_0403_ ;
 wire \hash/_0404_ ;
 wire \hash/_0405_ ;
 wire \hash/_0406_ ;
 wire \hash/_0407_ ;
 wire \hash/_0408_ ;
 wire \hash/_0409_ ;
 wire \hash/_0410_ ;
 wire \hash/_0411_ ;
 wire \hash/_0412_ ;
 wire \hash/_0413_ ;
 wire \hash/_0414_ ;
 wire \hash/_0415_ ;
 wire \hash/_0416_ ;
 wire \hash/_0417_ ;
 wire \hash/_0418_ ;
 wire \hash/_0419_ ;
 wire \hash/_0420_ ;
 wire \hash/_0421_ ;
 wire \hash/_0422_ ;
 wire \hash/_0423_ ;
 wire \hash/_0424_ ;
 wire \hash/_0425_ ;
 wire \hash/_0426_ ;
 wire \hash/_0427_ ;
 wire \hash/_0428_ ;
 wire \hash/_0429_ ;
 wire \hash/_0430_ ;
 wire \hash/_0431_ ;
 wire \hash/_0432_ ;
 wire \hash/_0433_ ;
 wire \hash/_0434_ ;
 wire \hash/_0436_ ;
 wire \hash/_0437_ ;
 wire \hash/_0438_ ;
 wire \hash/_0439_ ;
 wire \hash/_0440_ ;
 wire \hash/_0441_ ;
 wire \hash/_0442_ ;
 wire \hash/_0443_ ;
 wire \hash/_0444_ ;
 wire \hash/_0445_ ;
 wire \hash/_0446_ ;
 wire \hash/_0447_ ;
 wire \hash/_0448_ ;
 wire \hash/_0449_ ;
 wire \hash/_0450_ ;
 wire \hash/_0451_ ;
 wire \hash/_0452_ ;
 wire \hash/_0453_ ;
 wire \hash/_0454_ ;
 wire \hash/_0455_ ;
 wire \hash/_0456_ ;
 wire \hash/_0457_ ;
 wire \hash/_0458_ ;
 wire \hash/_0459_ ;
 wire \hash/_0460_ ;
 wire \hash/_0461_ ;
 wire \hash/_0462_ ;
 wire \hash/_0463_ ;
 wire \hash/_0464_ ;
 wire \hash/_0465_ ;
 wire \hash/_0466_ ;
 wire \hash/_0467_ ;
 wire \hash/_0468_ ;
 wire \hash/_0469_ ;
 wire \hash/_0470_ ;
 wire \hash/_0471_ ;
 wire \hash/_0472_ ;
 wire \hash/_0473_ ;
 wire \hash/_0474_ ;
 wire \hash/_0475_ ;
 wire \hash/_0476_ ;
 wire \hash/_0477_ ;
 wire \hash/_0478_ ;
 wire \hash/_0479_ ;
 wire \hash/_0480_ ;
 wire \hash/_0481_ ;
 wire \hash/_0482_ ;
 wire \hash/_0483_ ;
 wire \hash/_0484_ ;
 wire \hash/_0485_ ;
 wire \hash/_0486_ ;
 wire \hash/_0487_ ;
 wire \hash/_0488_ ;
 wire \hash/_0489_ ;
 wire \hash/_0490_ ;
 wire \hash/_0491_ ;
 wire \hash/_0492_ ;
 wire \hash/_0493_ ;
 wire \hash/_0494_ ;
 wire \hash/_0495_ ;
 wire \hash/_0496_ ;
 wire \hash/_0497_ ;
 wire \hash/_0498_ ;
 wire \hash/_0499_ ;
 wire \hash/_0500_ ;
 wire \hash/_0501_ ;
 wire \hash/_0502_ ;
 wire \hash/_0503_ ;
 wire \hash/_0504_ ;
 wire \hash/_0505_ ;
 wire \hash/_0506_ ;
 wire \hash/_0507_ ;
 wire \hash/_0508_ ;
 wire \hash/_0509_ ;
 wire \hash/_0510_ ;
 wire \hash/_0511_ ;
 wire \hash/_0512_ ;
 wire \hash/_0513_ ;
 wire \hash/_0514_ ;
 wire \hash/_0515_ ;
 wire \hash/_0516_ ;
 wire \hash/_0517_ ;
 wire \hash/_0518_ ;
 wire \hash/_0519_ ;
 wire \hash/_0520_ ;
 wire \hash/_0521_ ;
 wire \hash/_0522_ ;
 wire \hash/_0523_ ;
 wire \hash/_0524_ ;
 wire \hash/_0525_ ;
 wire \hash/_0526_ ;
 wire \hash/_0527_ ;
 wire \hash/_0528_ ;
 wire \hash/_0529_ ;
 wire \hash/_0530_ ;
 wire \hash/_0531_ ;
 wire \hash/_0532_ ;
 wire \hash/_0533_ ;
 wire \hash/_0534_ ;
 wire \hash/_0535_ ;
 wire \hash/_0536_ ;
 wire \hash/_0537_ ;
 wire \hash/_0538_ ;
 wire \hash/_0539_ ;
 wire \hash/_0540_ ;
 wire \hash/_0541_ ;
 wire \hash/_0542_ ;
 wire \hash/_0543_ ;
 wire \hash/_0544_ ;
 wire \hash/_0545_ ;
 wire \hash/_0546_ ;
 wire \hash/_0547_ ;
 wire \hash/_0548_ ;
 wire \hash/_0549_ ;
 wire \hash/_0550_ ;
 wire \hash/_0551_ ;
 wire \hash/_0552_ ;
 wire \hash/_0553_ ;
 wire \hash/_0554_ ;
 wire \hash/_0555_ ;
 wire \hash/_0556_ ;
 wire \hash/_0557_ ;
 wire \hash/_0558_ ;
 wire \hash/_0559_ ;
 wire \hash/_0560_ ;
 wire \hash/_0561_ ;
 wire \hash/_0562_ ;
 wire \hash/_0563_ ;
 wire \hash/_0564_ ;
 wire \hash/_0565_ ;
 wire \hash/_0567_ ;
 wire \hash/_0568_ ;
 wire \hash/_0569_ ;
 wire \hash/_0570_ ;
 wire \hash/_0571_ ;
 wire \hash/_0572_ ;
 wire \hash/_0574_ ;
 wire \hash/_0575_ ;
 wire \hash/_0576_ ;
 wire \hash/_0577_ ;
 wire \hash/_0578_ ;
 wire \hash/_0579_ ;
 wire \hash/_0580_ ;
 wire \hash/_0581_ ;
 wire \hash/_0582_ ;
 wire \hash/_0583_ ;
 wire \hash/_0584_ ;
 wire \hash/_0585_ ;
 wire \hash/_0586_ ;
 wire \hash/_0587_ ;
 wire \hash/_0589_ ;
 wire \hash/_0590_ ;
 wire \hash/_0591_ ;
 wire \hash/_0592_ ;
 wire \hash/_0593_ ;
 wire \hash/_0594_ ;
 wire \hash/_0595_ ;
 wire \hash/_0596_ ;
 wire \hash/_0597_ ;
 wire \hash/_0598_ ;
 wire \hash/_0599_ ;
 wire \hash/_0600_ ;
 wire \hash/_0601_ ;
 wire \hash/_0602_ ;
 wire \hash/_0603_ ;
 wire \hash/_0604_ ;
 wire \hash/_0605_ ;
 wire \hash/_0606_ ;
 wire \hash/_0607_ ;
 wire \hash/_0608_ ;
 wire \hash/_0609_ ;
 wire \hash/_0610_ ;
 wire \hash/_0611_ ;
 wire \hash/_0612_ ;
 wire \hash/_0613_ ;
 wire \hash/_0614_ ;
 wire \hash/_0615_ ;
 wire \hash/_0616_ ;
 wire \hash/_0617_ ;
 wire \hash/_0618_ ;
 wire \hash/_0619_ ;
 wire \hash/_0620_ ;
 wire \hash/_0621_ ;
 wire \hash/_0622_ ;
 wire \hash/_0623_ ;
 wire \hash/_0624_ ;
 wire \hash/_0625_ ;
 wire \hash/_0626_ ;
 wire \hash/_0627_ ;
 wire \hash/_0628_ ;
 wire \hash/_0629_ ;
 wire \hash/_0630_ ;
 wire \hash/_0631_ ;
 wire \hash/_0632_ ;
 wire \hash/_0633_ ;
 wire \hash/_0634_ ;
 wire \hash/_0635_ ;
 wire \hash/_0636_ ;
 wire \hash/_0637_ ;
 wire \hash/_0638_ ;
 wire \hash/_0639_ ;
 wire \hash/_0640_ ;
 wire \hash/_0641_ ;
 wire \hash/_0642_ ;
 wire \hash/_0643_ ;
 wire \hash/_0644_ ;
 wire \hash/_0645_ ;
 wire \hash/_0646_ ;
 wire \hash/_0647_ ;
 wire \hash/_0648_ ;
 wire \hash/_0649_ ;
 wire \hash/_0650_ ;
 wire \hash/_0651_ ;
 wire \hash/_0652_ ;
 wire \hash/_0653_ ;
 wire \hash/_0654_ ;
 wire \hash/_0655_ ;
 wire \hash/_0656_ ;
 wire \hash/_0657_ ;
 wire \hash/_0658_ ;
 wire \hash/_0659_ ;
 wire \hash/_0660_ ;
 wire \hash/_0661_ ;
 wire \hash/_0662_ ;
 wire \hash/_0664_ ;
 wire \hash/_0665_ ;
 wire \hash/_0666_ ;
 wire \hash/_0667_ ;
 wire \hash/_0668_ ;
 wire \hash/_0669_ ;
 wire \hash/_0670_ ;
 wire \hash/_0671_ ;
 wire \hash/_0672_ ;
 wire \hash/_0673_ ;
 wire \hash/_0674_ ;
 wire \hash/_0675_ ;
 wire \hash/_0676_ ;
 wire \hash/_0677_ ;
 wire \hash/_0679_ ;
 wire \hash/_0680_ ;
 wire \hash/_0681_ ;
 wire \hash/_0682_ ;
 wire \hash/_0683_ ;
 wire \hash/_0684_ ;
 wire \hash/_0685_ ;
 wire \hash/_0686_ ;
 wire \hash/_0687_ ;
 wire \hash/_0688_ ;
 wire \hash/_0689_ ;
 wire \hash/_0690_ ;
 wire \hash/_0691_ ;
 wire \hash/_0692_ ;
 wire \hash/_0693_ ;
 wire \hash/_0694_ ;
 wire \hash/_0695_ ;
 wire \hash/_0696_ ;
 wire \hash/_0697_ ;
 wire \hash/_0698_ ;
 wire \hash/_0699_ ;
 wire \hash/_0700_ ;
 wire \hash/_0701_ ;
 wire \hash/_0702_ ;
 wire \hash/_0703_ ;
 wire \hash/_0704_ ;
 wire \hash/_0705_ ;
 wire \hash/_0706_ ;
 wire \hash/_0707_ ;
 wire \hash/_0708_ ;
 wire \hash/_0709_ ;
 wire \hash/_0710_ ;
 wire \hash/_0711_ ;
 wire \hash/_0712_ ;
 wire \hash/_0713_ ;
 wire \hash/_0714_ ;
 wire \hash/_0715_ ;
 wire \hash/_0716_ ;
 wire \hash/_0717_ ;
 wire \hash/_0718_ ;
 wire \hash/_0719_ ;
 wire \hash/_0720_ ;
 wire \hash/_0721_ ;
 wire \hash/_0722_ ;
 wire \hash/_0723_ ;
 wire \hash/_0724_ ;
 wire \hash/_0725_ ;
 wire \hash/_0726_ ;
 wire \hash/_0727_ ;
 wire \hash/_0728_ ;
 wire \hash/_0729_ ;
 wire \hash/_0730_ ;
 wire \hash/_0731_ ;
 wire \hash/_0732_ ;
 wire \hash/_0733_ ;
 wire \hash/_0734_ ;
 wire \hash/_0735_ ;
 wire \hash/_0736_ ;
 wire \hash/_0737_ ;
 wire \hash/_0738_ ;
 wire \hash/_0739_ ;
 wire \hash/_0740_ ;
 wire \hash/_0741_ ;
 wire \hash/_0742_ ;
 wire \hash/_0743_ ;
 wire \hash/_0744_ ;
 wire \hash/_0745_ ;
 wire \hash/_0746_ ;
 wire \hash/_0747_ ;
 wire \hash/_0748_ ;
 wire \hash/_0749_ ;
 wire \hash/_0750_ ;
 wire \hash/_0751_ ;
 wire \hash/_0752_ ;
 wire \hash/_0753_ ;
 wire \hash/_0754_ ;
 wire \hash/_0755_ ;
 wire \hash/_0756_ ;
 wire \hash/_0757_ ;
 wire \hash/_0758_ ;
 wire \hash/_0759_ ;
 wire \hash/_0760_ ;
 wire \hash/_0761_ ;
 wire \hash/_0762_ ;
 wire \hash/_0763_ ;
 wire \hash/_0764_ ;
 wire \hash/_0765_ ;
 wire \hash/_0766_ ;
 wire \hash/_0767_ ;
 wire \hash/_0768_ ;
 wire \hash/_0769_ ;
 wire \hash/_0770_ ;
 wire \hash/_0771_ ;
 wire \hash/_0772_ ;
 wire \hash/_0774_ ;
 wire \hash/_0775_ ;
 wire \hash/_0776_ ;
 wire \hash/_0777_ ;
 wire \hash/_0778_ ;
 wire \hash/_0779_ ;
 wire \hash/_0780_ ;
 wire \hash/_0781_ ;
 wire \hash/_0782_ ;
 wire \hash/_0783_ ;
 wire \hash/_0785_ ;
 wire \hash/_0786_ ;
 wire \hash/_0787_ ;
 wire \hash/_0788_ ;
 wire \hash/_0789_ ;
 wire \hash/_0790_ ;
 wire \hash/_0791_ ;
 wire \hash/_0792_ ;
 wire \hash/_0793_ ;
 wire \hash/_0794_ ;
 wire \hash/_0795_ ;
 wire \hash/_0796_ ;
 wire \hash/_0797_ ;
 wire \hash/_0798_ ;
 wire \hash/_0799_ ;
 wire \hash/_0800_ ;
 wire \hash/_0801_ ;
 wire \hash/_0802_ ;
 wire \hash/_0803_ ;
 wire \hash/_0804_ ;
 wire \hash/_0805_ ;
 wire \hash/_0806_ ;
 wire \hash/_0807_ ;
 wire \hash/_0808_ ;
 wire \hash/_0809_ ;
 wire \hash/_0810_ ;
 wire \hash/_0811_ ;
 wire \hash/_0812_ ;
 wire \hash/_0813_ ;
 wire \hash/_0814_ ;
 wire \hash/_0815_ ;
 wire \hash/_0816_ ;
 wire \hash/_0817_ ;
 wire \hash/_0818_ ;
 wire \hash/_0819_ ;
 wire \hash/_0820_ ;
 wire \hash/_0821_ ;
 wire \hash/_0822_ ;
 wire \hash/_0823_ ;
 wire \hash/_0824_ ;
 wire \hash/_0825_ ;
 wire \hash/_0826_ ;
 wire \hash/_0827_ ;
 wire \hash/_0829_ ;
 wire \hash/_0830_ ;
 wire \hash/_0831_ ;
 wire \hash/_0832_ ;
 wire \hash/_0833_ ;
 wire \hash/_0834_ ;
 wire \hash/_0835_ ;
 wire \hash/_0836_ ;
 wire \hash/_0837_ ;
 wire \hash/_0838_ ;
 wire \hash/_0839_ ;
 wire \hash/_0840_ ;
 wire \hash/_0841_ ;
 wire \hash/_0842_ ;
 wire \hash/_0843_ ;
 wire \hash/_0844_ ;
 wire \hash/_0845_ ;
 wire \hash/_0846_ ;
 wire \hash/_0847_ ;
 wire \hash/_0848_ ;
 wire \hash/_0849_ ;
 wire \hash/_0850_ ;
 wire \hash/_0851_ ;
 wire \hash/_0852_ ;
 wire \hash/_0853_ ;
 wire \hash/_0854_ ;
 wire \hash/_0855_ ;
 wire \hash/_0856_ ;
 wire \hash/_0857_ ;
 wire \hash/_0858_ ;
 wire \hash/_0859_ ;
 wire \hash/_0860_ ;
 wire \hash/_0861_ ;
 wire \hash/_0862_ ;
 wire \hash/_0863_ ;
 wire \hash/_0864_ ;
 wire \hash/_0865_ ;
 wire \hash/_0866_ ;
 wire \hash/_0867_ ;
 wire \hash/_0868_ ;
 wire \hash/_0869_ ;
 wire \hash/_0870_ ;
 wire \hash/_0871_ ;
 wire \hash/_0872_ ;
 wire \hash/_0873_ ;
 wire \hash/_0874_ ;
 wire \hash/_0875_ ;
 wire \hash/_0877_ ;
 wire \hash/_0878_ ;
 wire \hash/_0879_ ;
 wire \hash/_0880_ ;
 wire \hash/_0881_ ;
 wire \hash/_0882_ ;
 wire \hash/_0883_ ;
 wire \hash/_0884_ ;
 wire \hash/_0885_ ;
 wire \hash/_0886_ ;
 wire \hash/_0887_ ;
 wire \hash/_0888_ ;
 wire \hash/_0889_ ;
 wire \hash/_0890_ ;
 wire \hash/_0891_ ;
 wire \hash/_0892_ ;
 wire \hash/_0893_ ;
 wire \hash/_0894_ ;
 wire \hash/_0895_ ;
 wire \hash/_0896_ ;
 wire \hash/_0897_ ;
 wire \hash/_0898_ ;
 wire \hash/_0900_ ;
 wire \hash/_0901_ ;
 wire \hash/_0902_ ;
 wire \hash/_0903_ ;
 wire \hash/_0904_ ;
 wire \hash/_0905_ ;
 wire \hash/_0906_ ;
 wire \hash/_0907_ ;
 wire \hash/_0908_ ;
 wire \hash/_0909_ ;
 wire \hash/_0910_ ;
 wire \hash/_0911_ ;
 wire \hash/_0912_ ;
 wire \hash/_0913_ ;
 wire \hash/_0914_ ;
 wire \hash/_0915_ ;
 wire \hash/_0917_ ;
 wire \hash/_0918_ ;
 wire \hash/_0919_ ;
 wire \hash/_0920_ ;
 wire \hash/_0921_ ;
 wire \hash/_0922_ ;
 wire \hash/_0923_ ;
 wire \hash/_0924_ ;
 wire \hash/_0925_ ;
 wire \hash/_0926_ ;
 wire \hash/_0927_ ;
 wire \hash/_0928_ ;
 wire \hash/_0929_ ;
 wire \hash/_0930_ ;
 wire \hash/_0931_ ;
 wire \hash/_0932_ ;
 wire \hash/_0933_ ;
 wire \hash/_0934_ ;
 wire \hash/_0935_ ;
 wire \hash/_0936_ ;
 wire \hash/_0937_ ;
 wire \hash/_0938_ ;
 wire \hash/_0939_ ;
 wire \hash/_0940_ ;
 wire \hash/_0941_ ;
 wire \hash/_0942_ ;
 wire \hash/_0943_ ;
 wire \hash/_0944_ ;
 wire \hash/_0945_ ;
 wire \hash/_0946_ ;
 wire \hash/_0947_ ;
 wire \hash/_0948_ ;
 wire \hash/_0949_ ;
 wire \hash/_0950_ ;
 wire \hash/_0951_ ;
 wire \hash/_0952_ ;
 wire \hash/_0953_ ;
 wire \hash/_0954_ ;
 wire \hash/_0955_ ;
 wire \hash/_0956_ ;
 wire \hash/_0957_ ;
 wire \hash/_0958_ ;
 wire \hash/_0959_ ;
 wire \hash/_0960_ ;
 wire \hash/_0961_ ;
 wire \hash/_0962_ ;
 wire \hash/_0963_ ;
 wire \hash/_0964_ ;
 wire \hash/_0965_ ;
 wire \hash/_0966_ ;
 wire \hash/_0967_ ;
 wire \hash/_0968_ ;
 wire \hash/_0969_ ;
 wire \hash/_0970_ ;
 wire \hash/_0971_ ;
 wire \hash/_0972_ ;
 wire \hash/_0973_ ;
 wire \hash/_0974_ ;
 wire \hash/_0975_ ;
 wire \hash/_0976_ ;
 wire \hash/_0977_ ;
 wire \hash/_0978_ ;
 wire \hash/_0979_ ;
 wire \hash/_0980_ ;
 wire \hash/_0981_ ;
 wire \hash/_0982_ ;
 wire \hash/_0983_ ;
 wire \hash/_0984_ ;
 wire \hash/_0985_ ;
 wire \hash/_0986_ ;
 wire \hash/_0987_ ;
 wire \hash/_0988_ ;
 wire \hash/_0989_ ;
 wire \hash/_0990_ ;
 wire \hash/_0991_ ;
 wire \hash/_0992_ ;
 wire \hash/_0993_ ;
 wire \hash/_0994_ ;
 wire \hash/_0995_ ;
 wire \hash/_0996_ ;
 wire \hash/_0997_ ;
 wire \hash/_0998_ ;
 wire \hash/_0999_ ;
 wire \hash/_1000_ ;
 wire \hash/_1002_ ;
 wire \hash/_1003_ ;
 wire \hash/_1004_ ;
 wire \hash/_1005_ ;
 wire \hash/_1006_ ;
 wire \hash/_1007_ ;
 wire \hash/_1008_ ;
 wire \hash/_1009_ ;
 wire \hash/_1010_ ;
 wire \hash/_1011_ ;
 wire \hash/_1012_ ;
 wire \hash/_1013_ ;
 wire \hash/_1015_ ;
 wire \hash/_1016_ ;
 wire \hash/_1017_ ;
 wire \hash/_1018_ ;
 wire \hash/_1019_ ;
 wire \hash/_1020_ ;
 wire \hash/_1021_ ;
 wire \hash/_1022_ ;
 wire \hash/_1023_ ;
 wire \hash/_1024_ ;
 wire \hash/_1025_ ;
 wire \hash/_1026_ ;
 wire \hash/_1027_ ;
 wire \hash/_1028_ ;
 wire \hash/_1029_ ;
 wire \hash/_1030_ ;
 wire \hash/_1031_ ;
 wire \hash/_1032_ ;
 wire \hash/_1033_ ;
 wire \hash/_1034_ ;
 wire \hash/_1035_ ;
 wire \hash/_1036_ ;
 wire \hash/_1037_ ;
 wire \hash/_1038_ ;
 wire \hash/_1039_ ;
 wire \hash/_1040_ ;
 wire \hash/_1041_ ;
 wire \hash/_1042_ ;
 wire \hash/_1043_ ;
 wire \hash/_1044_ ;
 wire \hash/_1045_ ;
 wire \hash/_1046_ ;
 wire \hash/_1047_ ;
 wire \hash/_1048_ ;
 wire \hash/_1049_ ;
 wire \hash/_1050_ ;
 wire \hash/_1051_ ;
 wire \hash/_1052_ ;
 wire \hash/_1053_ ;
 wire \hash/_1054_ ;
 wire \hash/_1055_ ;
 wire \hash/_1056_ ;
 wire \hash/_1057_ ;
 wire \hash/_1058_ ;
 wire \hash/_1059_ ;
 wire \hash/_1060_ ;
 wire \hash/_1061_ ;
 wire \hash/_1062_ ;
 wire \hash/_1063_ ;
 wire \hash/_1064_ ;
 wire \hash/_1065_ ;
 wire \hash/_1066_ ;
 wire \hash/_1067_ ;
 wire \hash/_1068_ ;
 wire \hash/_1069_ ;
 wire \hash/_1071_ ;
 wire \hash/_1072_ ;
 wire \hash/_1073_ ;
 wire \hash/_1074_ ;
 wire \hash/_1075_ ;
 wire \hash/_1076_ ;
 wire \hash/_1077_ ;
 wire \hash/_1078_ ;
 wire \hash/_1079_ ;
 wire \hash/_1080_ ;
 wire \hash/_1081_ ;
 wire \hash/_1082_ ;
 wire \hash/_1083_ ;
 wire \hash/_1084_ ;
 wire \hash/_1085_ ;
 wire \hash/_1086_ ;
 wire \hash/_1087_ ;
 wire \hash/_1088_ ;
 wire \hash/_1089_ ;
 wire \hash/_1090_ ;
 wire \hash/_1091_ ;
 wire \hash/_1092_ ;
 wire \hash/_1093_ ;
 wire \hash/_1094_ ;
 wire \hash/_1095_ ;
 wire \hash/_1096_ ;
 wire \hash/_1097_ ;
 wire \hash/_1098_ ;
 wire \hash/_1099_ ;
 wire \hash/_1100_ ;
 wire \hash/_1101_ ;
 wire \hash/_1102_ ;
 wire \hash/_1103_ ;
 wire \hash/_1104_ ;
 wire \hash/_1105_ ;
 wire \hash/_1106_ ;
 wire \hash/_1107_ ;
 wire \hash/_1108_ ;
 wire \hash/_1109_ ;
 wire \hash/_1110_ ;
 wire \hash/_1111_ ;
 wire \hash/_1112_ ;
 wire \hash/_1113_ ;
 wire \hash/_1114_ ;
 wire \hash/_1115_ ;
 wire \hash/_1116_ ;
 wire \hash/_1117_ ;
 wire \hash/_1118_ ;
 wire \hash/_1119_ ;
 wire \hash/_1120_ ;
 wire \hash/_1121_ ;
 wire \hash/_1122_ ;
 wire \hash/_1123_ ;
 wire \hash/_1124_ ;
 wire \hash/_1125_ ;
 wire \hash/_1126_ ;
 wire \hash/_1127_ ;
 wire \hash/_1128_ ;
 wire \hash/_1129_ ;
 wire \hash/_1130_ ;
 wire \hash/_1131_ ;
 wire \hash/_1132_ ;
 wire \hash/_1133_ ;
 wire \hash/_1134_ ;
 wire \hash/_1135_ ;
 wire \hash/_1136_ ;
 wire \hash/_1137_ ;
 wire \hash/_1138_ ;
 wire \hash/_1139_ ;
 wire \hash/_1140_ ;
 wire \hash/_1141_ ;
 wire \hash/_1142_ ;
 wire \hash/_1143_ ;
 wire \hash/_1144_ ;
 wire \hash/_1145_ ;
 wire \hash/_1146_ ;
 wire \hash/_1147_ ;
 wire \hash/_1148_ ;
 wire \hash/_1149_ ;
 wire \hash/_1150_ ;
 wire \hash/_1151_ ;
 wire \hash/_1152_ ;
 wire \hash/_1153_ ;
 wire \hash/_1154_ ;
 wire \hash/_1155_ ;
 wire \hash/_1156_ ;
 wire \hash/_1157_ ;
 wire \hash/_1158_ ;
 wire \hash/_1159_ ;
 wire \hash/_1160_ ;
 wire \hash/_1161_ ;
 wire \hash/_1162_ ;
 wire \hash/_1163_ ;
 wire \hash/_1164_ ;
 wire \hash/_1165_ ;
 wire \hash/_1166_ ;
 wire \hash/_1167_ ;
 wire \hash/_1168_ ;
 wire \hash/_1169_ ;
 wire \hash/_1170_ ;
 wire \hash/_1171_ ;
 wire \hash/_1172_ ;
 wire \hash/_1173_ ;
 wire \hash/_1174_ ;
 wire \hash/_1175_ ;
 wire \hash/_1176_ ;
 wire \hash/_1177_ ;
 wire \hash/_1178_ ;
 wire \hash/_1179_ ;
 wire \hash/_1180_ ;
 wire \hash/_1181_ ;
 wire \hash/_1182_ ;
 wire \hash/_1183_ ;
 wire \hash/_1184_ ;
 wire \hash/_1185_ ;
 wire \hash/_1186_ ;
 wire \hash/_1187_ ;
 wire \hash/_1188_ ;
 wire \hash/_1189_ ;
 wire \hash/_1190_ ;
 wire \hash/_1191_ ;
 wire \hash/_1192_ ;
 wire \hash/_1193_ ;
 wire \hash/_1194_ ;
 wire \hash/_1195_ ;
 wire \hash/_1196_ ;
 wire \hash/_1197_ ;
 wire \hash/_1198_ ;
 wire \hash/_1199_ ;
 wire \hash/_1200_ ;
 wire \hash/_1201_ ;
 wire \hash/_1202_ ;
 wire \hash/_1203_ ;
 wire \hash/_1204_ ;
 wire \hash/_1205_ ;
 wire \hash/_1206_ ;
 wire \hash/_1207_ ;
 wire \hash/_1208_ ;
 wire \hash/_1209_ ;
 wire \hash/_1210_ ;
 wire \hash/_1211_ ;
 wire \hash/_1212_ ;
 wire \hash/_1213_ ;
 wire \hash/_1214_ ;
 wire \hash/_1215_ ;
 wire \hash/_1216_ ;
 wire \hash/_1217_ ;
 wire \hash/_1218_ ;
 wire \hash/_1219_ ;
 wire \hash/_1220_ ;
 wire \hash/_1221_ ;
 wire \hash/_1222_ ;
 wire \hash/_1223_ ;
 wire \hash/_1224_ ;
 wire \hash/_1225_ ;
 wire \hash/_1226_ ;
 wire \hash/_1227_ ;
 wire \hash/_1228_ ;
 wire \hash/_1229_ ;
 wire \hash/_1230_ ;
 wire \hash/_1231_ ;
 wire \hash/_1232_ ;
 wire \hash/_1233_ ;
 wire \hash/_1234_ ;
 wire \hash/_1235_ ;
 wire \hash/_1236_ ;
 wire \hash/_1237_ ;
 wire \hash/_1238_ ;
 wire \hash/_1239_ ;
 wire \hash/_1240_ ;
 wire \hash/_1241_ ;
 wire \hash/_1242_ ;
 wire \hash/_1243_ ;
 wire \hash/_1244_ ;
 wire \hash/_1245_ ;
 wire \hash/_1246_ ;
 wire \hash/_1247_ ;
 wire \hash/_1248_ ;
 wire \hash/_1249_ ;
 wire \hash/_1250_ ;
 wire \hash/_1251_ ;
 wire \hash/_1252_ ;
 wire \hash/_1253_ ;
 wire \hash/_1254_ ;
 wire \hash/_1255_ ;
 wire \hash/_1256_ ;
 wire \hash/_1257_ ;
 wire \hash/_1258_ ;
 wire \hash/_1259_ ;
 wire \hash/_1260_ ;
 wire \hash/_1261_ ;
 wire \hash/_1262_ ;
 wire \hash/_1263_ ;
 wire \hash/_1264_ ;
 wire \hash/_1265_ ;
 wire \hash/_1266_ ;
 wire \hash/_1267_ ;
 wire \hash/_1268_ ;
 wire \hash/_1269_ ;
 wire \hash/_1270_ ;
 wire \hash/_1271_ ;
 wire \hash/_1272_ ;
 wire \hash/_1273_ ;
 wire \hash/_1274_ ;
 wire \hash/_1275_ ;
 wire \hash/_1276_ ;
 wire \hash/_1277_ ;
 wire \hash/_1278_ ;
 wire \hash/_1279_ ;
 wire \hash/_1280_ ;
 wire \hash/_1281_ ;
 wire \hash/_1282_ ;
 wire \hash/_1283_ ;
 wire \hash/_1284_ ;
 wire \hash/_1285_ ;
 wire \hash/_1286_ ;
 wire \hash/_1287_ ;
 wire \hash/_1288_ ;
 wire \hash/_1289_ ;
 wire \hash/_1290_ ;
 wire \hash/_1291_ ;
 wire \hash/_1292_ ;
 wire \hash/_1293_ ;
 wire \hash/_1294_ ;
 wire \hash/_1295_ ;
 wire \hash/_1296_ ;
 wire \hash/_1297_ ;
 wire \hash/_1298_ ;
 wire \hash/_1299_ ;
 wire \hash/_1300_ ;
 wire \hash/_1301_ ;
 wire \hash/_1302_ ;
 wire \hash/_1303_ ;
 wire \hash/_1304_ ;
 wire \hash/_1305_ ;
 wire \hash/_1306_ ;
 wire \hash/_1307_ ;
 wire \hash/_1308_ ;
 wire \hash/_1309_ ;
 wire \hash/_1310_ ;
 wire \hash/_1311_ ;
 wire \hash/_1312_ ;
 wire \hash/_1313_ ;
 wire \hash/_1314_ ;
 wire \hash/_1315_ ;
 wire \hash/_1316_ ;
 wire \hash/_1317_ ;
 wire \hash/_1318_ ;
 wire \hash/_1319_ ;
 wire \hash/_1320_ ;
 wire \hash/_1321_ ;
 wire \hash/_1322_ ;
 wire \hash/_1323_ ;
 wire \hash/_1324_ ;
 wire \hash/_1325_ ;
 wire \hash/_1326_ ;
 wire \hash/_1327_ ;
 wire \hash/_1328_ ;
 wire \hash/_1329_ ;
 wire \hash/_1330_ ;
 wire \hash/_1331_ ;
 wire \hash/_1332_ ;
 wire \hash/_1333_ ;
 wire \hash/_1334_ ;
 wire \hash/_1335_ ;
 wire \hash/_1336_ ;
 wire \hash/_1337_ ;
 wire \hash/_1338_ ;
 wire \hash/_1339_ ;
 wire \hash/_1340_ ;
 wire \hash/_1341_ ;
 wire \hash/_1342_ ;
 wire \hash/_1343_ ;
 wire \hash/_1344_ ;
 wire \hash/_1345_ ;
 wire \hash/_1346_ ;
 wire \hash/_1347_ ;
 wire \hash/_1348_ ;
 wire \hash/_1349_ ;
 wire \hash/_1350_ ;
 wire \hash/_1351_ ;
 wire \hash/_1352_ ;
 wire \hash/_1353_ ;
 wire \hash/_1354_ ;
 wire \hash/_1355_ ;
 wire \hash/_1356_ ;
 wire \hash/_1357_ ;
 wire \hash/_1358_ ;
 wire \hash/_1359_ ;
 wire \hash/_1360_ ;
 wire \hash/_1361_ ;
 wire \hash/_1362_ ;
 wire \hash/_1363_ ;
 wire \hash/_1364_ ;
 wire \hash/_1365_ ;
 wire \hash/_1366_ ;
 wire \hash/_1367_ ;
 wire \hash/_1368_ ;
 wire \hash/_1369_ ;
 wire \hash/_1370_ ;
 wire \hash/_1371_ ;
 wire \hash/_1372_ ;
 wire \hash/_1373_ ;
 wire \hash/_1374_ ;
 wire \hash/_1375_ ;
 wire \hash/_1376_ ;
 wire \hash/_1377_ ;
 wire \hash/_1378_ ;
 wire \hash/_1379_ ;
 wire \hash/_1380_ ;
 wire \hash/_1381_ ;
 wire \hash/_1382_ ;
 wire \hash/_1383_ ;
 wire \hash/_1384_ ;
 wire \hash/_1385_ ;
 wire \hash/_1386_ ;
 wire \hash/_1387_ ;
 wire \hash/_1388_ ;
 wire \hash/_1389_ ;
 wire \hash/_1390_ ;
 wire \hash/_1391_ ;
 wire \hash/_1392_ ;
 wire \hash/_1393_ ;
 wire \hash/_1394_ ;
 wire \hash/_1395_ ;
 wire \hash/_1396_ ;
 wire \hash/_1397_ ;
 wire \hash/_1398_ ;
 wire \hash/_1399_ ;
 wire \hash/_1400_ ;
 wire \hash/_1401_ ;
 wire \hash/_1402_ ;
 wire \hash/_1403_ ;
 wire \hash/_1404_ ;
 wire \hash/_1405_ ;
 wire \hash/_1406_ ;
 wire \hash/_1407_ ;
 wire \hash/_1408_ ;
 wire \hash/_1409_ ;
 wire \hash/_1410_ ;
 wire \hash/_1411_ ;
 wire \hash/_1412_ ;
 wire \hash/_1413_ ;
 wire \hash/_1414_ ;
 wire \hash/_1415_ ;
 wire \hash/_1416_ ;
 wire \hash/_1417_ ;
 wire \hash/_1418_ ;
 wire \hash/_1445_ ;
 wire \hash/_1446_ ;
 wire \hash/_1447_ ;
 wire \hash/_1448_ ;
 wire \hash/_1449_ ;
 wire \hash/_1450_ ;
 wire \hash/_1451_ ;
 wire \hash/_1452_ ;
 wire \hash/_1453_ ;
 wire \hash/_1454_ ;
 wire \hash/_1455_ ;
 wire \hash/_1456_ ;
 wire \hash/_1457_ ;
 wire \hash/_1458_ ;
 wire \hash/_1459_ ;
 wire \hash/_1460_ ;
 wire \hash/_1461_ ;
 wire \hash/_1462_ ;
 wire \hash/_1463_ ;
 wire \hash/_1464_ ;
 wire \hash/_1465_ ;
 wire \hash/_1466_ ;
 wire \hash/_1467_ ;
 wire \hash/_1468_ ;
 wire \hash/_1469_ ;
 wire \hash/_1470_ ;
 wire \hash/_1471_ ;
 wire \hash/_1472_ ;
 wire \hash/_1473_ ;
 wire \hash/_1474_ ;
 wire \hash/_1475_ ;
 wire \hash/_1476_ ;
 wire \hash/_1477_ ;
 wire \hash/_1478_ ;
 wire \hash/_1479_ ;
 wire \hash/_1480_ ;
 wire \hash/_1481_ ;
 wire \hash/_1482_ ;
 wire \hash/_1483_ ;
 wire \hash/_1484_ ;
 wire \hash/_1485_ ;
 wire \hash/_1486_ ;
 wire \hash/_1487_ ;
 wire \hash/_1488_ ;
 wire \hash/_1489_ ;
 wire \hash/_1490_ ;
 wire \hash/_1491_ ;
 wire \hash/_1492_ ;
 wire \hash/_1493_ ;
 wire \hash/_1494_ ;
 wire \hash/_1495_ ;
 wire \hash/_1496_ ;
 wire \hash/_1497_ ;
 wire \hash/_1498_ ;
 wire \hash/_1499_ ;
 wire \hash/_1500_ ;
 wire \hash/_1501_ ;
 wire \hash/_1502_ ;
 wire \hash/_1503_ ;
 wire \hash/_1504_ ;
 wire \hash/_1505_ ;
 wire \hash/_1506_ ;
 wire \hash/_1507_ ;
 wire \hash/_1508_ ;
 wire \hash/_1509_ ;
 wire \hash/_1510_ ;
 wire \hash/_1511_ ;
 wire \hash/_1512_ ;
 wire \hash/_1513_ ;
 wire \hash/_1514_ ;
 wire \hash/_1515_ ;
 wire \hash/_1516_ ;
 wire \hash/_1517_ ;
 wire \hash/_1518_ ;
 wire \hash/_1519_ ;
 wire \hash/_1520_ ;
 wire \hash/_1521_ ;
 wire \hash/_1522_ ;
 wire \hash/_1523_ ;
 wire \hash/_1524_ ;
 wire \hash/_1525_ ;
 wire \hash/_1526_ ;
 wire \hash/_1527_ ;
 wire \hash/_1528_ ;
 wire \hash/_1529_ ;
 wire \hash/_1530_ ;
 wire \hash/_1531_ ;
 wire \hash/_1532_ ;
 wire \hash/_1533_ ;
 wire \hash/_1534_ ;
 wire \hash/_1535_ ;
 wire \hash/_1536_ ;
 wire \hash/_1537_ ;
 wire \hash/_1538_ ;
 wire \hash/_1539_ ;
 wire \hash/_1540_ ;
 wire \hash/_1541_ ;
 wire \hash/_1542_ ;
 wire \hash/_1543_ ;
 wire \hash/_1544_ ;
 wire \hash/_1545_ ;
 wire \hash/_1546_ ;
 wire \hash/_1547_ ;
 wire \hash/_1548_ ;
 wire \hash/_1549_ ;
 wire \hash/_1550_ ;
 wire \hash/_1551_ ;
 wire \hash/_1552_ ;
 wire \hash/_1553_ ;
 wire \hash/_1554_ ;
 wire \hash/_1555_ ;
 wire \hash/_1556_ ;
 wire \hash/_1557_ ;
 wire \hash/_1558_ ;
 wire \hash/_1559_ ;
 wire \hash/_1560_ ;
 wire \hash/_1561_ ;
 wire \hash/_1562_ ;
 wire \hash/_1563_ ;
 wire \hash/_1564_ ;
 wire \hash/_1565_ ;
 wire \hash/_1566_ ;
 wire \hash/_1567_ ;
 wire \hash/_1568_ ;
 wire \hash/_1569_ ;
 wire \hash/_1570_ ;
 wire \hash/_1571_ ;
 wire \hash/_1572_ ;
 wire \hash/_1573_ ;
 wire \hash/_1574_ ;
 wire \hash/_1575_ ;
 wire \hash/_1576_ ;
 wire \hash/_1577_ ;
 wire \hash/_1578_ ;
 wire \hash/_1579_ ;
 wire \hash/_1580_ ;
 wire \hash/_1581_ ;
 wire \hash/_1582_ ;
 wire \hash/_1583_ ;
 wire \hash/_1584_ ;
 wire \hash/_1585_ ;
 wire \hash/_1586_ ;
 wire \hash/_1587_ ;
 wire \hash/_1588_ ;
 wire \hash/_1589_ ;
 wire \hash/_1590_ ;
 wire \hash/_1591_ ;
 wire \hash/_1592_ ;
 wire \hash/_1593_ ;
 wire \hash/_1594_ ;
 wire \hash/_1595_ ;
 wire \hash/_1596_ ;
 wire \hash/_1597_ ;
 wire \hash/_1598_ ;
 wire \hash/_1599_ ;
 wire \hash/_1600_ ;
 wire \hash/_1601_ ;
 wire \hash/_1602_ ;
 wire \hash/_1603_ ;
 wire \hash/_1604_ ;
 wire \hash/_1605_ ;
 wire \hash/_1606_ ;
 wire \hash/_1607_ ;
 wire \hash/_1608_ ;
 wire \hash/_1609_ ;
 wire \hash/_1610_ ;
 wire \hash/_1611_ ;
 wire \hash/_1612_ ;
 wire \hash/_1613_ ;
 wire \hash/_1614_ ;
 wire \hash/_1615_ ;
 wire \hash/_1616_ ;
 wire \hash/_1617_ ;
 wire \hash/_1618_ ;
 wire \hash/_1619_ ;
 wire \hash/_1620_ ;
 wire \hash/_1621_ ;
 wire \hash/_1622_ ;
 wire \hash/_1623_ ;
 wire \hash/_1624_ ;
 wire \hash/_1625_ ;
 wire \hash/_1626_ ;
 wire \hash/_1627_ ;
 wire \hash/_1628_ ;
 wire \hash/_1629_ ;
 wire \hash/_1630_ ;
 wire \hash/_1631_ ;
 wire \hash/_1632_ ;
 wire \hash/_1633_ ;
 wire \hash/_1634_ ;
 wire \hash/_1635_ ;
 wire \hash/_1636_ ;
 wire \hash/_1637_ ;
 wire \hash/_1638_ ;
 wire \hash/_1639_ ;
 wire \hash/_1640_ ;
 wire \hash/_1641_ ;
 wire \hash/_1642_ ;
 wire \hash/_1643_ ;
 wire \hash/_1644_ ;
 wire \hash/_1645_ ;
 wire \hash/_1646_ ;
 wire \hash/_1647_ ;
 wire \hash/_1648_ ;
 wire \hash/_1649_ ;
 wire \hash/_1650_ ;
 wire \hash/_1651_ ;
 wire \hash/_1652_ ;
 wire \hash/_1653_ ;
 wire \hash/_1654_ ;
 wire \hash/_1655_ ;
 wire \hash/_1656_ ;
 wire \hash/_1657_ ;
 wire \hash/_1658_ ;
 wire \hash/_1659_ ;
 wire \hash/_1660_ ;
 wire \hash/_1661_ ;
 wire \hash/_1662_ ;
 wire \hash/_1663_ ;
 wire \hash/_1664_ ;
 wire \hash/_1665_ ;
 wire \hash/_1666_ ;
 wire \hash/_1667_ ;
 wire \hash/_1668_ ;
 wire \hash/_1669_ ;
 wire \hash/_1670_ ;
 wire \hash/_1671_ ;
 wire \hash/_1672_ ;
 wire \hash/_1673_ ;
 wire \hash/_1674_ ;
 wire \hash/_1675_ ;
 wire \hash/_1676_ ;
 wire \hash/_1677_ ;
 wire \hash/_1678_ ;
 wire \hash/_1679_ ;
 wire \hash/_1680_ ;
 wire \hash/_1681_ ;
 wire \hash/_1682_ ;
 wire \hash/_1683_ ;
 wire \hash/_1684_ ;
 wire \hash/_1685_ ;
 wire \hash/_1686_ ;
 wire \hash/_1687_ ;
 wire \hash/_1688_ ;
 wire \hash/_1689_ ;
 wire \hash/_1690_ ;
 wire \hash/_1691_ ;
 wire \hash/_1692_ ;
 wire \hash/_1693_ ;
 wire \hash/_1694_ ;
 wire \hash/_1695_ ;
 wire \hash/_1696_ ;
 wire \hash/_1697_ ;
 wire \hash/_1698_ ;
 wire \hash/_1699_ ;
 wire \hash/_1700_ ;
 wire \hash/_1701_ ;
 wire \hash/_1702_ ;
 wire \hash/_1703_ ;
 wire \hash/_1704_ ;
 wire \hash/_1705_ ;
 wire \hash/_1706_ ;
 wire \hash/_1707_ ;
 wire \hash/_1708_ ;
 wire \hash/_1709_ ;
 wire \hash/_1710_ ;
 wire \hash/_1711_ ;
 wire \hash/_1712_ ;
 wire \hash/_1713_ ;
 wire \hash/_1714_ ;
 wire \hash/_1715_ ;
 wire \hash/_1716_ ;
 wire \hash/_1717_ ;
 wire \hash/_1718_ ;
 wire \hash/_1719_ ;
 wire \hash/_1720_ ;
 wire \hash/_1721_ ;
 wire \hash/_1722_ ;
 wire \hash/_1723_ ;
 wire \hash/_1724_ ;
 wire \hash/_1725_ ;
 wire \hash/_1726_ ;
 wire \hash/_1727_ ;
 wire \hash/_1728_ ;
 wire \hash/_1729_ ;
 wire \hash/_1730_ ;
 wire \hash/_1731_ ;
 wire \hash/_1732_ ;
 wire \hash/_1733_ ;
 wire \hash/_1734_ ;
 wire \hash/_1735_ ;
 wire \hash/_1736_ ;
 wire \hash/_1737_ ;
 wire \hash/_1738_ ;
 wire \hash/_1739_ ;
 wire \hash/_1740_ ;
 wire \hash/_1741_ ;
 wire \hash/_1742_ ;
 wire \hash/_1743_ ;
 wire \hash/_1744_ ;
 wire \hash/_1745_ ;
 wire \hash/_1746_ ;
 wire \hash/_1747_ ;
 wire \hash/_1748_ ;
 wire \hash/_1749_ ;
 wire \hash/_1750_ ;
 wire \hash/_1751_ ;
 wire \hash/_1752_ ;
 wire \hash/_1753_ ;
 wire \hash/_1754_ ;
 wire \hash/_1755_ ;
 wire \hash/_1756_ ;
 wire \hash/_1757_ ;
 wire \hash/_1758_ ;
 wire \hash/_1759_ ;
 wire \hash/_1760_ ;
 wire \hash/_1761_ ;
 wire \hash/_1762_ ;
 wire \hash/_1763_ ;
 wire \hash/_1764_ ;
 wire \hash/_1765_ ;
 wire \hash/_1766_ ;
 wire \hash/_1767_ ;
 wire \hash/_1768_ ;
 wire \hash/_1769_ ;
 wire \hash/_1770_ ;
 wire \hash/_1771_ ;
 wire \hash/_1772_ ;
 wire \hash/_1773_ ;
 wire \hash/_1774_ ;
 wire \hash/_1775_ ;
 wire \hash/_1776_ ;
 wire \hash/_1777_ ;
 wire \hash/_1778_ ;
 wire \hash/_1779_ ;
 wire \hash/_1780_ ;
 wire \hash/_1781_ ;
 wire \hash/_1782_ ;
 wire \hash/_1783_ ;
 wire \hash/_1784_ ;
 wire \hash/_1785_ ;
 wire \hash/_1786_ ;
 wire \hash/_1787_ ;
 wire \hash/_1788_ ;
 wire \hash/_1789_ ;
 wire \hash/_1790_ ;
 wire \hash/_1791_ ;
 wire \hash/_1792_ ;
 wire \hash/_1793_ ;
 wire \hash/_1794_ ;
 wire \hash/_1795_ ;
 wire \hash/_1796_ ;
 wire \hash/_1797_ ;
 wire \hash/_1798_ ;
 wire \hash/_1799_ ;
 wire \hash/_1800_ ;
 wire \hash/_1801_ ;
 wire \hash/_1802_ ;
 wire \hash/_1803_ ;
 wire \hash/_1804_ ;
 wire \hash/_1805_ ;
 wire \hash/_1806_ ;
 wire \hash/_1807_ ;
 wire \hash/_1808_ ;
 wire \hash/_1809_ ;
 wire \hash/_1810_ ;
 wire \hash/_1811_ ;
 wire \hash/_1812_ ;
 wire \hash/_1813_ ;
 wire \hash/_1814_ ;
 wire \hash/_1815_ ;
 wire \hash/_1816_ ;
 wire \hash/_1817_ ;
 wire \hash/_1818_ ;
 wire \hash/_1819_ ;
 wire \hash/_1820_ ;
 wire \hash/_1821_ ;
 wire \hash/_1822_ ;
 wire \hash/_1823_ ;
 wire \hash/_1824_ ;
 wire \hash/_1825_ ;
 wire \hash/_1826_ ;
 wire \hash/_1827_ ;
 wire \hash/_1828_ ;
 wire \hash/_1829_ ;
 wire \hash/_1830_ ;
 wire \hash/_1831_ ;
 wire \hash/_1832_ ;
 wire \hash/_1833_ ;
 wire \hash/_1834_ ;
 wire \hash/_1835_ ;
 wire \hash/_1836_ ;
 wire \hash/_1837_ ;
 wire \hash/_1838_ ;
 wire \hash/_1839_ ;
 wire \hash/_1840_ ;
 wire \hash/_1841_ ;
 wire \hash/_1842_ ;
 wire \hash/_1843_ ;
 wire \hash/_1844_ ;
 wire \hash/_1845_ ;
 wire \hash/_1846_ ;
 wire \hash/_1847_ ;
 wire \hash/_1848_ ;
 wire \hash/_1849_ ;
 wire \hash/_1850_ ;
 wire \hash/_1851_ ;
 wire \hash/_1852_ ;
 wire \hash/_1853_ ;
 wire \hash/_1854_ ;
 wire \hash/_1855_ ;
 wire \hash/_1856_ ;
 wire \hash/_1857_ ;
 wire \hash/_1858_ ;
 wire \hash/_1859_ ;
 wire \hash/_1860_ ;
 wire \hash/_1861_ ;
 wire \hash/_1862_ ;
 wire \hash/_1863_ ;
 wire \hash/_1864_ ;
 wire \hash/_1865_ ;
 wire \hash/_1866_ ;
 wire \hash/_1867_ ;
 wire \hash/_1868_ ;
 wire \hash/_1869_ ;
 wire \hash/_1870_ ;
 wire \hash/_1871_ ;
 wire \hash/_1872_ ;
 wire \hash/_1873_ ;
 wire \hash/_1874_ ;
 wire \hash/_1875_ ;
 wire \hash/_1876_ ;
 wire \hash/_1877_ ;
 wire \hash/_1878_ ;
 wire \hash/_1879_ ;
 wire \hash/_1880_ ;
 wire \hash/_1881_ ;
 wire \hash/_1882_ ;
 wire \hash/_1883_ ;
 wire \hash/_1884_ ;
 wire \hash/_1885_ ;
 wire \hash/_1886_ ;
 wire \hash/_1887_ ;
 wire \hash/_1888_ ;
 wire \hash/_1889_ ;
 wire \hash/_1890_ ;
 wire \hash/_1891_ ;
 wire \hash/_1892_ ;
 wire \hash/_1893_ ;
 wire \hash/_1894_ ;
 wire \hash/_1895_ ;
 wire \hash/_1896_ ;
 wire \hash/_1897_ ;
 wire \hash/_1898_ ;
 wire \hash/_1899_ ;
 wire \hash/_1900_ ;
 wire \hash/_1901_ ;
 wire \hash/_1902_ ;
 wire \hash/_1903_ ;
 wire \hash/_1904_ ;
 wire \hash/_1905_ ;
 wire \hash/_1906_ ;
 wire \hash/_1907_ ;
 wire \hash/_1908_ ;
 wire \hash/_1909_ ;
 wire \hash/_1910_ ;
 wire \hash/_1911_ ;
 wire \hash/_1912_ ;
 wire \hash/_1913_ ;
 wire \hash/_1914_ ;
 wire \hash/_1915_ ;
 wire \hash/_1916_ ;
 wire \hash/_1917_ ;
 wire \hash/_1918_ ;
 wire \hash/_1919_ ;
 wire \hash/_1920_ ;
 wire \hash/_1921_ ;
 wire \hash/_1922_ ;
 wire \hash/_1923_ ;
 wire \hash/_1924_ ;
 wire \hash/_1925_ ;
 wire \hash/_1926_ ;
 wire \hash/_1927_ ;
 wire \hash/_1928_ ;
 wire \hash/_1929_ ;
 wire \hash/_1930_ ;
 wire \hash/_1931_ ;
 wire \hash/_1932_ ;
 wire \hash/_1933_ ;
 wire \hash/_1934_ ;
 wire \hash/_1935_ ;
 wire \hash/_1936_ ;
 wire \hash/_1937_ ;
 wire \hash/_1938_ ;
 wire \hash/_1939_ ;
 wire \hash/_1940_ ;
 wire \hash/_1941_ ;
 wire \hash/_1942_ ;
 wire \hash/_1943_ ;
 wire \hash/_1944_ ;
 wire \hash/_1945_ ;
 wire \hash/_1946_ ;
 wire \hash/_1947_ ;
 wire \hash/_1948_ ;
 wire \hash/_1949_ ;
 wire \hash/_1950_ ;
 wire \hash/_1951_ ;
 wire \hash/_1952_ ;
 wire \hash/_1953_ ;
 wire \hash/_1954_ ;
 wire \hash/_1955_ ;
 wire \hash/_1956_ ;
 wire \hash/a[0] ;
 wire \hash/a[10] ;
 wire \hash/a[11] ;
 wire \hash/a[12] ;
 wire \hash/a[13] ;
 wire \hash/a[14] ;
 wire \hash/a[15] ;
 wire \hash/a[16] ;
 wire \hash/a[17] ;
 wire \hash/a[18] ;
 wire \hash/a[19] ;
 wire \hash/a[1] ;
 wire \hash/a[20] ;
 wire \hash/a[21] ;
 wire \hash/a[22] ;
 wire \hash/a[23] ;
 wire \hash/a[24] ;
 wire \hash/a[25] ;
 wire \hash/a[26] ;
 wire \hash/a[27] ;
 wire \hash/a[28] ;
 wire \hash/a[29] ;
 wire \hash/a[2] ;
 wire \hash/a[30] ;
 wire \hash/a[31] ;
 wire \hash/a[3] ;
 wire \hash/a[4] ;
 wire \hash/a[5] ;
 wire \hash/a[6] ;
 wire \hash/a[7] ;
 wire \hash/a[8] ;
 wire \hash/a[9] ;
 wire \hash/a_cap[0] ;
 wire \hash/a_cap[10] ;
 wire \hash/a_cap[11] ;
 wire \hash/a_cap[12] ;
 wire \hash/a_cap[13] ;
 wire \hash/a_cap[14] ;
 wire \hash/a_cap[15] ;
 wire \hash/a_cap[16] ;
 wire \hash/a_cap[17] ;
 wire \hash/a_cap[18] ;
 wire \hash/a_cap[19] ;
 wire \hash/a_cap[1] ;
 wire \hash/a_cap[20] ;
 wire \hash/a_cap[21] ;
 wire \hash/a_cap[22] ;
 wire \hash/a_cap[23] ;
 wire \hash/a_cap[24] ;
 wire \hash/a_cap[25] ;
 wire \hash/a_cap[26] ;
 wire \hash/a_cap[27] ;
 wire \hash/a_cap[28] ;
 wire \hash/a_cap[29] ;
 wire \hash/a_cap[2] ;
 wire \hash/a_cap[30] ;
 wire \hash/a_cap[31] ;
 wire \hash/a_cap[3] ;
 wire \hash/a_cap[4] ;
 wire \hash/a_cap[5] ;
 wire \hash/a_cap[6] ;
 wire \hash/a_cap[7] ;
 wire \hash/a_cap[8] ;
 wire \hash/a_cap[9] ;
 wire \hash/a_new[0] ;
 wire \hash/a_new[10] ;
 wire \hash/a_new[11] ;
 wire \hash/a_new[12] ;
 wire \hash/a_new[13] ;
 wire \hash/a_new[14] ;
 wire \hash/a_new[15] ;
 wire \hash/a_new[16] ;
 wire \hash/a_new[17] ;
 wire \hash/a_new[18] ;
 wire \hash/a_new[19] ;
 wire \hash/a_new[1] ;
 wire \hash/a_new[20] ;
 wire \hash/a_new[21] ;
 wire \hash/a_new[22] ;
 wire \hash/a_new[23] ;
 wire \hash/a_new[24] ;
 wire \hash/a_new[25] ;
 wire \hash/a_new[26] ;
 wire \hash/a_new[27] ;
 wire \hash/a_new[28] ;
 wire \hash/a_new[29] ;
 wire \hash/a_new[2] ;
 wire \hash/a_new[30] ;
 wire \hash/a_new[31] ;
 wire \hash/a_new[3] ;
 wire \hash/a_new[4] ;
 wire \hash/a_new[5] ;
 wire \hash/a_new[6] ;
 wire \hash/a_new[7] ;
 wire \hash/a_new[8] ;
 wire \hash/a_new[9] ;
 wire \hash/b[0] ;
 wire \hash/b[10] ;
 wire \hash/b[11] ;
 wire \hash/b[12] ;
 wire \hash/b[13] ;
 wire \hash/b[14] ;
 wire \hash/b[15] ;
 wire \hash/b[16] ;
 wire \hash/b[17] ;
 wire \hash/b[18] ;
 wire \hash/b[19] ;
 wire \hash/b[1] ;
 wire \hash/b[20] ;
 wire \hash/b[21] ;
 wire \hash/b[22] ;
 wire \hash/b[23] ;
 wire \hash/b[24] ;
 wire \hash/b[25] ;
 wire \hash/b[26] ;
 wire \hash/b[27] ;
 wire \hash/b[28] ;
 wire \hash/b[29] ;
 wire \hash/b[2] ;
 wire \hash/b[30] ;
 wire \hash/b[31] ;
 wire \hash/b[3] ;
 wire \hash/b[4] ;
 wire \hash/b[5] ;
 wire \hash/b[6] ;
 wire \hash/b[7] ;
 wire \hash/b[8] ;
 wire \hash/b[9] ;
 wire \hash/b_cap[0] ;
 wire \hash/b_cap[10] ;
 wire \hash/b_cap[11] ;
 wire \hash/b_cap[12] ;
 wire \hash/b_cap[13] ;
 wire \hash/b_cap[14] ;
 wire \hash/b_cap[15] ;
 wire \hash/b_cap[16] ;
 wire \hash/b_cap[17] ;
 wire \hash/b_cap[18] ;
 wire \hash/b_cap[19] ;
 wire \hash/b_cap[1] ;
 wire \hash/b_cap[20] ;
 wire \hash/b_cap[21] ;
 wire \hash/b_cap[22] ;
 wire \hash/b_cap[23] ;
 wire \hash/b_cap[24] ;
 wire \hash/b_cap[25] ;
 wire \hash/b_cap[26] ;
 wire \hash/b_cap[27] ;
 wire \hash/b_cap[28] ;
 wire \hash/b_cap[29] ;
 wire \hash/b_cap[2] ;
 wire \hash/b_cap[30] ;
 wire \hash/b_cap[31] ;
 wire \hash/b_cap[3] ;
 wire \hash/b_cap[4] ;
 wire \hash/b_cap[5] ;
 wire \hash/b_cap[6] ;
 wire \hash/b_cap[7] ;
 wire \hash/b_cap[8] ;
 wire \hash/b_cap[9] ;
 wire \hash/b_new[0] ;
 wire \hash/b_new[10] ;
 wire \hash/b_new[11] ;
 wire \hash/b_new[12] ;
 wire \hash/b_new[13] ;
 wire \hash/b_new[14] ;
 wire \hash/b_new[15] ;
 wire \hash/b_new[16] ;
 wire \hash/b_new[17] ;
 wire \hash/b_new[18] ;
 wire \hash/b_new[19] ;
 wire \hash/b_new[1] ;
 wire \hash/b_new[20] ;
 wire \hash/b_new[21] ;
 wire \hash/b_new[22] ;
 wire \hash/b_new[23] ;
 wire \hash/b_new[24] ;
 wire \hash/b_new[25] ;
 wire \hash/b_new[26] ;
 wire \hash/b_new[27] ;
 wire \hash/b_new[28] ;
 wire \hash/b_new[29] ;
 wire \hash/b_new[2] ;
 wire \hash/b_new[30] ;
 wire \hash/b_new[31] ;
 wire \hash/b_new[3] ;
 wire \hash/b_new[4] ;
 wire \hash/b_new[5] ;
 wire \hash/b_new[6] ;
 wire \hash/b_new[7] ;
 wire \hash/b_new[8] ;
 wire \hash/b_new[9] ;
 wire \hash/c[0] ;
 wire \hash/c[10] ;
 wire \hash/c[11] ;
 wire \hash/c[12] ;
 wire \hash/c[13] ;
 wire \hash/c[14] ;
 wire \hash/c[15] ;
 wire \hash/c[16] ;
 wire \hash/c[17] ;
 wire \hash/c[18] ;
 wire \hash/c[19] ;
 wire \hash/c[1] ;
 wire \hash/c[20] ;
 wire \hash/c[21] ;
 wire \hash/c[22] ;
 wire \hash/c[23] ;
 wire \hash/c[24] ;
 wire \hash/c[25] ;
 wire \hash/c[26] ;
 wire \hash/c[27] ;
 wire \hash/c[28] ;
 wire \hash/c[29] ;
 wire \hash/c[2] ;
 wire \hash/c[30] ;
 wire \hash/c[31] ;
 wire \hash/c[3] ;
 wire \hash/c[4] ;
 wire \hash/c[5] ;
 wire \hash/c[6] ;
 wire \hash/c[7] ;
 wire \hash/c[8] ;
 wire \hash/c[9] ;
 wire \hash/d[0] ;
 wire \hash/d[10] ;
 wire \hash/d[11] ;
 wire \hash/d[12] ;
 wire \hash/d[13] ;
 wire \hash/d[14] ;
 wire \hash/d[15] ;
 wire \hash/d[16] ;
 wire \hash/d[17] ;
 wire \hash/d[18] ;
 wire \hash/d[19] ;
 wire \hash/d[1] ;
 wire \hash/d[20] ;
 wire \hash/d[21] ;
 wire \hash/d[22] ;
 wire \hash/d[23] ;
 wire \hash/d[24] ;
 wire \hash/d[25] ;
 wire \hash/d[26] ;
 wire \hash/d[27] ;
 wire \hash/d[28] ;
 wire \hash/d[29] ;
 wire \hash/d[2] ;
 wire \hash/d[30] ;
 wire \hash/d[31] ;
 wire \hash/d[3] ;
 wire \hash/d[4] ;
 wire \hash/d[5] ;
 wire \hash/d[6] ;
 wire \hash/d[7] ;
 wire \hash/d[8] ;
 wire \hash/d[9] ;
 wire \hash/e[0] ;
 wire \hash/e[10] ;
 wire \hash/e[11] ;
 wire \hash/e[12] ;
 wire \hash/e[13] ;
 wire \hash/e[14] ;
 wire \hash/e[15] ;
 wire \hash/e[16] ;
 wire \hash/e[17] ;
 wire \hash/e[18] ;
 wire \hash/e[19] ;
 wire \hash/e[1] ;
 wire \hash/e[20] ;
 wire \hash/e[21] ;
 wire \hash/e[22] ;
 wire \hash/e[23] ;
 wire \hash/e[24] ;
 wire \hash/e[25] ;
 wire \hash/e[26] ;
 wire \hash/e[27] ;
 wire \hash/e[28] ;
 wire \hash/e[29] ;
 wire \hash/e[2] ;
 wire \hash/e[30] ;
 wire \hash/e[31] ;
 wire \hash/e[3] ;
 wire \hash/e[4] ;
 wire \hash/e[5] ;
 wire \hash/e[6] ;
 wire \hash/e[7] ;
 wire \hash/e[8] ;
 wire \hash/e[9] ;
 wire \hash/e_cap[0] ;
 wire \hash/e_cap[10] ;
 wire \hash/e_cap[11] ;
 wire \hash/e_cap[12] ;
 wire \hash/e_cap[13] ;
 wire \hash/e_cap[14] ;
 wire \hash/e_cap[15] ;
 wire \hash/e_cap[16] ;
 wire \hash/e_cap[17] ;
 wire \hash/e_cap[18] ;
 wire \hash/e_cap[19] ;
 wire \hash/e_cap[1] ;
 wire \hash/e_cap[20] ;
 wire \hash/e_cap[21] ;
 wire \hash/e_cap[22] ;
 wire \hash/e_cap[23] ;
 wire \hash/e_cap[24] ;
 wire \hash/e_cap[25] ;
 wire \hash/e_cap[26] ;
 wire \hash/e_cap[27] ;
 wire \hash/e_cap[28] ;
 wire \hash/e_cap[29] ;
 wire \hash/e_cap[2] ;
 wire \hash/e_cap[30] ;
 wire \hash/e_cap[31] ;
 wire \hash/e_cap[3] ;
 wire \hash/e_cap[4] ;
 wire \hash/e_cap[5] ;
 wire \hash/e_cap[6] ;
 wire \hash/e_cap[7] ;
 wire \hash/e_cap[8] ;
 wire \hash/e_cap[9] ;
 wire \hash/e_new[0] ;
 wire \hash/e_new[10] ;
 wire \hash/e_new[11] ;
 wire \hash/e_new[12] ;
 wire \hash/e_new[13] ;
 wire \hash/e_new[14] ;
 wire \hash/e_new[15] ;
 wire \hash/e_new[16] ;
 wire \hash/e_new[17] ;
 wire \hash/e_new[18] ;
 wire \hash/e_new[19] ;
 wire \hash/e_new[1] ;
 wire \hash/e_new[20] ;
 wire \hash/e_new[21] ;
 wire \hash/e_new[22] ;
 wire \hash/e_new[23] ;
 wire \hash/e_new[24] ;
 wire \hash/e_new[25] ;
 wire \hash/e_new[26] ;
 wire \hash/e_new[27] ;
 wire \hash/e_new[28] ;
 wire \hash/e_new[29] ;
 wire \hash/e_new[2] ;
 wire \hash/e_new[30] ;
 wire \hash/e_new[31] ;
 wire \hash/e_new[3] ;
 wire \hash/e_new[4] ;
 wire \hash/e_new[5] ;
 wire \hash/e_new[6] ;
 wire \hash/e_new[7] ;
 wire \hash/e_new[8] ;
 wire \hash/e_new[9] ;
 wire \hash/f[0] ;
 wire \hash/f[10] ;
 wire \hash/f[11] ;
 wire \hash/f[12] ;
 wire \hash/f[13] ;
 wire \hash/f[14] ;
 wire \hash/f[15] ;
 wire \hash/f[16] ;
 wire \hash/f[17] ;
 wire \hash/f[18] ;
 wire \hash/f[19] ;
 wire \hash/f[1] ;
 wire \hash/f[20] ;
 wire \hash/f[21] ;
 wire \hash/f[22] ;
 wire \hash/f[23] ;
 wire \hash/f[24] ;
 wire \hash/f[25] ;
 wire \hash/f[26] ;
 wire \hash/f[27] ;
 wire \hash/f[28] ;
 wire \hash/f[29] ;
 wire \hash/f[2] ;
 wire \hash/f[30] ;
 wire \hash/f[31] ;
 wire \hash/f[3] ;
 wire \hash/f[4] ;
 wire \hash/f[5] ;
 wire \hash/f[6] ;
 wire \hash/f[7] ;
 wire \hash/f[8] ;
 wire \hash/f[9] ;
 wire \hash/f_cap[0] ;
 wire \hash/f_cap[10] ;
 wire \hash/f_cap[11] ;
 wire \hash/f_cap[12] ;
 wire \hash/f_cap[13] ;
 wire \hash/f_cap[14] ;
 wire \hash/f_cap[15] ;
 wire \hash/f_cap[16] ;
 wire \hash/f_cap[17] ;
 wire \hash/f_cap[18] ;
 wire \hash/f_cap[19] ;
 wire \hash/f_cap[1] ;
 wire \hash/f_cap[20] ;
 wire \hash/f_cap[21] ;
 wire \hash/f_cap[22] ;
 wire \hash/f_cap[23] ;
 wire \hash/f_cap[24] ;
 wire \hash/f_cap[25] ;
 wire \hash/f_cap[26] ;
 wire \hash/f_cap[27] ;
 wire \hash/f_cap[28] ;
 wire \hash/f_cap[29] ;
 wire \hash/f_cap[2] ;
 wire \hash/f_cap[30] ;
 wire \hash/f_cap[31] ;
 wire \hash/f_cap[3] ;
 wire \hash/f_cap[4] ;
 wire \hash/f_cap[5] ;
 wire \hash/f_cap[6] ;
 wire \hash/f_cap[7] ;
 wire \hash/f_cap[8] ;
 wire \hash/f_cap[9] ;
 wire \hash/g[0] ;
 wire \hash/g[10] ;
 wire \hash/g[11] ;
 wire \hash/g[12] ;
 wire \hash/g[13] ;
 wire \hash/g[14] ;
 wire \hash/g[15] ;
 wire \hash/g[16] ;
 wire \hash/g[17] ;
 wire \hash/g[18] ;
 wire \hash/g[19] ;
 wire \hash/g[1] ;
 wire \hash/g[20] ;
 wire \hash/g[21] ;
 wire \hash/g[22] ;
 wire \hash/g[23] ;
 wire \hash/g[24] ;
 wire \hash/g[25] ;
 wire \hash/g[26] ;
 wire \hash/g[27] ;
 wire \hash/g[28] ;
 wire \hash/g[29] ;
 wire \hash/g[2] ;
 wire \hash/g[30] ;
 wire \hash/g[31] ;
 wire \hash/g[3] ;
 wire \hash/g[4] ;
 wire \hash/g[5] ;
 wire \hash/g[6] ;
 wire \hash/g[7] ;
 wire \hash/g[8] ;
 wire \hash/g[9] ;
 wire \hash/h[0] ;
 wire \hash/h[10] ;
 wire \hash/h[11] ;
 wire \hash/h[12] ;
 wire \hash/h[13] ;
 wire \hash/h[14] ;
 wire \hash/h[15] ;
 wire \hash/h[16] ;
 wire \hash/h[17] ;
 wire \hash/h[18] ;
 wire \hash/h[19] ;
 wire \hash/h[1] ;
 wire \hash/h[20] ;
 wire \hash/h[21] ;
 wire \hash/h[22] ;
 wire \hash/h[23] ;
 wire \hash/h[24] ;
 wire \hash/h[25] ;
 wire \hash/h[26] ;
 wire \hash/h[27] ;
 wire \hash/h[28] ;
 wire \hash/h[29] ;
 wire \hash/h[2] ;
 wire \hash/h[30] ;
 wire \hash/h[31] ;
 wire \hash/h[3] ;
 wire \hash/h[4] ;
 wire \hash/h[5] ;
 wire \hash/h[6] ;
 wire \hash/h[7] ;
 wire \hash/h[8] ;
 wire \hash/h[9] ;
 wire \hash/p1[0] ;
 wire \hash/p1[10] ;
 wire \hash/p1[11] ;
 wire \hash/p1[12] ;
 wire \hash/p1[13] ;
 wire \hash/p1[14] ;
 wire \hash/p1[15] ;
 wire \hash/p1[16] ;
 wire \hash/p1[17] ;
 wire \hash/p1[18] ;
 wire \hash/p1[19] ;
 wire \hash/p1[1] ;
 wire \hash/p1[20] ;
 wire \hash/p1[21] ;
 wire \hash/p1[22] ;
 wire \hash/p1[23] ;
 wire \hash/p1[24] ;
 wire \hash/p1[25] ;
 wire \hash/p1[26] ;
 wire \hash/p1[27] ;
 wire \hash/p1[28] ;
 wire \hash/p1[29] ;
 wire \hash/p1[2] ;
 wire \hash/p1[30] ;
 wire \hash/p1[31] ;
 wire \hash/p1[3] ;
 wire \hash/p1[4] ;
 wire \hash/p1[5] ;
 wire \hash/p1[6] ;
 wire \hash/p1[7] ;
 wire \hash/p1[8] ;
 wire \hash/p1[9] ;
 wire \hash/p1_cap[0] ;
 wire \hash/p1_cap[10] ;
 wire \hash/p1_cap[11] ;
 wire \hash/p1_cap[12] ;
 wire \hash/p1_cap[13] ;
 wire \hash/p1_cap[14] ;
 wire \hash/p1_cap[15] ;
 wire \hash/p1_cap[16] ;
 wire \hash/p1_cap[17] ;
 wire \hash/p1_cap[18] ;
 wire \hash/p1_cap[19] ;
 wire \hash/p1_cap[1] ;
 wire \hash/p1_cap[20] ;
 wire \hash/p1_cap[21] ;
 wire \hash/p1_cap[22] ;
 wire \hash/p1_cap[23] ;
 wire \hash/p1_cap[24] ;
 wire \hash/p1_cap[25] ;
 wire \hash/p1_cap[26] ;
 wire \hash/p1_cap[27] ;
 wire \hash/p1_cap[28] ;
 wire \hash/p1_cap[29] ;
 wire \hash/p1_cap[2] ;
 wire \hash/p1_cap[30] ;
 wire \hash/p1_cap[31] ;
 wire \hash/p1_cap[3] ;
 wire \hash/p1_cap[4] ;
 wire \hash/p1_cap[5] ;
 wire \hash/p1_cap[6] ;
 wire \hash/p1_cap[7] ;
 wire \hash/p1_cap[8] ;
 wire \hash/p1_cap[9] ;
 wire \hash/p2[0] ;
 wire \hash/p2[10] ;
 wire \hash/p2[11] ;
 wire \hash/p2[12] ;
 wire \hash/p2[13] ;
 wire \hash/p2[14] ;
 wire \hash/p2[15] ;
 wire \hash/p2[16] ;
 wire \hash/p2[17] ;
 wire \hash/p2[18] ;
 wire \hash/p2[19] ;
 wire \hash/p2[1] ;
 wire \hash/p2[20] ;
 wire \hash/p2[21] ;
 wire \hash/p2[22] ;
 wire \hash/p2[23] ;
 wire \hash/p2[24] ;
 wire \hash/p2[25] ;
 wire \hash/p2[26] ;
 wire \hash/p2[27] ;
 wire \hash/p2[28] ;
 wire \hash/p2[29] ;
 wire \hash/p2[2] ;
 wire \hash/p2[30] ;
 wire \hash/p2[31] ;
 wire \hash/p2[3] ;
 wire \hash/p2[4] ;
 wire \hash/p2[5] ;
 wire \hash/p2[6] ;
 wire \hash/p2[7] ;
 wire \hash/p2[8] ;
 wire \hash/p2[9] ;
 wire \hash/p2_cap[0] ;
 wire \hash/p2_cap[10] ;
 wire \hash/p2_cap[11] ;
 wire \hash/p2_cap[12] ;
 wire \hash/p2_cap[13] ;
 wire \hash/p2_cap[14] ;
 wire \hash/p2_cap[15] ;
 wire \hash/p2_cap[16] ;
 wire \hash/p2_cap[17] ;
 wire \hash/p2_cap[18] ;
 wire \hash/p2_cap[19] ;
 wire \hash/p2_cap[1] ;
 wire \hash/p2_cap[20] ;
 wire \hash/p2_cap[21] ;
 wire \hash/p2_cap[22] ;
 wire \hash/p2_cap[23] ;
 wire \hash/p2_cap[24] ;
 wire \hash/p2_cap[25] ;
 wire \hash/p2_cap[26] ;
 wire \hash/p2_cap[27] ;
 wire \hash/p2_cap[28] ;
 wire \hash/p2_cap[29] ;
 wire \hash/p2_cap[2] ;
 wire \hash/p2_cap[30] ;
 wire \hash/p2_cap[31] ;
 wire \hash/p2_cap[3] ;
 wire \hash/p2_cap[4] ;
 wire \hash/p2_cap[5] ;
 wire \hash/p2_cap[6] ;
 wire \hash/p2_cap[7] ;
 wire \hash/p2_cap[8] ;
 wire \hash/p2_cap[9] ;
 wire \hash/p3[0] ;
 wire \hash/p3[10] ;
 wire \hash/p3[11] ;
 wire \hash/p3[12] ;
 wire \hash/p3[13] ;
 wire \hash/p3[14] ;
 wire \hash/p3[15] ;
 wire \hash/p3[16] ;
 wire \hash/p3[17] ;
 wire \hash/p3[18] ;
 wire \hash/p3[19] ;
 wire \hash/p3[1] ;
 wire \hash/p3[20] ;
 wire \hash/p3[21] ;
 wire \hash/p3[22] ;
 wire \hash/p3[23] ;
 wire \hash/p3[24] ;
 wire \hash/p3[25] ;
 wire \hash/p3[26] ;
 wire \hash/p3[27] ;
 wire \hash/p3[28] ;
 wire \hash/p3[29] ;
 wire \hash/p3[2] ;
 wire \hash/p3[30] ;
 wire \hash/p3[31] ;
 wire \hash/p3[3] ;
 wire \hash/p3[4] ;
 wire \hash/p3[5] ;
 wire \hash/p3[6] ;
 wire \hash/p3[7] ;
 wire \hash/p3[8] ;
 wire \hash/p3[9] ;
 wire \hash/p3_cap[0] ;
 wire \hash/p3_cap[10] ;
 wire \hash/p3_cap[11] ;
 wire \hash/p3_cap[12] ;
 wire \hash/p3_cap[13] ;
 wire \hash/p3_cap[14] ;
 wire \hash/p3_cap[15] ;
 wire \hash/p3_cap[16] ;
 wire \hash/p3_cap[17] ;
 wire \hash/p3_cap[18] ;
 wire \hash/p3_cap[19] ;
 wire \hash/p3_cap[1] ;
 wire \hash/p3_cap[20] ;
 wire \hash/p3_cap[21] ;
 wire \hash/p3_cap[22] ;
 wire \hash/p3_cap[23] ;
 wire \hash/p3_cap[24] ;
 wire \hash/p3_cap[25] ;
 wire \hash/p3_cap[26] ;
 wire \hash/p3_cap[27] ;
 wire \hash/p3_cap[28] ;
 wire \hash/p3_cap[29] ;
 wire \hash/p3_cap[2] ;
 wire \hash/p3_cap[30] ;
 wire \hash/p3_cap[31] ;
 wire \hash/p3_cap[3] ;
 wire \hash/p3_cap[4] ;
 wire \hash/p3_cap[5] ;
 wire \hash/p3_cap[6] ;
 wire \hash/p3_cap[7] ;
 wire \hash/p3_cap[8] ;
 wire \hash/p3_cap[9] ;
 wire \hash/p4[0] ;
 wire \hash/p4[10] ;
 wire \hash/p4[11] ;
 wire \hash/p4[12] ;
 wire \hash/p4[13] ;
 wire \hash/p4[14] ;
 wire \hash/p4[15] ;
 wire \hash/p4[16] ;
 wire \hash/p4[17] ;
 wire \hash/p4[18] ;
 wire \hash/p4[19] ;
 wire \hash/p4[1] ;
 wire \hash/p4[20] ;
 wire \hash/p4[21] ;
 wire \hash/p4[22] ;
 wire \hash/p4[23] ;
 wire \hash/p4[24] ;
 wire \hash/p4[25] ;
 wire \hash/p4[26] ;
 wire \hash/p4[27] ;
 wire \hash/p4[28] ;
 wire \hash/p4[29] ;
 wire \hash/p4[2] ;
 wire \hash/p4[30] ;
 wire \hash/p4[31] ;
 wire \hash/p4[3] ;
 wire \hash/p4[4] ;
 wire \hash/p4[5] ;
 wire \hash/p4[6] ;
 wire \hash/p4[7] ;
 wire \hash/p4[8] ;
 wire \hash/p4[9] ;
 wire \hash/p4_cap[0] ;
 wire \hash/p4_cap[10] ;
 wire \hash/p4_cap[11] ;
 wire \hash/p4_cap[12] ;
 wire \hash/p4_cap[13] ;
 wire \hash/p4_cap[14] ;
 wire \hash/p4_cap[15] ;
 wire \hash/p4_cap[16] ;
 wire \hash/p4_cap[17] ;
 wire \hash/p4_cap[18] ;
 wire \hash/p4_cap[19] ;
 wire \hash/p4_cap[1] ;
 wire \hash/p4_cap[20] ;
 wire \hash/p4_cap[21] ;
 wire \hash/p4_cap[22] ;
 wire \hash/p4_cap[23] ;
 wire \hash/p4_cap[24] ;
 wire \hash/p4_cap[25] ;
 wire \hash/p4_cap[26] ;
 wire \hash/p4_cap[27] ;
 wire \hash/p4_cap[28] ;
 wire \hash/p4_cap[29] ;
 wire \hash/p4_cap[2] ;
 wire \hash/p4_cap[30] ;
 wire \hash/p4_cap[31] ;
 wire \hash/p4_cap[3] ;
 wire \hash/p4_cap[4] ;
 wire \hash/p4_cap[5] ;
 wire \hash/p4_cap[6] ;
 wire \hash/p4_cap[7] ;
 wire \hash/p4_cap[8] ;
 wire \hash/p4_cap[9] ;
 wire \hash/p5[0] ;
 wire \hash/p5[10] ;
 wire \hash/p5[11] ;
 wire \hash/p5[12] ;
 wire \hash/p5[13] ;
 wire \hash/p5[14] ;
 wire \hash/p5[15] ;
 wire \hash/p5[16] ;
 wire \hash/p5[17] ;
 wire \hash/p5[18] ;
 wire \hash/p5[19] ;
 wire \hash/p5[1] ;
 wire \hash/p5[20] ;
 wire \hash/p5[21] ;
 wire \hash/p5[22] ;
 wire \hash/p5[23] ;
 wire \hash/p5[24] ;
 wire \hash/p5[25] ;
 wire \hash/p5[26] ;
 wire \hash/p5[27] ;
 wire \hash/p5[28] ;
 wire \hash/p5[29] ;
 wire \hash/p5[2] ;
 wire \hash/p5[30] ;
 wire \hash/p5[31] ;
 wire \hash/p5[3] ;
 wire \hash/p5[4] ;
 wire \hash/p5[5] ;
 wire \hash/p5[6] ;
 wire \hash/p5[7] ;
 wire \hash/p5[8] ;
 wire \hash/p5[9] ;
 wire \hash/p5_cap[0] ;
 wire \hash/p5_cap[10] ;
 wire \hash/p5_cap[11] ;
 wire \hash/p5_cap[12] ;
 wire \hash/p5_cap[13] ;
 wire \hash/p5_cap[14] ;
 wire \hash/p5_cap[15] ;
 wire \hash/p5_cap[16] ;
 wire \hash/p5_cap[17] ;
 wire \hash/p5_cap[18] ;
 wire \hash/p5_cap[19] ;
 wire \hash/p5_cap[1] ;
 wire \hash/p5_cap[20] ;
 wire \hash/p5_cap[21] ;
 wire \hash/p5_cap[22] ;
 wire \hash/p5_cap[23] ;
 wire \hash/p5_cap[24] ;
 wire \hash/p5_cap[25] ;
 wire \hash/p5_cap[26] ;
 wire \hash/p5_cap[27] ;
 wire \hash/p5_cap[28] ;
 wire \hash/p5_cap[29] ;
 wire \hash/p5_cap[2] ;
 wire \hash/p5_cap[30] ;
 wire \hash/p5_cap[31] ;
 wire \hash/p5_cap[3] ;
 wire \hash/p5_cap[4] ;
 wire \hash/p5_cap[5] ;
 wire \hash/p5_cap[6] ;
 wire \hash/p5_cap[7] ;
 wire \hash/p5_cap[8] ;
 wire \hash/p5_cap[9] ;
 wire \hash/CA1/_0000_ ;
 wire \hash/CA1/_0001_ ;
 wire \hash/CA1/_0002_ ;
 wire \hash/CA1/_0003_ ;
 wire \hash/CA1/_0004_ ;
 wire \hash/CA1/_0005_ ;
 wire \hash/CA1/_0006_ ;
 wire \hash/CA1/_0007_ ;
 wire \hash/CA1/_0008_ ;
 wire \hash/CA1/_0009_ ;
 wire \hash/CA1/_0010_ ;
 wire \hash/CA1/_0011_ ;
 wire \hash/CA1/_0012_ ;
 wire \hash/CA1/_0013_ ;
 wire \hash/CA1/_0014_ ;
 wire \hash/CA1/_0015_ ;
 wire \hash/CA1/_0016_ ;
 wire \hash/CA1/_0017_ ;
 wire \hash/CA1/_0018_ ;
 wire \hash/CA1/_0019_ ;
 wire \hash/CA1/_0020_ ;
 wire \hash/CA1/_0021_ ;
 wire \hash/CA1/_0022_ ;
 wire \hash/CA1/_0023_ ;
 wire \hash/CA1/_0024_ ;
 wire \hash/CA1/_0025_ ;
 wire \hash/CA1/_0026_ ;
 wire \hash/CA1/_0027_ ;
 wire \hash/CA1/_0028_ ;
 wire \hash/CA1/_0029_ ;
 wire \hash/CA1/_0030_ ;
 wire \hash/CA1/_0031_ ;
 wire \hash/CA1/_0032_ ;
 wire \hash/CA1/_0033_ ;
 wire \hash/CA1/_0034_ ;
 wire \hash/CA1/_0035_ ;
 wire \hash/CA1/_0036_ ;
 wire \hash/CA1/_0037_ ;
 wire \hash/CA1/_0038_ ;
 wire \hash/CA1/_0039_ ;
 wire \hash/CA1/_0040_ ;
 wire \hash/CA1/_0041_ ;
 wire \hash/CA1/_0042_ ;
 wire \hash/CA1/_0043_ ;
 wire \hash/CA1/_0044_ ;
 wire \hash/CA1/_0045_ ;
 wire \hash/CA1/_0046_ ;
 wire \hash/CA1/_0047_ ;
 wire \hash/CA1/_0048_ ;
 wire \hash/CA1/_0049_ ;
 wire \hash/CA1/_0050_ ;
 wire \hash/CA1/_0051_ ;
 wire \hash/CA1/_0052_ ;
 wire \hash/CA1/_0053_ ;
 wire \hash/CA1/_0054_ ;
 wire \hash/CA1/_0055_ ;
 wire \hash/CA1/_0056_ ;
 wire \hash/CA1/_0057_ ;
 wire \hash/CA1/_0058_ ;
 wire \hash/CA1/_0059_ ;
 wire \hash/CA1/_0060_ ;
 wire \hash/CA1/_0061_ ;
 wire \hash/CA1/_0062_ ;
 wire \hash/CA1/_0063_ ;
 wire \hash/CA1/_0064_ ;
 wire \hash/CA1/_0065_ ;
 wire \hash/CA1/_0066_ ;
 wire \hash/CA1/_0067_ ;
 wire \hash/CA1/_0068_ ;
 wire \hash/CA1/_0069_ ;
 wire \hash/CA1/_0070_ ;
 wire \hash/CA1/_0071_ ;
 wire \hash/CA1/_0073_ ;
 wire \hash/CA1/_0074_ ;
 wire \hash/CA1/_0075_ ;
 wire \hash/CA1/_0076_ ;
 wire \hash/CA1/_0077_ ;
 wire \hash/CA1/_0078_ ;
 wire \hash/CA1/_0079_ ;
 wire \hash/CA1/_0080_ ;
 wire \hash/CA1/_0081_ ;
 wire \hash/CA1/_0082_ ;
 wire \hash/CA1/_0083_ ;
 wire \hash/CA1/_0084_ ;
 wire \hash/CA1/_0085_ ;
 wire \hash/CA1/_0086_ ;
 wire \hash/CA1/_0087_ ;
 wire \hash/CA1/_0088_ ;
 wire \hash/CA1/_0090_ ;
 wire \hash/CA1/_0091_ ;
 wire \hash/CA1/_0092_ ;
 wire \hash/CA1/_0093_ ;
 wire \hash/CA1/_0094_ ;
 wire \hash/CA1/_0095_ ;
 wire \hash/CA1/_0096_ ;
 wire \hash/CA1/_0097_ ;
 wire \hash/CA1/_0098_ ;
 wire \hash/CA1/_0099_ ;
 wire \hash/CA1/_0100_ ;
 wire \hash/CA1/_0101_ ;
 wire \hash/CA1/_0102_ ;
 wire \hash/CA1/_0103_ ;
 wire \hash/CA1/_0104_ ;
 wire \hash/CA1/_0105_ ;
 wire \hash/CA1/_0106_ ;
 wire \hash/CA1/_0107_ ;
 wire \hash/CA1/_0108_ ;
 wire \hash/CA1/_0109_ ;
 wire \hash/CA1/_0110_ ;
 wire \hash/CA1/_0111_ ;
 wire \hash/CA1/_0112_ ;
 wire \hash/CA1/_0113_ ;
 wire \hash/CA1/_0114_ ;
 wire \hash/CA1/_0115_ ;
 wire \hash/CA1/_0116_ ;
 wire \hash/CA1/_0117_ ;
 wire \hash/CA1/_0118_ ;
 wire \hash/CA1/_0120_ ;
 wire \hash/CA1/_0121_ ;
 wire \hash/CA1/_0122_ ;
 wire \hash/CA1/_0123_ ;
 wire \hash/CA1/_0124_ ;
 wire \hash/CA1/_0125_ ;
 wire \hash/CA1/_0126_ ;
 wire \hash/CA1/_0127_ ;
 wire \hash/CA1/_0128_ ;
 wire \hash/CA1/_0129_ ;
 wire \hash/CA1/_0130_ ;
 wire \hash/CA1/_0131_ ;
 wire \hash/CA1/_0132_ ;
 wire \hash/CA1/_0133_ ;
 wire \hash/CA1/_0134_ ;
 wire \hash/CA1/_0135_ ;
 wire \hash/CA1/_0136_ ;
 wire \hash/CA1/_0137_ ;
 wire \hash/CA1/_0138_ ;
 wire \hash/CA1/_0139_ ;
 wire \hash/CA1/_0141_ ;
 wire \hash/CA1/_0142_ ;
 wire \hash/CA1/_0143_ ;
 wire \hash/CA1/_0144_ ;
 wire \hash/CA1/_0145_ ;
 wire \hash/CA1/_0146_ ;
 wire \hash/CA1/_0147_ ;
 wire \hash/CA1/_0148_ ;
 wire \hash/CA1/_0149_ ;
 wire \hash/CA1/_0151_ ;
 wire \hash/CA1/_0152_ ;
 wire \hash/CA1/_0153_ ;
 wire \hash/CA1/_0154_ ;
 wire \hash/CA1/_0156_ ;
 wire \hash/CA1/_0157_ ;
 wire \hash/CA1/_0158_ ;
 wire \hash/CA1/_0159_ ;
 wire \hash/CA1/_0160_ ;
 wire \hash/CA1/_0161_ ;
 wire \hash/CA1/_0162_ ;
 wire \hash/CA1/_0163_ ;
 wire \hash/CA1/_0164_ ;
 wire \hash/CA1/_0165_ ;
 wire \hash/CA1/_0166_ ;
 wire \hash/CA1/_0167_ ;
 wire \hash/CA1/_0168_ ;
 wire \hash/CA1/_0169_ ;
 wire \hash/CA1/_0170_ ;
 wire \hash/CA1/_0171_ ;
 wire \hash/CA1/_0172_ ;
 wire \hash/CA1/_0173_ ;
 wire \hash/CA1/_0174_ ;
 wire \hash/CA1/_0175_ ;
 wire \hash/CA1/_0176_ ;
 wire \hash/CA1/_0177_ ;
 wire \hash/CA1/_0178_ ;
 wire \hash/CA1/_0179_ ;
 wire \hash/CA1/_0180_ ;
 wire \hash/CA1/_0181_ ;
 wire \hash/CA1/_0182_ ;
 wire \hash/CA1/_0183_ ;
 wire \hash/CA1/_0184_ ;
 wire \hash/CA1/_0185_ ;
 wire \hash/CA1/_0187_ ;
 wire \hash/CA1/_0188_ ;
 wire \hash/CA1/_0189_ ;
 wire \hash/CA1/_0190_ ;
 wire \hash/CA1/_0191_ ;
 wire \hash/CA1/_0192_ ;
 wire \hash/CA1/_0193_ ;
 wire \hash/CA1/_0194_ ;
 wire \hash/CA1/_0195_ ;
 wire \hash/CA1/_0196_ ;
 wire \hash/CA1/_0197_ ;
 wire \hash/CA1/_0198_ ;
 wire \hash/CA1/_0199_ ;
 wire \hash/CA1/_0200_ ;
 wire \hash/CA1/_0201_ ;
 wire \hash/CA1/_0202_ ;
 wire \hash/CA1/_0203_ ;
 wire \hash/CA1/_0204_ ;
 wire \hash/CA1/_0205_ ;
 wire \hash/CA1/_0206_ ;
 wire \hash/CA1/_0208_ ;
 wire \hash/CA1/_0209_ ;
 wire \hash/CA1/_0210_ ;
 wire \hash/CA1/_0211_ ;
 wire \hash/CA1/_0212_ ;
 wire \hash/CA1/_0213_ ;
 wire \hash/CA1/_0214_ ;
 wire \hash/CA1/_0215_ ;
 wire \hash/CA1/_0217_ ;
 wire \hash/CA1/_0218_ ;
 wire \hash/CA1/_0219_ ;
 wire \hash/CA1/_0220_ ;
 wire \hash/CA1/_0221_ ;
 wire \hash/CA1/_0222_ ;
 wire \hash/CA1/_0223_ ;
 wire \hash/CA1/_0224_ ;
 wire \hash/CA1/_0225_ ;
 wire \hash/CA1/_0226_ ;
 wire \hash/CA1/_0227_ ;
 wire \hash/CA1/_0228_ ;
 wire \hash/CA1/_0229_ ;
 wire \hash/CA1/_0230_ ;
 wire \hash/CA1/_0231_ ;
 wire \hash/CA1/_0232_ ;
 wire \hash/CA1/_0233_ ;
 wire \hash/CA1/_0234_ ;
 wire \hash/CA1/_0235_ ;
 wire \hash/CA1/_0236_ ;
 wire \hash/CA1/_0237_ ;
 wire \hash/CA1/_0238_ ;
 wire \hash/CA1/_0239_ ;
 wire \hash/CA1/_0240_ ;
 wire \hash/CA1/_0241_ ;
 wire \hash/CA1/_0242_ ;
 wire \hash/CA1/_0243_ ;
 wire \hash/CA1/_0244_ ;
 wire \hash/CA1/_0245_ ;
 wire \hash/CA1/_0246_ ;
 wire \hash/CA1/_0247_ ;
 wire \hash/CA1/_0248_ ;
 wire \hash/CA1/_0249_ ;
 wire \hash/CA1/_0250_ ;
 wire \hash/CA1/_0251_ ;
 wire \hash/CA1/_0252_ ;
 wire \hash/CA1/_0253_ ;
 wire \hash/CA1/_0254_ ;
 wire \hash/CA1/_0255_ ;
 wire \hash/CA1/_0256_ ;
 wire \hash/CA1/_0257_ ;
 wire \hash/CA1/_0258_ ;
 wire \hash/CA1/_0259_ ;
 wire \hash/CA1/_0260_ ;
 wire \hash/CA1/_0261_ ;
 wire \hash/CA1/_0262_ ;
 wire \hash/CA1/_0263_ ;
 wire \hash/CA1/_0264_ ;
 wire \hash/CA1/_0265_ ;
 wire \hash/CA1/_0266_ ;
 wire \hash/CA1/_0267_ ;
 wire \hash/CA1/_0268_ ;
 wire \hash/CA1/_0269_ ;
 wire \hash/CA1/_0270_ ;
 wire \hash/CA1/_0271_ ;
 wire \hash/CA1/_0272_ ;
 wire \hash/CA1/_0273_ ;
 wire \hash/CA1/_0274_ ;
 wire \hash/CA1/_0275_ ;
 wire \hash/CA1/_0276_ ;
 wire \hash/CA1/_0277_ ;
 wire \hash/CA1/_0278_ ;
 wire \hash/CA1/_0279_ ;
 wire \hash/CA1/_0280_ ;
 wire \hash/CA1/_0281_ ;
 wire \hash/CA1/_0282_ ;
 wire \hash/CA1/_0283_ ;
 wire \hash/CA1/_0284_ ;
 wire \hash/CA1/_0285_ ;
 wire \hash/CA1/_0286_ ;
 wire \hash/CA1/_0287_ ;
 wire \hash/CA1/_0288_ ;
 wire \hash/CA1/_0289_ ;
 wire \hash/CA1/_0290_ ;
 wire \hash/CA1/_0291_ ;
 wire \hash/CA1/_0292_ ;
 wire \hash/CA1/_0293_ ;
 wire \hash/CA1/_0294_ ;
 wire \hash/CA1/_0295_ ;
 wire \hash/CA1/_0296_ ;
 wire \hash/CA1/_0297_ ;
 wire \hash/CA1/_0298_ ;
 wire \hash/CA1/_0299_ ;
 wire \hash/CA1/_0300_ ;
 wire \hash/CA1/_0301_ ;
 wire \hash/CA1/_0302_ ;
 wire \hash/CA1/_0303_ ;
 wire \hash/CA1/_0304_ ;
 wire \hash/CA1/_0305_ ;
 wire \hash/CA1/_0306_ ;
 wire \hash/CA1/_0307_ ;
 wire \hash/CA1/_0308_ ;
 wire \hash/CA1/_0309_ ;
 wire \hash/CA1/_0310_ ;
 wire \hash/CA1/_0311_ ;
 wire \hash/CA1/_0312_ ;
 wire \hash/CA1/_0313_ ;
 wire \hash/CA1/_0314_ ;
 wire \hash/CA1/_0315_ ;
 wire \hash/CA1/_0316_ ;
 wire \hash/CA1/_0317_ ;
 wire \hash/CA1/_0318_ ;
 wire \hash/CA1/_0319_ ;
 wire \hash/CA1/_0320_ ;
 wire \hash/CA1/_0321_ ;
 wire \hash/CA1/_0322_ ;
 wire \hash/CA1/_0323_ ;
 wire \hash/CA1/_0324_ ;
 wire \hash/CA1/_0325_ ;
 wire \hash/CA1/_0326_ ;
 wire \hash/CA1/_0327_ ;
 wire \hash/CA1/_0328_ ;
 wire \hash/CA1/_0329_ ;
 wire \hash/CA1/_0330_ ;
 wire \hash/CA1/_0331_ ;
 wire \hash/CA1/_0332_ ;
 wire \hash/CA1/_0333_ ;
 wire \hash/CA1/_0334_ ;
 wire \hash/CA1/_0335_ ;
 wire \hash/CA1/_0336_ ;
 wire \hash/CA1/_0337_ ;
 wire \hash/CA1/_0338_ ;
 wire \hash/CA1/_0339_ ;
 wire \hash/CA1/_0340_ ;
 wire \hash/CA1/_0341_ ;
 wire \hash/CA1/_0342_ ;
 wire \hash/CA1/_0343_ ;
 wire \hash/CA1/_0344_ ;
 wire \hash/CA1/_0345_ ;
 wire \hash/CA1/_0346_ ;
 wire \hash/CA1/_0347_ ;
 wire \hash/CA1/_0348_ ;
 wire \hash/CA1/_0349_ ;
 wire \hash/CA1/_0350_ ;
 wire \hash/CA1/_0351_ ;
 wire \hash/CA1/_0352_ ;
 wire \hash/CA1/_0353_ ;
 wire \hash/CA1/_0354_ ;
 wire \hash/CA1/_0355_ ;
 wire \hash/CA1/_0356_ ;
 wire \hash/CA1/_0357_ ;
 wire \hash/CA1/_0358_ ;
 wire \hash/CA1/_0359_ ;
 wire \hash/CA1/_0360_ ;
 wire \hash/CA1/_0361_ ;
 wire \hash/CA1/_0362_ ;
 wire \hash/CA1/_0363_ ;
 wire \hash/CA1/_0364_ ;
 wire \hash/CA1/_0365_ ;
 wire \hash/CA1/_0366_ ;
 wire \hash/CA1/_0367_ ;
 wire \hash/CA1/_0368_ ;
 wire \hash/CA1/_0369_ ;
 wire \hash/CA1/_0370_ ;
 wire \hash/CA1/_0371_ ;
 wire \hash/CA1/_0372_ ;
 wire \hash/CA1/_0373_ ;
 wire \hash/CA1/_0374_ ;
 wire \hash/CA1/_0375_ ;
 wire \hash/CA1/_0376_ ;
 wire \hash/CA1/_0377_ ;
 wire \hash/CA1/_0378_ ;
 wire \hash/CA1/_0379_ ;
 wire \hash/CA1/_0380_ ;
 wire \hash/CA1/_0381_ ;
 wire \hash/CA1/_0382_ ;
 wire \hash/CA1/_0383_ ;
 wire \hash/CA1/_0384_ ;
 wire \hash/CA1/_0385_ ;
 wire \hash/CA1/_0386_ ;
 wire \hash/CA1/_0387_ ;
 wire \hash/CA1/_0388_ ;
 wire \hash/CA1/_0389_ ;
 wire \hash/CA1/_0390_ ;
 wire \hash/CA1/_0391_ ;
 wire \hash/CA1/_0392_ ;
 wire \hash/CA1/_0393_ ;
 wire \hash/CA1/_0394_ ;
 wire \hash/CA1/_0395_ ;
 wire \hash/CA1/_0396_ ;
 wire \hash/CA1/_0397_ ;
 wire \hash/CA1/_0398_ ;
 wire \hash/CA1/_0399_ ;
 wire \hash/CA1/_0400_ ;
 wire \hash/CA1/_0401_ ;
 wire \hash/CA1/_0402_ ;
 wire \hash/CA1/_0403_ ;
 wire \hash/CA1/_0404_ ;
 wire \hash/CA1/_0405_ ;
 wire \hash/CA1/_0406_ ;
 wire \hash/CA1/_0407_ ;
 wire \hash/CA1/_0408_ ;
 wire \hash/CA1/_0409_ ;
 wire \hash/CA1/_0410_ ;
 wire \hash/CA1/_0411_ ;
 wire \hash/CA1/_0412_ ;
 wire \hash/CA1/_0413_ ;
 wire \hash/CA1/_0414_ ;
 wire \hash/CA1/_0415_ ;
 wire \hash/CA1/_0416_ ;
 wire \hash/CA1/_0417_ ;
 wire \hash/CA1/_0418_ ;
 wire \hash/CA1/_0419_ ;
 wire \hash/CA1/_0420_ ;
 wire \hash/CA1/_0421_ ;
 wire \hash/CA1/_0422_ ;
 wire \hash/CA1/_0423_ ;
 wire \hash/CA1/_0424_ ;
 wire \hash/CA1/_0425_ ;
 wire \hash/CA1/_0426_ ;
 wire \hash/CA1/_0427_ ;
 wire \hash/CA1/_0428_ ;
 wire \hash/CA1/_0429_ ;
 wire \hash/CA1/_0430_ ;
 wire \hash/CA1/_0431_ ;
 wire \hash/CA1/_0432_ ;
 wire \hash/CA1/_0433_ ;
 wire \hash/CA1/_0434_ ;
 wire \hash/CA1/_0435_ ;
 wire \hash/CA1/_0436_ ;
 wire \hash/CA1/_0437_ ;
 wire \hash/CA1/_0438_ ;
 wire \hash/CA1/_0439_ ;
 wire \hash/CA1/_0440_ ;
 wire \hash/CA1/_0441_ ;
 wire \hash/CA1/_0442_ ;
 wire \hash/CA1/_0443_ ;
 wire \hash/CA1/_0444_ ;
 wire \hash/CA1/_0445_ ;
 wire \hash/CA1/_0446_ ;
 wire \hash/CA1/_0447_ ;
 wire \hash/CA1/_0448_ ;
 wire \hash/CA1/_0449_ ;
 wire \hash/CA1/_0450_ ;
 wire \hash/CA1/_0451_ ;
 wire \hash/CA1/_0452_ ;
 wire \hash/CA1/_0453_ ;
 wire \hash/CA1/_0454_ ;
 wire \hash/CA1/_0455_ ;
 wire \hash/CA1/_0456_ ;
 wire \hash/CA1/_0457_ ;
 wire \hash/CA1/_0458_ ;
 wire \hash/CA1/_0459_ ;
 wire \hash/CA1/_0460_ ;
 wire \hash/CA1/_0461_ ;
 wire \hash/CA1/_0462_ ;
 wire \hash/CA1/_0463_ ;
 wire \hash/CA1/_0464_ ;
 wire \hash/CA1/_0465_ ;
 wire \hash/CA1/_0466_ ;
 wire \hash/CA1/_0467_ ;
 wire \hash/CA1/_0468_ ;
 wire \hash/CA1/_0469_ ;
 wire \hash/CA1/_0470_ ;
 wire \hash/CA1/_0471_ ;
 wire \hash/CA1/_0472_ ;
 wire \hash/CA1/_0473_ ;
 wire \hash/CA1/_0474_ ;
 wire \hash/CA1/_0475_ ;
 wire \hash/CA1/_0476_ ;
 wire \hash/CA1/_0477_ ;
 wire \hash/CA1/_0478_ ;
 wire \hash/CA1/_0479_ ;
 wire \hash/CA1/_0480_ ;
 wire \hash/CA1/_0481_ ;
 wire \hash/CA1/_0482_ ;
 wire \hash/CA1/_0483_ ;
 wire \hash/CA1/_0484_ ;
 wire \hash/CA1/_0485_ ;
 wire \hash/CA1/_0486_ ;
 wire \hash/CA1/_0487_ ;
 wire \hash/CA1/_0488_ ;
 wire \hash/CA1/_0489_ ;
 wire \hash/CA1/_0490_ ;
 wire \hash/CA1/_0491_ ;
 wire \hash/CA1/_0492_ ;
 wire \hash/CA1/_0493_ ;
 wire \hash/CA1/_0494_ ;
 wire \hash/CA1/_0495_ ;
 wire \hash/CA1/_0496_ ;
 wire \hash/CA1/_0497_ ;
 wire \hash/CA1/_0498_ ;
 wire \hash/CA1/_0499_ ;
 wire \hash/CA1/_0500_ ;
 wire \hash/CA1/_0501_ ;
 wire \hash/CA1/_0502_ ;
 wire \hash/CA1/_0503_ ;
 wire \hash/CA1/_0504_ ;
 wire \hash/CA1/_0505_ ;
 wire \hash/CA1/_0506_ ;
 wire \hash/CA1/_0507_ ;
 wire \hash/CA1/_0508_ ;
 wire \hash/CA1/_0509_ ;
 wire \hash/CA1/_0510_ ;
 wire \hash/CA1/_0511_ ;
 wire \hash/CA1/_0512_ ;
 wire \hash/CA1/_0513_ ;
 wire \hash/CA1/_0514_ ;
 wire \hash/CA1/_0515_ ;
 wire \hash/CA1/_0516_ ;
 wire \hash/CA1/_0517_ ;
 wire \hash/CA1/_0518_ ;
 wire \hash/CA1/_0519_ ;
 wire \hash/CA1/_0520_ ;
 wire \hash/CA1/_0521_ ;
 wire \hash/CA1/_0522_ ;
 wire \hash/CA1/_0523_ ;
 wire \hash/CA1/_0524_ ;
 wire \hash/CA1/_0525_ ;
 wire \hash/CA1/_0526_ ;
 wire \hash/CA1/_0527_ ;
 wire \hash/CA1/_0528_ ;
 wire \hash/CA1/_0529_ ;
 wire \hash/CA1/_0530_ ;
 wire \hash/CA1/_0531_ ;
 wire \hash/CA1/_0532_ ;
 wire \hash/CA1/_0533_ ;
 wire \hash/CA1/_0534_ ;
 wire \hash/CA1/_0535_ ;
 wire \hash/CA1/_0536_ ;
 wire \hash/CA1/_0537_ ;
 wire \hash/CA1/_0538_ ;
 wire \hash/CA1/_0539_ ;
 wire \hash/CA1/_0540_ ;
 wire \hash/CA1/_0541_ ;
 wire \hash/CA1/_0542_ ;
 wire \hash/CA1/_0543_ ;
 wire \hash/CA1/_0544_ ;
 wire \hash/CA1/_0545_ ;
 wire \hash/CA1/_0546_ ;
 wire \hash/CA1/_0547_ ;
 wire \hash/CA1/_0548_ ;
 wire \hash/CA1/_0549_ ;
 wire \hash/CA1/_0550_ ;
 wire \hash/CA1/_0551_ ;
 wire \hash/CA1/_0552_ ;
 wire \hash/CA1/_0553_ ;
 wire \hash/CA1/_0554_ ;
 wire \hash/CA1/_0555_ ;
 wire \hash/CA1/_0556_ ;
 wire \hash/CA1/_0557_ ;
 wire \hash/CA1/_0558_ ;
 wire \hash/CA1/_0559_ ;
 wire \hash/CA1/_0560_ ;
 wire \hash/CA1/_0561_ ;
 wire \hash/CA1/_0562_ ;
 wire \hash/CA1/_0563_ ;
 wire \hash/CA1/_0564_ ;
 wire \hash/CA1/_0565_ ;
 wire \hash/CA1/_0566_ ;
 wire \hash/CA1/_0567_ ;
 wire \hash/CA1/_0568_ ;
 wire \hash/CA1/_0569_ ;
 wire \hash/CA1/_0570_ ;
 wire \hash/CA1/_0571_ ;
 wire \hash/CA1/_0572_ ;
 wire \hash/CA1/_0573_ ;
 wire \hash/CA1/_0574_ ;
 wire \hash/CA1/_0575_ ;
 wire \hash/CA1/_0576_ ;
 wire \hash/CA1/_0577_ ;
 wire \hash/CA1/_0578_ ;
 wire \hash/CA1/_0579_ ;
 wire \hash/CA1/_0580_ ;
 wire \hash/CA1/_0581_ ;
 wire \hash/CA1/_0582_ ;
 wire \hash/CA1/_0583_ ;
 wire \hash/CA1/_0584_ ;
 wire \hash/CA1/_0585_ ;
 wire \hash/CA1/_0586_ ;
 wire \hash/CA1/_0587_ ;
 wire \hash/CA1/_0588_ ;
 wire \hash/CA1/_0589_ ;
 wire \hash/CA1/_0590_ ;
 wire \hash/CA1/_0591_ ;
 wire \hash/CA1/_0592_ ;
 wire \hash/CA1/_0593_ ;
 wire \hash/CA1/_0594_ ;
 wire \hash/CA1/_0595_ ;
 wire \hash/CA1/_0596_ ;
 wire \hash/CA1/_0597_ ;
 wire \hash/CA1/_0598_ ;
 wire \hash/CA1/_0599_ ;
 wire \hash/CA1/_0600_ ;
 wire \hash/CA1/_0601_ ;
 wire \hash/CA1/_0602_ ;
 wire \hash/CA1/_0603_ ;
 wire \hash/CA1/_0604_ ;
 wire \hash/CA1/_0605_ ;
 wire \hash/CA1/_0606_ ;
 wire \hash/CA1/_0607_ ;
 wire \hash/CA1/_0608_ ;
 wire \hash/CA1/_0609_ ;
 wire \hash/CA1/_0610_ ;
 wire \hash/CA1/_0611_ ;
 wire \hash/CA1/_0613_ ;
 wire \hash/CA1/_0614_ ;
 wire \hash/CA1/_0615_ ;
 wire \hash/CA1/_0616_ ;
 wire \hash/CA1/_0617_ ;
 wire \hash/CA1/_0618_ ;
 wire \hash/CA1/_0619_ ;
 wire \hash/CA1/_0620_ ;
 wire \hash/CA1/_0621_ ;
 wire \hash/CA1/_0622_ ;
 wire \hash/CA1/_0623_ ;
 wire \hash/CA1/_0624_ ;
 wire \hash/CA1/_0625_ ;
 wire \hash/CA1/_0626_ ;
 wire \hash/CA1/_0627_ ;
 wire \hash/CA1/_0628_ ;
 wire \hash/CA1/_0629_ ;
 wire \hash/CA1/_0630_ ;
 wire \hash/CA1/_0631_ ;
 wire \hash/CA1/_0632_ ;
 wire \hash/CA1/_0633_ ;
 wire \hash/CA1/_0634_ ;
 wire \hash/CA1/_0635_ ;
 wire \hash/CA1/_0636_ ;
 wire \hash/CA1/_0637_ ;
 wire \hash/CA1/_0638_ ;
 wire \hash/CA1/_0639_ ;
 wire \hash/CA1/_0640_ ;
 wire \hash/CA1/_0641_ ;
 wire \hash/CA1/_0642_ ;
 wire \hash/CA1/_0643_ ;
 wire \hash/CA1/_0644_ ;
 wire \hash/CA1/_0645_ ;
 wire \hash/CA1/_0646_ ;
 wire \hash/CA1/_0647_ ;
 wire \hash/CA1/_0648_ ;
 wire \hash/CA1/_0649_ ;
 wire \hash/CA1/_0650_ ;
 wire \hash/CA1/_0651_ ;
 wire \hash/CA1/_0652_ ;
 wire \hash/CA1/_0653_ ;
 wire \hash/CA1/_0654_ ;
 wire \hash/CA1/_0655_ ;
 wire \hash/CA1/_0656_ ;
 wire \hash/CA1/_0657_ ;
 wire \hash/CA1/_0658_ ;
 wire \hash/CA1/_0659_ ;
 wire \hash/CA1/_0660_ ;
 wire \hash/CA1/_0661_ ;
 wire \hash/CA1/_0662_ ;
 wire \hash/CA1/_0663_ ;
 wire \hash/CA1/_0664_ ;
 wire \hash/CA1/_0665_ ;
 wire \hash/CA1/_0666_ ;
 wire \hash/CA1/_0667_ ;
 wire \hash/CA1/_0668_ ;
 wire \hash/CA1/_0669_ ;
 wire \hash/CA1/_0670_ ;
 wire \hash/CA1/_0671_ ;
 wire \hash/CA1/_0672_ ;
 wire \hash/CA1/_0673_ ;
 wire \hash/CA1/_0674_ ;
 wire \hash/CA1/_0675_ ;
 wire \hash/CA1/_0676_ ;
 wire \hash/CA1/_0677_ ;
 wire \hash/CA1/_0678_ ;
 wire \hash/CA1/_0679_ ;
 wire \hash/CA1/_0680_ ;
 wire \hash/CA1/_0681_ ;
 wire \hash/CA1/_0682_ ;
 wire \hash/CA1/_0683_ ;
 wire \hash/CA1/_0684_ ;
 wire \hash/CA1/_0685_ ;
 wire \hash/CA1/_0686_ ;
 wire \hash/CA1/_0687_ ;
 wire \hash/CA1/_0688_ ;
 wire \hash/CA1/_0689_ ;
 wire \hash/CA1/_0690_ ;
 wire \hash/CA1/_0691_ ;
 wire \hash/CA1/_0692_ ;
 wire \hash/CA1/_0694_ ;
 wire \hash/CA1/_0695_ ;
 wire \hash/CA1/_0696_ ;
 wire \hash/CA1/_0697_ ;
 wire \hash/CA1/_0698_ ;
 wire \hash/CA1/_0699_ ;
 wire \hash/CA1/_0700_ ;
 wire \hash/CA1/_0701_ ;
 wire \hash/CA1/_0702_ ;
 wire \hash/CA1/_0703_ ;
 wire \hash/CA1/_0704_ ;
 wire \hash/CA1/_0705_ ;
 wire \hash/CA1/_0706_ ;
 wire \hash/CA1/_0707_ ;
 wire \hash/CA1/_0708_ ;
 wire \hash/CA1/_0709_ ;
 wire \hash/CA1/_0710_ ;
 wire \hash/CA1/_0711_ ;
 wire \hash/CA1/_0712_ ;
 wire \hash/CA1/_0713_ ;
 wire \hash/CA1/_0714_ ;
 wire \hash/CA1/_0715_ ;
 wire \hash/CA1/_0716_ ;
 wire \hash/CA1/_0717_ ;
 wire \hash/CA1/_0718_ ;
 wire \hash/CA1/_0719_ ;
 wire \hash/CA1/_0720_ ;
 wire \hash/CA1/_0721_ ;
 wire \hash/CA1/_0722_ ;
 wire \hash/CA1/_0723_ ;
 wire \hash/CA1/_0724_ ;
 wire \hash/CA1/_0725_ ;
 wire \hash/CA1/_0726_ ;
 wire \hash/CA1/_0727_ ;
 wire \hash/CA1/_0728_ ;
 wire \hash/CA1/_0729_ ;
 wire \hash/CA1/_0730_ ;
 wire \hash/CA1/_0731_ ;
 wire \hash/CA1/_0732_ ;
 wire \hash/CA1/_0733_ ;
 wire \hash/CA1/_0734_ ;
 wire \hash/CA1/_0735_ ;
 wire \hash/CA1/_0736_ ;
 wire \hash/CA1/_0737_ ;
 wire \hash/CA1/_0738_ ;
 wire \hash/CA1/_0739_ ;
 wire \hash/CA1/_0740_ ;
 wire \hash/CA1/_0741_ ;
 wire \hash/CA1/_0742_ ;
 wire \hash/CA1/_0743_ ;
 wire \hash/CA1/_0744_ ;
 wire \hash/CA1/_0745_ ;
 wire \hash/CA1/_0746_ ;
 wire \hash/CA1/_0747_ ;
 wire \hash/CA1/_0748_ ;
 wire \hash/CA1/_0749_ ;
 wire \hash/CA1/_0750_ ;
 wire \hash/CA1/_0751_ ;
 wire \hash/CA1/_0752_ ;
 wire \hash/CA1/_0753_ ;
 wire \hash/CA1/_0754_ ;
 wire \hash/CA1/_0755_ ;
 wire \hash/CA1/_0756_ ;
 wire \hash/CA1/_0757_ ;
 wire \hash/CA1/_0758_ ;
 wire \hash/CA1/_0759_ ;
 wire \hash/CA1/_0760_ ;
 wire \hash/CA1/_0761_ ;
 wire \hash/CA1/_0762_ ;
 wire \hash/CA1/_0763_ ;
 wire \hash/CA1/_0764_ ;
 wire \hash/CA1/_0765_ ;
 wire \hash/CA1/_0766_ ;
 wire \hash/CA1/_0767_ ;
 wire \hash/CA1/_0768_ ;
 wire \hash/CA1/_0769_ ;
 wire \hash/CA1/_0770_ ;
 wire \hash/CA1/_0771_ ;
 wire \hash/CA1/_0772_ ;
 wire \hash/CA1/_0773_ ;
 wire \hash/CA1/_0774_ ;
 wire \hash/CA1/_0775_ ;
 wire \hash/CA1/_0776_ ;
 wire \hash/CA1/_0777_ ;
 wire \hash/CA1/_0778_ ;
 wire \hash/CA1/_0779_ ;
 wire \hash/CA1/_0780_ ;
 wire \hash/CA1/_0781_ ;
 wire \hash/CA1/_0782_ ;
 wire \hash/CA1/_0783_ ;
 wire \hash/CA1/_0784_ ;
 wire \hash/CA1/_0785_ ;
 wire \hash/CA1/_0786_ ;
 wire \hash/CA1/_0787_ ;
 wire \hash/CA1/_0788_ ;
 wire \hash/CA1/_0789_ ;
 wire \hash/CA1/_0790_ ;
 wire \hash/CA1/_0792_ ;
 wire \hash/CA1/_0793_ ;
 wire \hash/CA1/_0794_ ;
 wire \hash/CA1/_0795_ ;
 wire \hash/CA1/_0796_ ;
 wire \hash/CA1/_0797_ ;
 wire \hash/CA1/_0798_ ;
 wire \hash/CA1/_0799_ ;
 wire \hash/CA1/_0800_ ;
 wire \hash/CA1/_0801_ ;
 wire \hash/CA1/_0802_ ;
 wire \hash/CA1/_0803_ ;
 wire \hash/CA1/_0804_ ;
 wire \hash/CA1/_0805_ ;
 wire \hash/CA1/_0806_ ;
 wire \hash/CA1/_0807_ ;
 wire \hash/CA1/_0808_ ;
 wire \hash/CA1/_0809_ ;
 wire \hash/CA1/_0810_ ;
 wire \hash/CA1/_0811_ ;
 wire \hash/CA1/_0812_ ;
 wire \hash/CA1/_0813_ ;
 wire \hash/CA1/_0814_ ;
 wire \hash/CA1/_0815_ ;
 wire \hash/CA1/_0816_ ;
 wire \hash/CA1/_0817_ ;
 wire \hash/CA1/_0818_ ;
 wire \hash/CA1/_0819_ ;
 wire \hash/CA1/_0820_ ;
 wire \hash/CA1/_0821_ ;
 wire \hash/CA1/_0822_ ;
 wire \hash/CA1/_0823_ ;
 wire \hash/CA1/_0824_ ;
 wire \hash/CA1/_0825_ ;
 wire \hash/CA1/_0826_ ;
 wire \hash/CA1/_0827_ ;
 wire \hash/CA1/_0828_ ;
 wire \hash/CA1/_0829_ ;
 wire \hash/CA1/_0830_ ;
 wire \hash/CA1/_0831_ ;
 wire \hash/CA1/_0832_ ;
 wire \hash/CA1/_0833_ ;
 wire \hash/CA1/_0834_ ;
 wire \hash/CA1/_0835_ ;
 wire \hash/CA1/_0836_ ;
 wire \hash/CA1/_0837_ ;
 wire \hash/CA1/_0838_ ;
 wire \hash/CA1/_0839_ ;
 wire \hash/CA1/_0840_ ;
 wire \hash/CA1/_0841_ ;
 wire \hash/CA1/_0842_ ;
 wire \hash/CA1/_0843_ ;
 wire \hash/CA1/_0844_ ;
 wire \hash/CA1/_0845_ ;
 wire \hash/CA1/_0846_ ;
 wire \hash/CA1/_0847_ ;
 wire \hash/CA1/_0848_ ;
 wire \hash/CA1/_0849_ ;
 wire \hash/CA1/_0850_ ;
 wire \hash/CA1/_0851_ ;
 wire \hash/CA1/_0852_ ;
 wire \hash/CA1/_0853_ ;
 wire \hash/CA1/_0854_ ;
 wire \hash/CA1/_0855_ ;
 wire \hash/CA1/_0856_ ;
 wire \hash/CA1/_0857_ ;
 wire \hash/CA1/_0858_ ;
 wire \hash/CA1/_0859_ ;
 wire \hash/CA1/_0860_ ;
 wire \hash/CA1/_0861_ ;
 wire \hash/CA1/_0862_ ;
 wire \hash/CA1/_0863_ ;
 wire \hash/CA1/_0864_ ;
 wire \hash/CA1/_0865_ ;
 wire \hash/CA1/_0866_ ;
 wire \hash/CA1/_0867_ ;
 wire \hash/CA1/_0868_ ;
 wire \hash/CA1/_0869_ ;
 wire \hash/CA1/_0870_ ;
 wire \hash/CA1/_0871_ ;
 wire \hash/CA1/_0872_ ;
 wire \hash/CA1/_0873_ ;
 wire \hash/CA1/_0874_ ;
 wire \hash/CA1/_0875_ ;
 wire \hash/CA1/_0876_ ;
 wire \hash/CA1/_0877_ ;
 wire \hash/CA1/_0878_ ;
 wire \hash/CA1/_0879_ ;
 wire \hash/CA1/_0880_ ;
 wire \hash/CA1/_0881_ ;
 wire \hash/CA1/_0882_ ;
 wire \hash/CA1/_0883_ ;
 wire \hash/CA1/_0884_ ;
 wire \hash/CA1/_0885_ ;
 wire \hash/CA1/_0886_ ;
 wire \hash/CA1/_0887_ ;
 wire \hash/CA1/_0888_ ;
 wire \hash/CA1/_0889_ ;
 wire \hash/CA1/_0890_ ;
 wire \hash/CA1/_0891_ ;
 wire \hash/CA1/_0893_ ;
 wire \hash/CA1/_0894_ ;
 wire \hash/CA1/_0895_ ;
 wire \hash/CA1/_0896_ ;
 wire \hash/CA1/_0897_ ;
 wire \hash/CA1/_0898_ ;
 wire \hash/CA1/_0899_ ;
 wire \hash/CA1/_0900_ ;
 wire \hash/CA1/_0901_ ;
 wire \hash/CA1/_0902_ ;
 wire \hash/CA1/_0903_ ;
 wire \hash/CA1/_0904_ ;
 wire \hash/CA1/_0905_ ;
 wire \hash/CA1/_0906_ ;
 wire \hash/CA1/_0907_ ;
 wire \hash/CA1/_0908_ ;
 wire \hash/CA1/_0909_ ;
 wire \hash/CA1/_0910_ ;
 wire \hash/CA1/_0911_ ;
 wire \hash/CA1/_0912_ ;
 wire \hash/CA1/_0913_ ;
 wire \hash/CA1/_0914_ ;
 wire \hash/CA1/_0915_ ;
 wire \hash/CA1/_0916_ ;
 wire \hash/CA1/_0917_ ;
 wire \hash/CA1/_0918_ ;
 wire \hash/CA1/_0919_ ;
 wire \hash/CA1/_0920_ ;
 wire \hash/CA1/_0921_ ;
 wire \hash/CA1/_0922_ ;
 wire \hash/CA1/_0923_ ;
 wire \hash/CA1/_0924_ ;
 wire \hash/CA1/_0925_ ;
 wire \hash/CA1/_0926_ ;
 wire \hash/CA1/_0927_ ;
 wire \hash/CA1/_0928_ ;
 wire \hash/CA1/_0929_ ;
 wire \hash/CA1/_0930_ ;
 wire \hash/CA1/_0931_ ;
 wire \hash/CA1/_0932_ ;
 wire \hash/CA1/_0933_ ;
 wire \hash/CA1/_0934_ ;
 wire \hash/CA1/_0935_ ;
 wire \hash/CA1/_0936_ ;
 wire \hash/CA1/_0937_ ;
 wire \hash/CA1/_0938_ ;
 wire \hash/CA1/_0939_ ;
 wire \hash/CA1/_0940_ ;
 wire \hash/CA1/_0941_ ;
 wire \hash/CA1/_0942_ ;
 wire \hash/CA1/_0943_ ;
 wire \hash/CA1/_0944_ ;
 wire \hash/CA1/_0945_ ;
 wire \hash/CA1/_0946_ ;
 wire \hash/CA1/_0947_ ;
 wire \hash/CA1/_0948_ ;
 wire \hash/CA1/_0949_ ;
 wire \hash/CA1/_0950_ ;
 wire \hash/CA1/_0951_ ;
 wire \hash/CA1/_0952_ ;
 wire \hash/CA1/_0953_ ;
 wire \hash/CA1/_0954_ ;
 wire \hash/CA1/_0955_ ;
 wire \hash/CA1/_0956_ ;
 wire \hash/CA1/_0957_ ;
 wire \hash/CA1/_0958_ ;
 wire \hash/CA1/_0959_ ;
 wire \hash/CA1/_0960_ ;
 wire \hash/CA1/_0961_ ;
 wire \hash/CA1/_0962_ ;
 wire \hash/CA1/_0963_ ;
 wire \hash/CA1/_0964_ ;
 wire \hash/CA1/_0965_ ;
 wire \hash/CA1/_0966_ ;
 wire \hash/CA1/_0967_ ;
 wire \hash/CA1/_0968_ ;
 wire \hash/CA1/_0969_ ;
 wire \hash/CA1/_0970_ ;
 wire \hash/CA1/_0971_ ;
 wire \hash/CA1/_0972_ ;
 wire \hash/CA1/_0973_ ;
 wire \hash/CA1/_0974_ ;
 wire \hash/CA1/_0975_ ;
 wire \hash/CA1/_0976_ ;
 wire \hash/CA1/_0977_ ;
 wire \hash/CA1/_0978_ ;
 wire \hash/CA1/_0979_ ;
 wire \hash/CA1/_0980_ ;
 wire \hash/CA1/_0981_ ;
 wire \hash/CA1/_0982_ ;
 wire \hash/CA1/_0983_ ;
 wire \hash/CA1/_0984_ ;
 wire \hash/CA1/_0985_ ;
 wire \hash/CA1/_0986_ ;
 wire \hash/CA1/_0987_ ;
 wire \hash/CA1/_0988_ ;
 wire \hash/CA1/_0989_ ;
 wire \hash/CA1/_0990_ ;
 wire \hash/CA1/_0991_ ;
 wire \hash/CA1/_0992_ ;
 wire \hash/CA1/_0993_ ;
 wire \hash/CA1/_0994_ ;
 wire \hash/CA1/_0995_ ;
 wire \hash/CA1/_0996_ ;
 wire \hash/CA1/_0997_ ;
 wire \hash/CA1/_0998_ ;
 wire \hash/CA1/_0999_ ;
 wire \hash/CA1/_1000_ ;
 wire \hash/CA1/_1001_ ;
 wire \hash/CA1/_1002_ ;
 wire \hash/CA1/_1003_ ;
 wire \hash/CA1/_1004_ ;
 wire \hash/CA1/_1005_ ;
 wire \hash/CA1/_1006_ ;
 wire \hash/CA1/_1007_ ;
 wire \hash/CA1/_1008_ ;
 wire \hash/CA1/_1009_ ;
 wire \hash/CA1/_1010_ ;
 wire \hash/CA1/_1011_ ;
 wire \hash/CA1/_1012_ ;
 wire \hash/CA1/_1013_ ;
 wire \hash/CA1/_1014_ ;
 wire \hash/CA1/_1015_ ;
 wire \hash/CA1/_1016_ ;
 wire \hash/CA1/_1017_ ;
 wire \hash/CA1/_1018_ ;
 wire \hash/CA1/_1019_ ;
 wire \hash/CA1/_1020_ ;
 wire \hash/CA1/_1021_ ;
 wire \hash/CA1/_1022_ ;
 wire \hash/CA1/_1023_ ;
 wire \hash/CA1/_1024_ ;
 wire \hash/CA1/_1025_ ;
 wire \hash/CA1/_1026_ ;
 wire \hash/CA1/_1027_ ;
 wire \hash/CA1/_1028_ ;
 wire \hash/CA1/_1029_ ;
 wire \hash/CA1/_1030_ ;
 wire \hash/CA1/_1031_ ;
 wire \hash/CA1/_1032_ ;
 wire \hash/CA1/_1033_ ;
 wire \hash/CA1/_1034_ ;
 wire \hash/CA1/_1035_ ;
 wire \hash/CA1/_1036_ ;
 wire \hash/CA1/_1037_ ;
 wire \hash/CA1/_1038_ ;
 wire \hash/CA1/_1039_ ;
 wire \hash/CA1/_1040_ ;
 wire \hash/CA1/_1041_ ;
 wire \hash/CA1/_1042_ ;
 wire \hash/CA1/_1043_ ;
 wire \hash/CA1/_1044_ ;
 wire \hash/CA1/_1045_ ;
 wire \hash/CA1/_1046_ ;
 wire \hash/CA1/_1047_ ;
 wire \hash/CA1/_1048_ ;
 wire \hash/CA1/_1049_ ;
 wire \hash/CA1/_1050_ ;
 wire \hash/CA1/_1051_ ;
 wire \hash/CA1/_1052_ ;
 wire \hash/CA1/_1053_ ;
 wire \hash/CA1/_1054_ ;
 wire \hash/CA1/_1055_ ;
 wire \hash/CA1/_1056_ ;
 wire \hash/CA1/_1057_ ;
 wire \hash/CA1/_1058_ ;
 wire \hash/CA1/_1059_ ;
 wire \hash/CA1/_1060_ ;
 wire \hash/CA1/_1061_ ;
 wire \hash/CA1/_1062_ ;
 wire \hash/CA1/_1063_ ;
 wire \hash/CA1/_1064_ ;
 wire \hash/CA1/_1065_ ;
 wire \hash/CA1/_1066_ ;
 wire \hash/CA1/_1067_ ;
 wire \hash/CA1/_1068_ ;
 wire \hash/CA1/_1069_ ;
 wire \hash/CA1/_1070_ ;
 wire \hash/CA1/_1071_ ;
 wire \hash/CA1/_1072_ ;
 wire \hash/CA1/_1073_ ;
 wire \hash/CA1/_1074_ ;
 wire \hash/CA1/_1075_ ;
 wire \hash/CA1/_1076_ ;
 wire \hash/CA1/_1077_ ;
 wire \hash/CA1/_1078_ ;
 wire \hash/CA1/_1079_ ;
 wire \hash/CA1/_1080_ ;
 wire \hash/CA1/_1081_ ;
 wire \hash/CA1/_1082_ ;
 wire \hash/CA1/_1083_ ;
 wire \hash/CA1/_1084_ ;
 wire \hash/CA1/_1085_ ;
 wire \hash/CA1/_1086_ ;
 wire \hash/CA1/_1087_ ;
 wire \hash/CA1/_1088_ ;
 wire \hash/CA1/_1089_ ;
 wire \hash/CA1/_1090_ ;
 wire \hash/CA1/_1091_ ;
 wire \hash/CA1/_1092_ ;
 wire \hash/CA1/_1093_ ;
 wire \hash/CA1/_1094_ ;
 wire \hash/CA1/_1095_ ;
 wire \hash/CA1/_1096_ ;
 wire \hash/CA1/_1097_ ;
 wire \hash/CA1/_1098_ ;
 wire \hash/CA1/_1099_ ;
 wire \hash/CA1/_1100_ ;
 wire \hash/CA1/_1101_ ;
 wire \hash/CA1/_1102_ ;
 wire \hash/CA1/_1103_ ;
 wire \hash/CA1/_1104_ ;
 wire \hash/CA1/_1105_ ;
 wire \hash/CA1/_1106_ ;
 wire \hash/CA1/_1107_ ;
 wire \hash/CA1/_1108_ ;
 wire \hash/CA1/_1109_ ;
 wire \hash/CA1/_1110_ ;
 wire \hash/CA1/_1111_ ;
 wire \hash/CA1/_1112_ ;
 wire \hash/CA1/_1113_ ;
 wire \hash/CA1/_1114_ ;
 wire \hash/CA1/_1115_ ;
 wire \hash/CA1/_1116_ ;
 wire \hash/CA1/_1117_ ;
 wire \hash/CA1/_1118_ ;
 wire \hash/CA1/_1119_ ;
 wire \hash/CA1/_1120_ ;
 wire \hash/CA1/_1121_ ;
 wire \hash/CA1/_1122_ ;
 wire \hash/CA1/_1123_ ;
 wire \hash/CA1/_1124_ ;
 wire \hash/CA1/_1125_ ;
 wire \hash/CA1/_1126_ ;
 wire \hash/CA1/_1127_ ;
 wire \hash/CA1/_1128_ ;
 wire \hash/CA1/_1129_ ;
 wire \hash/CA1/_1130_ ;
 wire \hash/CA1/_1131_ ;
 wire \hash/CA1/_1132_ ;
 wire \hash/CA1/_1133_ ;
 wire \hash/CA1/_1134_ ;
 wire \hash/CA1/_1135_ ;
 wire \hash/CA1/_1136_ ;
 wire \hash/CA1/_1137_ ;
 wire \hash/CA1/_1138_ ;
 wire \hash/CA1/_1139_ ;
 wire \hash/CA1/_1140_ ;
 wire \hash/CA1/_1141_ ;
 wire \hash/CA1/_1142_ ;
 wire \hash/CA1/_1143_ ;
 wire \hash/CA1/_1144_ ;
 wire \hash/CA1/_1145_ ;
 wire \hash/CA1/_1146_ ;
 wire \hash/CA1/_1147_ ;
 wire \hash/CA1/_1148_ ;
 wire \hash/CA1/_1149_ ;
 wire \hash/CA1/_1150_ ;
 wire \hash/CA1/_1151_ ;
 wire \hash/CA1/_1152_ ;
 wire \hash/CA1/_1153_ ;
 wire \hash/CA1/_1154_ ;
 wire \hash/CA1/_1155_ ;
 wire \hash/CA1/_1156_ ;
 wire \hash/CA1/_1157_ ;
 wire \hash/CA1/_1158_ ;
 wire \hash/CA1/_1159_ ;
 wire \hash/CA1/_1160_ ;
 wire \hash/CA1/_1161_ ;
 wire \hash/CA1/_1162_ ;
 wire \hash/CA1/_1163_ ;
 wire \hash/CA1/_1164_ ;
 wire \hash/CA1/_1165_ ;
 wire \hash/CA1/_1166_ ;
 wire \hash/CA1/_1167_ ;
 wire \hash/CA1/_1168_ ;
 wire \hash/CA1/_1169_ ;
 wire \hash/CA1/_1170_ ;
 wire \hash/CA1/_1171_ ;
 wire \hash/CA1/_1172_ ;
 wire \hash/CA1/_1173_ ;
 wire \hash/CA1/_1174_ ;
 wire \hash/CA1/_1175_ ;
 wire \hash/CA1/_1176_ ;
 wire \hash/CA1/_1177_ ;
 wire \hash/CA1/_1178_ ;
 wire \hash/CA1/_1179_ ;
 wire \hash/CA1/_1180_ ;
 wire \hash/CA1/_1181_ ;
 wire \hash/CA1/_1182_ ;
 wire \hash/CA1/_1183_ ;
 wire \hash/CA1/_1184_ ;
 wire \hash/CA1/_1185_ ;
 wire \hash/CA1/_1186_ ;
 wire \hash/CA1/_1187_ ;
 wire \hash/CA1/_1188_ ;
 wire \hash/CA1/_1189_ ;
 wire \hash/CA1/_1190_ ;
 wire \hash/CA1/_1191_ ;
 wire \hash/CA1/_1192_ ;
 wire \hash/CA1/_1193_ ;
 wire \hash/CA1/_1194_ ;
 wire \hash/CA1/_1195_ ;
 wire \hash/CA1/_1196_ ;
 wire \hash/CA1/_1197_ ;
 wire \hash/CA1/_1198_ ;
 wire \hash/CA1/_1199_ ;
 wire \hash/CA1/_1200_ ;
 wire \hash/CA1/_1201_ ;
 wire \hash/CA1/_1202_ ;
 wire \hash/CA1/_1203_ ;
 wire \hash/CA1/_1204_ ;
 wire \hash/CA1/_1205_ ;
 wire \hash/CA1/_1206_ ;
 wire \hash/CA1/_1207_ ;
 wire \hash/CA1/_1208_ ;
 wire \hash/CA1/_1209_ ;
 wire \hash/CA1/_1210_ ;
 wire \hash/CA1/_1211_ ;
 wire \hash/CA1/_1212_ ;
 wire \hash/CA1/_1213_ ;
 wire \hash/CA1/_1214_ ;
 wire \hash/CA1/_1215_ ;
 wire \hash/CA1/_1216_ ;
 wire \hash/CA1/_1217_ ;
 wire \hash/CA1/_1218_ ;
 wire \hash/CA1/_1219_ ;
 wire \hash/CA1/_1220_ ;
 wire \hash/CA1/_1221_ ;
 wire \hash/CA1/_1222_ ;
 wire \hash/CA1/_1223_ ;
 wire \hash/CA1/_1224_ ;
 wire \hash/CA1/_1225_ ;
 wire \hash/CA1/_1226_ ;
 wire \hash/CA1/_1227_ ;
 wire \hash/CA1/_1228_ ;
 wire \hash/CA1/_1229_ ;
 wire \hash/CA1/_1230_ ;
 wire \hash/CA1/_1231_ ;
 wire \hash/CA1/_1232_ ;
 wire \hash/CA1/_1233_ ;
 wire \hash/CA1/_1234_ ;
 wire \hash/CA1/_1235_ ;
 wire \hash/CA1/_1236_ ;
 wire \hash/CA1/_1237_ ;
 wire \hash/CA1/_1238_ ;
 wire \hash/CA1/_1239_ ;
 wire \hash/CA1/_1240_ ;
 wire \hash/CA1/_1241_ ;
 wire \hash/CA1/_1242_ ;
 wire \hash/CA1/_1243_ ;
 wire \hash/CA1/_1244_ ;
 wire \hash/CA1/_1245_ ;
 wire \hash/CA1/_1246_ ;
 wire \hash/CA1/_1247_ ;
 wire \hash/CA1/_1248_ ;
 wire \hash/CA1/_1249_ ;
 wire \hash/CA1/_1250_ ;
 wire \hash/CA1/_1251_ ;
 wire \hash/CA1/_1252_ ;
 wire \hash/CA1/_1253_ ;
 wire \hash/CA1/_1254_ ;
 wire \hash/CA1/_1255_ ;
 wire \hash/CA1/_1256_ ;
 wire \hash/CA1/_1257_ ;
 wire \hash/CA1/_1258_ ;
 wire \hash/CA1/_1259_ ;
 wire \hash/CA1/_1260_ ;
 wire \hash/CA1/_1261_ ;
 wire \hash/CA1/_1262_ ;
 wire \hash/CA1/_1263_ ;
 wire \hash/CA1/_1264_ ;
 wire \hash/CA1/_1265_ ;
 wire \hash/CA1/_1266_ ;
 wire \hash/CA1/_1267_ ;
 wire \hash/CA1/_1268_ ;
 wire \hash/CA1/_1269_ ;
 wire \hash/CA1/_1270_ ;
 wire \hash/CA1/_1271_ ;
 wire \hash/CA1/_1272_ ;
 wire \hash/CA1/_1273_ ;
 wire \hash/CA1/_1274_ ;
 wire \hash/CA1/_1275_ ;
 wire \hash/CA1/_1276_ ;
 wire \hash/CA1/_1277_ ;
 wire \hash/CA1/_1278_ ;
 wire \hash/CA1/_1279_ ;
 wire \hash/CA1/_1280_ ;
 wire \hash/CA1/_1281_ ;
 wire \hash/CA1/_1282_ ;
 wire \hash/CA1/_1283_ ;
 wire \hash/CA1/_1284_ ;
 wire \hash/CA1/_1285_ ;
 wire \hash/CA1/_1286_ ;
 wire \hash/CA1/_1287_ ;
 wire \hash/CA1/_1288_ ;
 wire \hash/CA1/_1289_ ;
 wire \hash/CA1/_1290_ ;
 wire \hash/CA1/_1291_ ;
 wire \hash/CA1/_1292_ ;
 wire \hash/CA1/_1293_ ;
 wire \hash/CA1/_1294_ ;
 wire \hash/CA1/_1295_ ;
 wire \hash/CA1/_1296_ ;
 wire \hash/CA1/_1297_ ;
 wire \hash/CA1/_1298_ ;
 wire \hash/CA1/_1299_ ;
 wire \hash/CA1/_1300_ ;
 wire \hash/CA1/_1301_ ;
 wire \hash/CA1/_1302_ ;
 wire \hash/CA1/_1303_ ;
 wire \hash/CA1/_1304_ ;
 wire \hash/CA1/_1305_ ;
 wire \hash/CA1/_1306_ ;
 wire \hash/CA1/_1307_ ;
 wire \hash/CA1/_1308_ ;
 wire \hash/CA1/_1309_ ;
 wire \hash/CA1/_1310_ ;
 wire \hash/CA1/_1311_ ;
 wire \hash/CA1/_1312_ ;
 wire \hash/CA1/_1313_ ;
 wire \hash/CA1/_1314_ ;
 wire \hash/CA1/_1315_ ;
 wire \hash/CA1/_1316_ ;
 wire \hash/CA1/_1317_ ;
 wire \hash/CA1/_1318_ ;
 wire \hash/CA1/_1319_ ;
 wire \hash/CA1/_1320_ ;
 wire \hash/CA1/_1321_ ;
 wire \hash/CA1/_1322_ ;
 wire \hash/CA1/_1323_ ;
 wire \hash/CA1/_1324_ ;
 wire \hash/CA1/_1325_ ;
 wire \hash/CA1/_1326_ ;
 wire \hash/CA1/_1327_ ;
 wire \hash/CA1/_1328_ ;
 wire \hash/CA1/_1329_ ;
 wire \hash/CA1/_1330_ ;
 wire \hash/CA1/_1331_ ;
 wire \hash/CA1/_1332_ ;
 wire \hash/CA1/_1333_ ;
 wire \hash/CA1/_1334_ ;
 wire \hash/CA1/_1335_ ;
 wire \hash/CA1/_1336_ ;
 wire \hash/CA1/_1337_ ;
 wire \hash/CA1/_1338_ ;
 wire \hash/CA1/_1339_ ;
 wire \hash/CA1/_1340_ ;
 wire \hash/CA1/_1341_ ;
 wire \hash/CA1/_1342_ ;
 wire \hash/CA1/_1343_ ;
 wire \hash/CA1/_1344_ ;
 wire \hash/CA1/_1345_ ;
 wire \hash/CA1/_1346_ ;
 wire \hash/CA1/_1347_ ;
 wire \hash/CA1/_1348_ ;
 wire \hash/CA1/_1349_ ;
 wire \hash/CA1/_1350_ ;
 wire \hash/CA1/_1351_ ;
 wire \hash/CA1/_1352_ ;
 wire \hash/CA1/_1353_ ;
 wire \hash/CA1/_1354_ ;
 wire \hash/CA1/_1355_ ;
 wire \hash/CA1/_1356_ ;
 wire \hash/CA1/_1357_ ;
 wire \hash/CA1/_1358_ ;
 wire \hash/CA1/_1359_ ;
 wire \hash/CA1/_1360_ ;
 wire \hash/CA1/_1361_ ;
 wire \hash/CA1/_1362_ ;
 wire \hash/CA1/_1363_ ;
 wire \hash/CA1/_1364_ ;
 wire \hash/CA1/_1365_ ;
 wire \hash/CA1/_1366_ ;
 wire \hash/CA1/_1367_ ;
 wire \hash/CA1/_1368_ ;
 wire \hash/CA1/_1369_ ;
 wire \hash/CA1/_1370_ ;
 wire \hash/CA1/_1371_ ;
 wire \hash/CA1/_1372_ ;
 wire \hash/CA1/_1373_ ;
 wire \hash/CA1/_1374_ ;
 wire \hash/CA1/_1375_ ;
 wire \hash/CA1/_1376_ ;
 wire \hash/CA1/_1377_ ;
 wire \hash/CA1/_1378_ ;
 wire \hash/CA1/_1379_ ;
 wire \hash/CA1/_1380_ ;
 wire \hash/CA1/_1381_ ;
 wire \hash/CA1/_1382_ ;
 wire \hash/CA1/_1383_ ;
 wire \hash/CA1/_1384_ ;
 wire \hash/CA1/_1385_ ;
 wire \hash/CA1/_1386_ ;
 wire \hash/CA1/_1387_ ;
 wire \hash/CA1/_1388_ ;
 wire \hash/CA1/_1389_ ;
 wire \hash/CA1/_1390_ ;
 wire \hash/CA1/_1391_ ;
 wire \hash/CA1/_1392_ ;
 wire \hash/CA1/_1393_ ;
 wire \hash/CA1/_1394_ ;
 wire \hash/CA1/_1395_ ;
 wire \hash/CA1/_1396_ ;
 wire \hash/CA1/_1397_ ;
 wire \hash/CA1/_1398_ ;
 wire \hash/CA1/_1399_ ;
 wire \hash/CA1/_1400_ ;
 wire \hash/CA1/_1401_ ;
 wire \hash/CA1/_1402_ ;
 wire \hash/CA1/_1403_ ;
 wire \hash/CA1/_1404_ ;
 wire \hash/CA1/_1405_ ;
 wire \hash/CA1/_1406_ ;
 wire \hash/CA1/_1407_ ;
 wire \hash/CA1/_1408_ ;
 wire \hash/CA1/_1409_ ;
 wire \hash/CA1/_1410_ ;
 wire \hash/CA1/_1411_ ;
 wire \hash/CA1/_1412_ ;
 wire \hash/CA1/_1413_ ;
 wire \hash/CA1/_1414_ ;
 wire \hash/CA1/_1415_ ;
 wire \hash/CA1/_1416_ ;
 wire \hash/CA1/_1417_ ;
 wire \hash/CA1/_1418_ ;
 wire \hash/CA1/_1419_ ;
 wire \hash/CA1/_1420_ ;
 wire \hash/CA1/_1421_ ;
 wire \hash/CA1/_1422_ ;
 wire \hash/CA1/_1423_ ;
 wire \hash/CA1/_1424_ ;
 wire \hash/CA1/_1425_ ;
 wire \hash/CA1/_1426_ ;
 wire \hash/CA1/_1427_ ;
 wire \hash/CA1/_1428_ ;
 wire \hash/CA1/_1429_ ;
 wire \hash/CA1/_1430_ ;
 wire \hash/CA1/_1431_ ;
 wire \hash/CA1/_1432_ ;
 wire \hash/CA1/_1433_ ;
 wire \hash/CA1/_1434_ ;
 wire \hash/CA1/_1435_ ;
 wire \hash/CA1/_1436_ ;
 wire \hash/CA1/_1437_ ;
 wire \hash/CA1/_1438_ ;
 wire \hash/CA1/_1439_ ;
 wire \hash/CA1/_1440_ ;
 wire \hash/CA1/_1441_ ;
 wire \hash/CA1/_1442_ ;
 wire \hash/CA1/_1443_ ;
 wire \hash/CA1/_1444_ ;
 wire \hash/CA1/_1445_ ;
 wire \hash/CA1/_1446_ ;
 wire \hash/CA1/_1447_ ;
 wire \hash/CA1/_1448_ ;
 wire \hash/CA1/_1449_ ;
 wire \hash/CA1/_1450_ ;
 wire \hash/CA1/_1451_ ;
 wire \hash/CA1/_1452_ ;
 wire \hash/CA1/_1453_ ;
 wire \hash/CA1/_1454_ ;
 wire \hash/CA1/_1455_ ;
 wire \hash/CA1/_1456_ ;
 wire \hash/CA1/_1457_ ;
 wire \hash/CA1/_1458_ ;
 wire \hash/CA1/_1459_ ;
 wire \hash/CA1/_1460_ ;
 wire \hash/CA1/_1461_ ;
 wire \hash/CA1/_1462_ ;
 wire \hash/CA1/_1463_ ;
 wire \hash/CA1/_1464_ ;
 wire \hash/CA1/_1465_ ;
 wire \hash/CA1/_1466_ ;
 wire \hash/CA1/_1467_ ;
 wire \hash/CA1/_1468_ ;
 wire \hash/CA1/_1469_ ;
 wire \hash/CA1/_1470_ ;
 wire \hash/CA1/_1471_ ;
 wire \hash/CA1/_1472_ ;
 wire \hash/CA1/_1473_ ;
 wire \hash/CA1/_1474_ ;
 wire \hash/CA1/_1475_ ;
 wire \hash/CA1/_1476_ ;
 wire \hash/CA1/_1477_ ;
 wire \hash/CA1/_1478_ ;
 wire \hash/CA1/_1479_ ;
 wire \hash/CA1/_1480_ ;
 wire \hash/CA1/_1481_ ;
 wire \hash/CA1/_1482_ ;
 wire \hash/CA1/_1483_ ;
 wire \hash/CA1/_1484_ ;
 wire \hash/CA1/_1485_ ;
 wire \hash/CA1/_1486_ ;
 wire \hash/CA1/_1487_ ;
 wire \hash/CA1/_1488_ ;
 wire \hash/CA1/_1489_ ;
 wire \hash/CA1/_1490_ ;
 wire \hash/CA1/_1491_ ;
 wire \hash/CA1/_1492_ ;
 wire \hash/CA1/_1493_ ;
 wire \hash/CA1/_1494_ ;
 wire \hash/CA1/_1495_ ;
 wire \hash/CA1/_1496_ ;
 wire \hash/CA1/_1497_ ;
 wire \hash/CA1/_1498_ ;
 wire \hash/CA1/_1499_ ;
 wire \hash/CA1/_1500_ ;
 wire \hash/CA1/_1501_ ;
 wire \hash/CA1/_1502_ ;
 wire \hash/CA1/_1503_ ;
 wire \hash/CA1/_1504_ ;
 wire \hash/CA1/_1505_ ;
 wire \hash/CA1/_1506_ ;
 wire \hash/CA1/_1507_ ;
 wire \hash/CA1/_1508_ ;
 wire \hash/CA1/_1509_ ;
 wire \hash/CA1/_1510_ ;
 wire \hash/CA1/_1511_ ;
 wire \hash/CA1/_1512_ ;
 wire \hash/CA1/_1513_ ;
 wire \hash/CA1/_1514_ ;
 wire \hash/CA1/_1515_ ;
 wire \hash/CA1/_1516_ ;
 wire \hash/CA1/_1517_ ;
 wire \hash/CA1/_1518_ ;
 wire \hash/CA1/_1519_ ;
 wire \hash/CA1/_1520_ ;
 wire \hash/CA1/_1521_ ;
 wire \hash/CA1/_1522_ ;
 wire \hash/CA1/_1523_ ;
 wire \hash/CA1/_1524_ ;
 wire \hash/CA1/_1525_ ;
 wire \hash/CA1/_1526_ ;
 wire \hash/CA1/_1527_ ;
 wire \hash/CA1/_1528_ ;
 wire \hash/CA1/_1529_ ;
 wire \hash/CA1/_1530_ ;
 wire \hash/CA1/_1531_ ;
 wire \hash/CA1/_1532_ ;
 wire \hash/CA1/_1533_ ;
 wire \hash/CA1/_1534_ ;
 wire \hash/CA1/_1535_ ;
 wire \hash/CA1/_1536_ ;
 wire \hash/CA1/_1537_ ;
 wire \hash/CA1/_1538_ ;
 wire \hash/CA1/_1539_ ;
 wire \hash/CA1/_1540_ ;
 wire \hash/CA1/_1541_ ;
 wire \hash/CA1/_1542_ ;
 wire \hash/CA1/_1543_ ;
 wire \hash/CA1/_1544_ ;
 wire \hash/CA1/_1545_ ;
 wire \hash/CA1/_1546_ ;
 wire \hash/CA1/_1547_ ;
 wire \hash/CA1/_1548_ ;
 wire \hash/CA1/_1549_ ;
 wire \hash/CA1/_1550_ ;
 wire \hash/CA1/_1551_ ;
 wire \hash/CA1/_1552_ ;
 wire \hash/CA1/_1553_ ;
 wire \hash/CA1/_1554_ ;
 wire \hash/CA1/_1555_ ;
 wire \hash/CA1/_1556_ ;
 wire \hash/CA1/_1557_ ;
 wire \hash/CA1/_1558_ ;
 wire \hash/CA1/_1559_ ;
 wire \hash/CA1/_1560_ ;
 wire \hash/CA1/_1561_ ;
 wire \hash/CA1/_1562_ ;
 wire \hash/CA1/_1563_ ;
 wire \hash/CA1/_1564_ ;
 wire \hash/CA1/_1565_ ;
 wire \hash/CA1/_1566_ ;
 wire \hash/CA1/_1567_ ;
 wire \hash/CA1/_1568_ ;
 wire \hash/CA1/_1569_ ;
 wire \hash/CA1/_1570_ ;
 wire \hash/CA1/_1571_ ;
 wire \hash/CA1/_1572_ ;
 wire \hash/CA1/_1573_ ;
 wire \hash/CA1/_1574_ ;
 wire \hash/CA1/_1575_ ;
 wire \hash/CA1/_1576_ ;
 wire \hash/CA1/_1577_ ;
 wire \hash/CA1/_1578_ ;
 wire \hash/CA1/_1579_ ;
 wire \hash/CA1/_1580_ ;
 wire \hash/CA1/_1581_ ;
 wire \hash/CA1/_1582_ ;
 wire \hash/CA1/_1583_ ;
 wire \hash/CA1/_1584_ ;
 wire \hash/CA1/_1585_ ;
 wire \hash/CA1/_1586_ ;
 wire \hash/CA1/_1587_ ;
 wire \hash/CA1/_1588_ ;
 wire \hash/CA1/_1589_ ;
 wire \hash/CA1/_1590_ ;
 wire \hash/CA1/_1591_ ;
 wire \hash/CA1/_1592_ ;
 wire \hash/CA1/_1593_ ;
 wire \hash/CA1/_1594_ ;
 wire \hash/CA1/_1595_ ;
 wire \hash/CA1/_1596_ ;
 wire \hash/CA1/_1597_ ;
 wire \hash/CA1/_1598_ ;
 wire \hash/CA1/_1599_ ;
 wire \hash/CA1/_1600_ ;
 wire \hash/CA1/_1601_ ;
 wire \hash/CA1/_1602_ ;
 wire \hash/CA1/_1603_ ;
 wire \hash/CA1/_1604_ ;
 wire \hash/CA1/_1605_ ;
 wire \hash/CA1/_1606_ ;
 wire \hash/CA1/_1607_ ;
 wire \hash/CA1/_1608_ ;
 wire \hash/CA1/_1609_ ;
 wire \hash/CA1/_1610_ ;
 wire \hash/CA1/_1611_ ;
 wire \hash/CA1/_1612_ ;
 wire \hash/CA1/_1613_ ;
 wire \hash/CA1/_1614_ ;
 wire \hash/CA1/_1615_ ;
 wire \hash/CA1/_1616_ ;
 wire \hash/CA1/_1617_ ;
 wire \hash/CA1/_1618_ ;
 wire \hash/CA1/_1619_ ;
 wire \hash/CA1/_1620_ ;
 wire \hash/CA1/_1621_ ;
 wire \hash/CA1/_1622_ ;
 wire \hash/CA1/_1623_ ;
 wire \hash/CA1/_1624_ ;
 wire \hash/CA1/_1625_ ;
 wire \hash/CA1/_1626_ ;
 wire \hash/CA1/_1627_ ;
 wire \hash/CA1/_1628_ ;
 wire \hash/CA1/_1629_ ;
 wire \hash/CA1/_1630_ ;
 wire \hash/CA1/_1631_ ;
 wire \hash/CA1/_1632_ ;
 wire \hash/CA1/_1633_ ;
 wire \hash/CA1/_1634_ ;
 wire \hash/CA1/_1635_ ;
 wire \hash/CA1/_1636_ ;
 wire \hash/CA1/_1637_ ;
 wire \hash/CA1/_1638_ ;
 wire \hash/CA1/_1639_ ;
 wire \hash/CA1/_1640_ ;
 wire \hash/CA1/_1641_ ;
 wire \hash/CA1/_1642_ ;
 wire \hash/CA1/_1643_ ;
 wire \hash/CA1/_1644_ ;
 wire \hash/CA1/_1645_ ;
 wire \hash/CA1/_1646_ ;
 wire \hash/CA1/_1647_ ;
 wire \hash/CA1/_1648_ ;
 wire \hash/CA1/_1649_ ;
 wire \hash/CA1/_1650_ ;
 wire \hash/CA1/_1651_ ;
 wire \hash/CA1/_1652_ ;
 wire \hash/CA1/_1653_ ;
 wire \hash/CA1/_1654_ ;
 wire \hash/CA1/_1655_ ;
 wire \hash/CA1/_1656_ ;
 wire \hash/CA1/_1657_ ;
 wire \hash/CA1/_1658_ ;
 wire \hash/CA1/_1659_ ;
 wire \hash/CA1/_1660_ ;
 wire \hash/CA1/_1661_ ;
 wire \hash/CA1/_1662_ ;
 wire \hash/CA1/_1663_ ;
 wire \hash/CA1/_1664_ ;
 wire \hash/CA1/_1665_ ;
 wire \hash/CA1/_1666_ ;
 wire \hash/CA1/_1667_ ;
 wire \hash/CA1/_1668_ ;
 wire \hash/CA1/_1669_ ;
 wire \hash/CA1/_1670_ ;
 wire \hash/CA1/_1671_ ;
 wire \hash/CA1/_1672_ ;
 wire \hash/CA1/_1673_ ;
 wire \hash/CA1/_1674_ ;
 wire \hash/CA1/_1675_ ;
 wire \hash/CA1/_1676_ ;
 wire \hash/CA1/_1677_ ;
 wire \hash/CA1/_1678_ ;
 wire \hash/CA1/_1679_ ;
 wire \hash/CA1/_1680_ ;
 wire \hash/CA1/_1681_ ;
 wire \hash/CA1/_1682_ ;
 wire \hash/CA1/_1683_ ;
 wire \hash/CA1/_1684_ ;
 wire \hash/CA1/_1685_ ;
 wire \hash/CA1/_1686_ ;
 wire \hash/CA1/_1687_ ;
 wire \hash/CA1/_1688_ ;
 wire \hash/CA1/_1689_ ;
 wire \hash/CA1/_1690_ ;
 wire \hash/CA1/_1691_ ;
 wire \hash/CA1/_1692_ ;
 wire \hash/CA1/_1693_ ;
 wire \hash/CA1/_1694_ ;
 wire \hash/CA1/_1695_ ;
 wire \hash/CA1/_1696_ ;
 wire \hash/CA1/_1697_ ;
 wire \hash/CA1/_1698_ ;
 wire \hash/CA1/_1699_ ;
 wire \hash/CA1/_1700_ ;
 wire \hash/CA1/_1701_ ;
 wire \hash/CA1/_1702_ ;
 wire \hash/CA1/_1703_ ;
 wire \hash/CA1/_1704_ ;
 wire \hash/CA1/_1705_ ;
 wire \hash/CA1/_1706_ ;
 wire \hash/CA1/_1707_ ;
 wire \hash/CA1/_1708_ ;
 wire \hash/CA1/_1709_ ;
 wire \hash/CA1/_1710_ ;
 wire \hash/CA1/_1711_ ;
 wire \hash/CA1/_1712_ ;
 wire \hash/CA1/_1713_ ;
 wire \hash/CA1/_1714_ ;
 wire \hash/CA1/_1715_ ;
 wire \hash/CA1/_1716_ ;
 wire \hash/CA1/_1717_ ;
 wire \hash/CA1/_1718_ ;
 wire \hash/CA1/_1719_ ;
 wire \hash/CA1/_1720_ ;
 wire \hash/CA1/_1721_ ;
 wire \hash/CA1/_1722_ ;
 wire \hash/CA1/_1723_ ;
 wire \hash/CA1/_1724_ ;
 wire \hash/CA1/_1725_ ;
 wire \hash/CA1/_1726_ ;
 wire \hash/CA1/_1727_ ;
 wire \hash/CA1/_1728_ ;
 wire \hash/CA1/_1729_ ;
 wire \hash/CA1/_1730_ ;
 wire \hash/CA1/_1731_ ;
 wire \hash/CA1/_1732_ ;
 wire \hash/CA1/_1733_ ;
 wire \hash/CA1/_1734_ ;
 wire \hash/CA1/_1735_ ;
 wire \hash/CA1/_1736_ ;
 wire \hash/CA1/_1737_ ;
 wire \hash/CA1/_1738_ ;
 wire \hash/CA1/_1739_ ;
 wire \hash/CA1/_1740_ ;
 wire \hash/CA1/_1741_ ;
 wire \hash/CA1/_1742_ ;
 wire \hash/CA1/_1743_ ;
 wire \hash/CA1/_1744_ ;
 wire \hash/CA1/_1745_ ;
 wire \hash/CA1/_1746_ ;
 wire \hash/CA1/_1747_ ;
 wire \hash/CA1/_1748_ ;
 wire \hash/CA1/_1749_ ;
 wire \hash/CA1/_1750_ ;
 wire \hash/CA1/_1751_ ;
 wire \hash/CA1/_1752_ ;
 wire \hash/CA1/_1753_ ;
 wire \hash/CA1/_1754_ ;
 wire \hash/CA1/_1755_ ;
 wire \hash/CA1/_1756_ ;
 wire \hash/CA1/_1757_ ;
 wire \hash/CA1/_1758_ ;
 wire \hash/CA1/_1759_ ;
 wire \hash/CA1/_1760_ ;
 wire \hash/CA1/_1761_ ;
 wire \hash/CA1/_1762_ ;
 wire \hash/CA1/_1763_ ;
 wire \hash/CA1/_1764_ ;
 wire \hash/CA1/_1765_ ;
 wire \hash/CA1/_1766_ ;
 wire \hash/CA1/_1767_ ;
 wire \hash/CA1/_1768_ ;
 wire \hash/CA1/_1769_ ;
 wire \hash/CA1/_1770_ ;
 wire \hash/CA1/_1771_ ;
 wire \hash/CA1/_1772_ ;
 wire \hash/CA1/_1773_ ;
 wire \hash/CA1/_1774_ ;
 wire \hash/CA1/_1775_ ;
 wire \hash/CA1/_1776_ ;
 wire \hash/CA1/_1777_ ;
 wire \hash/CA1/_1778_ ;
 wire \hash/CA1/_1779_ ;
 wire \hash/CA1/_1780_ ;
 wire \hash/CA1/_1781_ ;
 wire \hash/CA1/_1782_ ;
 wire \hash/CA1/_1783_ ;
 wire \hash/CA1/_1784_ ;
 wire \hash/CA1/_1785_ ;
 wire \hash/CA1/_1786_ ;
 wire \hash/CA1/_1787_ ;
 wire \hash/CA1/_1788_ ;
 wire \hash/CA1/_1789_ ;
 wire \hash/CA1/_1790_ ;
 wire \hash/CA1/_1791_ ;
 wire \hash/CA1/_1792_ ;
 wire \hash/CA1/_1793_ ;
 wire \hash/CA1/_1794_ ;
 wire \hash/CA1/_1795_ ;
 wire \hash/CA1/_1796_ ;
 wire \hash/CA1/_1797_ ;
 wire \hash/CA1/_1798_ ;
 wire \hash/CA1/_1799_ ;
 wire \hash/CA1/_1800_ ;
 wire \hash/CA1/_1801_ ;
 wire \hash/CA1/_1802_ ;
 wire \hash/CA1/_1803_ ;
 wire \hash/CA1/_1804_ ;
 wire \hash/CA1/_1805_ ;
 wire \hash/CA1/_1806_ ;
 wire \hash/CA1/_1807_ ;
 wire \hash/CA1/_1808_ ;
 wire \hash/CA1/_1809_ ;
 wire \hash/CA1/_1810_ ;
 wire \hash/CA1/_1811_ ;
 wire \hash/CA1/_1812_ ;
 wire \hash/CA1/_1813_ ;
 wire \hash/CA1/_1814_ ;
 wire \hash/CA1/_1815_ ;
 wire \hash/CA1/_1816_ ;
 wire \hash/CA1/_1817_ ;
 wire \hash/CA1/_1818_ ;
 wire \hash/CA1/_1819_ ;
 wire \hash/CA1/_1820_ ;
 wire \hash/CA1/_1821_ ;
 wire \hash/CA1/_1822_ ;
 wire \hash/CA1/_1823_ ;
 wire \hash/CA1/_1824_ ;
 wire \hash/CA1/_1825_ ;
 wire \hash/CA1/_1826_ ;
 wire \hash/CA1/_1827_ ;
 wire \hash/CA1/_1828_ ;
 wire \hash/CA1/_1829_ ;
 wire \hash/CA1/_1830_ ;
 wire \hash/CA1/_1831_ ;
 wire \hash/CA1/_1832_ ;
 wire \hash/CA1/_1833_ ;
 wire \hash/CA1/_1834_ ;
 wire \hash/CA1/_1835_ ;
 wire \hash/CA1/_1836_ ;
 wire \hash/CA1/_1837_ ;
 wire \hash/CA1/_1838_ ;
 wire \hash/CA1/_1839_ ;
 wire \hash/CA1/_1840_ ;
 wire \hash/CA1/_1841_ ;
 wire \hash/CA1/_1842_ ;
 wire \hash/CA1/_1843_ ;
 wire \hash/CA1/_1844_ ;
 wire \hash/CA1/_1845_ ;
 wire \hash/CA1/_1846_ ;
 wire \hash/CA1/_1847_ ;
 wire \hash/CA1/_1848_ ;
 wire \hash/CA1/_1849_ ;
 wire \hash/CA1/_1850_ ;
 wire \hash/CA1/_1851_ ;
 wire \hash/CA1/_1852_ ;
 wire \hash/CA1/_1853_ ;
 wire \hash/CA1/_1854_ ;
 wire \hash/CA1/_1855_ ;
 wire \hash/CA1/_1856_ ;
 wire \hash/CA1/_1857_ ;
 wire \hash/CA1/_1858_ ;
 wire \hash/CA1/_1859_ ;
 wire \hash/CA1/_1860_ ;
 wire \hash/CA1/_1861_ ;
 wire \hash/CA1/_1862_ ;
 wire \hash/CA1/_1863_ ;
 wire \hash/CA1/_1864_ ;
 wire \hash/CA1/_1865_ ;
 wire \hash/CA1/_1866_ ;
 wire \hash/CA1/_1867_ ;
 wire \hash/CA1/_1868_ ;
 wire \hash/CA1/_1869_ ;
 wire \hash/CA1/_1870_ ;
 wire \hash/CA1/_1871_ ;
 wire \hash/CA1/_1872_ ;
 wire \hash/CA1/_1873_ ;
 wire \hash/CA1/_1874_ ;
 wire \hash/CA1/_1875_ ;
 wire \hash/CA1/_1876_ ;
 wire \hash/CA1/_1877_ ;
 wire \hash/CA1/_1878_ ;
 wire \hash/CA1/_1879_ ;
 wire \hash/CA1/_1880_ ;
 wire \hash/CA1/_1881_ ;
 wire \hash/CA1/_1882_ ;
 wire \hash/CA1/_1883_ ;
 wire \hash/CA1/_1884_ ;
 wire \hash/CA1/_1885_ ;
 wire \hash/CA1/_1886_ ;
 wire \hash/CA1/_1887_ ;
 wire \hash/CA1/_1888_ ;
 wire \hash/CA1/_1889_ ;
 wire \hash/CA1/_1890_ ;
 wire \hash/CA1/_1891_ ;
 wire \hash/CA1/_1892_ ;
 wire \hash/CA1/_1893_ ;
 wire \hash/CA1/_1894_ ;
 wire \hash/CA1/_1895_ ;
 wire \hash/CA1/_1896_ ;
 wire \hash/CA1/_1897_ ;
 wire \hash/CA1/_1898_ ;
 wire \hash/CA1/_1899_ ;
 wire \hash/CA1/_1900_ ;
 wire \hash/CA1/_1901_ ;
 wire \hash/CA1/_1902_ ;
 wire \hash/CA1/_1903_ ;
 wire \hash/CA1/_1904_ ;
 wire \hash/CA1/_1905_ ;
 wire \hash/CA1/_1906_ ;
 wire \hash/CA1/_1907_ ;
 wire \hash/CA1/_1908_ ;
 wire \hash/CA1/_1909_ ;
 wire \hash/CA1/_1910_ ;
 wire \hash/CA1/_1911_ ;
 wire \hash/CA1/_1912_ ;
 wire \hash/CA1/_1913_ ;
 wire \hash/CA1/_1914_ ;
 wire \hash/CA1/_1915_ ;
 wire \hash/CA1/_1916_ ;
 wire \hash/CA1/_1917_ ;
 wire \hash/CA1/_1918_ ;
 wire \hash/CA1/_1919_ ;
 wire \hash/CA1/_1920_ ;
 wire \hash/CA1/_1921_ ;
 wire \hash/CA1/_1922_ ;
 wire \hash/CA1/_1923_ ;
 wire \hash/CA1/_1924_ ;
 wire \hash/CA1/_1925_ ;
 wire \hash/CA1/_1926_ ;
 wire \hash/CA1/_1927_ ;
 wire \hash/CA1/_1928_ ;
 wire \hash/CA1/_1929_ ;
 wire \hash/CA1/_1930_ ;
 wire \hash/CA1/_1931_ ;
 wire \hash/CA1/_1932_ ;
 wire \hash/CA1/_1933_ ;
 wire \hash/CA1/_1934_ ;
 wire \hash/CA1/_1935_ ;
 wire \hash/CA1/_1936_ ;
 wire \hash/CA1/_1937_ ;
 wire \hash/CA1/_1938_ ;
 wire \hash/CA1/_1939_ ;
 wire \hash/CA1/_1940_ ;
 wire \hash/CA1/_1941_ ;
 wire \hash/CA1/_1942_ ;
 wire \hash/CA1/_1943_ ;
 wire \hash/CA1/_1944_ ;
 wire \hash/CA1/_1945_ ;
 wire \hash/CA1/_1946_ ;
 wire \hash/CA1/_1947_ ;
 wire \hash/CA1/_1948_ ;
 wire \hash/CA1/_1949_ ;
 wire \hash/CA1/_1950_ ;
 wire \hash/CA1/_1951_ ;
 wire \hash/CA1/_1952_ ;
 wire \hash/CA1/_1953_ ;
 wire \hash/CA1/_1954_ ;
 wire \hash/CA1/_1955_ ;
 wire \hash/CA1/_1956_ ;
 wire \hash/CA1/_1957_ ;
 wire \hash/CA1/_1958_ ;
 wire \hash/CA1/_1959_ ;
 wire \hash/CA1/_1960_ ;
 wire \hash/CA1/_1961_ ;
 wire \hash/CA1/_1962_ ;
 wire \hash/CA1/_1963_ ;
 wire \hash/CA1/_1964_ ;
 wire \hash/CA1/_1965_ ;
 wire \hash/CA1/_1966_ ;
 wire \hash/CA1/_1967_ ;
 wire \hash/CA1/_1968_ ;
 wire \hash/CA1/_1969_ ;
 wire \hash/CA1/_1970_ ;
 wire \hash/CA1/_1971_ ;
 wire \hash/CA1/_1972_ ;
 wire \hash/CA1/_1973_ ;
 wire \hash/CA1/_1974_ ;
 wire \hash/CA1/_1975_ ;
 wire \hash/CA1/_1976_ ;
 wire \hash/CA1/s0[0] ;
 wire \hash/CA1/s0[10] ;
 wire \hash/CA1/s0[11] ;
 wire \hash/CA1/s0[12] ;
 wire \hash/CA1/s0[13] ;
 wire \hash/CA1/s0[14] ;
 wire \hash/CA1/s0[15] ;
 wire \hash/CA1/s0[16] ;
 wire \hash/CA1/s0[17] ;
 wire \hash/CA1/s0[18] ;
 wire \hash/CA1/s0[19] ;
 wire \hash/CA1/s0[1] ;
 wire \hash/CA1/s0[20] ;
 wire \hash/CA1/s0[21] ;
 wire \hash/CA1/s0[22] ;
 wire \hash/CA1/s0[23] ;
 wire \hash/CA1/s0[24] ;
 wire \hash/CA1/s0[25] ;
 wire \hash/CA1/s0[26] ;
 wire \hash/CA1/s0[27] ;
 wire \hash/CA1/s0[28] ;
 wire \hash/CA1/s0[29] ;
 wire \hash/CA1/s0[2] ;
 wire \hash/CA1/s0[30] ;
 wire \hash/CA1/s0[31] ;
 wire \hash/CA1/s0[3] ;
 wire \hash/CA1/s0[4] ;
 wire \hash/CA1/s0[5] ;
 wire \hash/CA1/s0[6] ;
 wire \hash/CA1/s0[7] ;
 wire \hash/CA1/s0[8] ;
 wire \hash/CA1/s0[9] ;
 wire \hash/CA1/s1[0] ;
 wire \hash/CA1/s1[10] ;
 wire \hash/CA1/s1[11] ;
 wire \hash/CA1/s1[12] ;
 wire \hash/CA1/s1[13] ;
 wire \hash/CA1/s1[14] ;
 wire \hash/CA1/s1[15] ;
 wire \hash/CA1/s1[16] ;
 wire \hash/CA1/s1[17] ;
 wire \hash/CA1/s1[18] ;
 wire \hash/CA1/s1[19] ;
 wire \hash/CA1/s1[1] ;
 wire \hash/CA1/s1[20] ;
 wire \hash/CA1/s1[21] ;
 wire \hash/CA1/s1[22] ;
 wire \hash/CA1/s1[23] ;
 wire \hash/CA1/s1[24] ;
 wire \hash/CA1/s1[25] ;
 wire \hash/CA1/s1[26] ;
 wire \hash/CA1/s1[27] ;
 wire \hash/CA1/s1[28] ;
 wire \hash/CA1/s1[29] ;
 wire \hash/CA1/s1[2] ;
 wire \hash/CA1/s1[30] ;
 wire \hash/CA1/s1[31] ;
 wire \hash/CA1/s1[3] ;
 wire \hash/CA1/s1[4] ;
 wire \hash/CA1/s1[5] ;
 wire \hash/CA1/s1[6] ;
 wire \hash/CA1/s1[7] ;
 wire \hash/CA1/s1[8] ;
 wire \hash/CA1/s1[9] ;
 wire \hash/CA2/_0000_ ;
 wire \hash/CA2/_0001_ ;
 wire \hash/CA2/_0002_ ;
 wire \hash/CA2/_0003_ ;
 wire \hash/CA2/_0004_ ;
 wire \hash/CA2/_0005_ ;
 wire \hash/CA2/_0006_ ;
 wire \hash/CA2/_0007_ ;
 wire \hash/CA2/_0008_ ;
 wire \hash/CA2/_0009_ ;
 wire \hash/CA2/_0010_ ;
 wire \hash/CA2/_0011_ ;
 wire \hash/CA2/_0012_ ;
 wire \hash/CA2/_0013_ ;
 wire \hash/CA2/_0014_ ;
 wire \hash/CA2/_0015_ ;
 wire \hash/CA2/_0016_ ;
 wire \hash/CA2/_0017_ ;
 wire \hash/CA2/_0018_ ;
 wire \hash/CA2/_0019_ ;
 wire \hash/CA2/_0020_ ;
 wire \hash/CA2/_0021_ ;
 wire \hash/CA2/_0022_ ;
 wire \hash/CA2/_0023_ ;
 wire \hash/CA2/_0024_ ;
 wire \hash/CA2/_0025_ ;
 wire \hash/CA2/_0026_ ;
 wire \hash/CA2/_0027_ ;
 wire \hash/CA2/_0028_ ;
 wire \hash/CA2/_0029_ ;
 wire \hash/CA2/_0030_ ;
 wire \hash/CA2/_0031_ ;
 wire \hash/CA2/_0032_ ;
 wire \hash/CA2/_0033_ ;
 wire \hash/CA2/_0034_ ;
 wire \hash/CA2/_0035_ ;
 wire \hash/CA2/_0036_ ;
 wire \hash/CA2/_0037_ ;
 wire \hash/CA2/_0038_ ;
 wire \hash/CA2/_0039_ ;
 wire \hash/CA2/_0040_ ;
 wire \hash/CA2/_0041_ ;
 wire \hash/CA2/_0042_ ;
 wire \hash/CA2/_0043_ ;
 wire \hash/CA2/_0044_ ;
 wire \hash/CA2/_0045_ ;
 wire \hash/CA2/_0046_ ;
 wire \hash/CA2/_0047_ ;
 wire \hash/CA2/_0048_ ;
 wire \hash/CA2/_0049_ ;
 wire \hash/CA2/_0050_ ;
 wire \hash/CA2/_0051_ ;
 wire \hash/CA2/_0052_ ;
 wire \hash/CA2/_0053_ ;
 wire \hash/CA2/_0054_ ;
 wire \hash/CA2/_0055_ ;
 wire \hash/CA2/_0056_ ;
 wire \hash/CA2/_0057_ ;
 wire \hash/CA2/_0058_ ;
 wire \hash/CA2/_0059_ ;
 wire \hash/CA2/_0060_ ;
 wire \hash/CA2/_0061_ ;
 wire \hash/CA2/_0062_ ;
 wire \hash/CA2/_0063_ ;
 wire \hash/CA2/_0064_ ;
 wire \hash/CA2/_0065_ ;
 wire \hash/CA2/_0066_ ;
 wire \hash/CA2/_0067_ ;
 wire \hash/CA2/_0068_ ;
 wire \hash/CA2/_0069_ ;
 wire \hash/CA2/_0070_ ;
 wire \hash/CA2/_0071_ ;
 wire \hash/CA2/_0072_ ;
 wire \hash/CA2/_0073_ ;
 wire \hash/CA2/_0074_ ;
 wire \hash/CA2/_0075_ ;
 wire \hash/CA2/_0076_ ;
 wire \hash/CA2/_0077_ ;
 wire \hash/CA2/_0078_ ;
 wire \hash/CA2/_0079_ ;
 wire \hash/CA2/_0080_ ;
 wire \hash/CA2/_0081_ ;
 wire \hash/CA2/_0082_ ;
 wire \hash/CA2/_0083_ ;
 wire \hash/CA2/_0084_ ;
 wire \hash/CA2/_0085_ ;
 wire \hash/CA2/_0086_ ;
 wire \hash/CA2/_0087_ ;
 wire \hash/CA2/_0088_ ;
 wire \hash/CA2/_0089_ ;
 wire \hash/CA2/_0090_ ;
 wire \hash/CA2/_0091_ ;
 wire \hash/CA2/_0092_ ;
 wire \hash/CA2/_0093_ ;
 wire \hash/CA2/_0094_ ;
 wire \hash/CA2/_0095_ ;
 wire \hash/CA2/_0096_ ;
 wire \hash/CA2/_0097_ ;
 wire \hash/CA2/_0098_ ;
 wire \hash/CA2/_0099_ ;
 wire \hash/CA2/_0100_ ;
 wire \hash/CA2/_0101_ ;
 wire \hash/CA2/_0102_ ;
 wire \hash/CA2/_0103_ ;
 wire \hash/CA2/_0104_ ;
 wire \hash/CA2/_0105_ ;
 wire \hash/CA2/_0106_ ;
 wire \hash/CA2/_0107_ ;
 wire \hash/CA2/_0108_ ;
 wire \hash/CA2/_0109_ ;
 wire \hash/CA2/_0110_ ;
 wire \hash/CA2/_0111_ ;
 wire \hash/CA2/_0112_ ;
 wire \hash/CA2/_0113_ ;
 wire \hash/CA2/_0114_ ;
 wire \hash/CA2/_0115_ ;
 wire \hash/CA2/_0116_ ;
 wire \hash/CA2/_0117_ ;
 wire \hash/CA2/_0118_ ;
 wire \hash/CA2/_0119_ ;
 wire \hash/CA2/_0120_ ;
 wire \hash/CA2/_0122_ ;
 wire \hash/CA2/_0123_ ;
 wire \hash/CA2/_0124_ ;
 wire \hash/CA2/_0125_ ;
 wire \hash/CA2/_0126_ ;
 wire \hash/CA2/_0127_ ;
 wire \hash/CA2/_0128_ ;
 wire \hash/CA2/_0129_ ;
 wire \hash/CA2/_0131_ ;
 wire \hash/CA2/_0132_ ;
 wire \hash/CA2/_0133_ ;
 wire \hash/CA2/_0134_ ;
 wire \hash/CA2/_0135_ ;
 wire \hash/CA2/_0136_ ;
 wire \hash/CA2/_0137_ ;
 wire \hash/CA2/_0138_ ;
 wire \hash/CA2/_0139_ ;
 wire \hash/CA2/_0140_ ;
 wire \hash/CA2/_0141_ ;
 wire \hash/CA2/_0142_ ;
 wire \hash/CA2/_0143_ ;
 wire \hash/CA2/_0144_ ;
 wire \hash/CA2/_0145_ ;
 wire \hash/CA2/_0146_ ;
 wire \hash/CA2/_0147_ ;
 wire \hash/CA2/_0148_ ;
 wire \hash/CA2/_0149_ ;
 wire \hash/CA2/_0150_ ;
 wire \hash/CA2/_0151_ ;
 wire \hash/CA2/_0153_ ;
 wire \hash/CA2/_0154_ ;
 wire \hash/CA2/_0155_ ;
 wire \hash/CA2/_0156_ ;
 wire \hash/CA2/_0157_ ;
 wire \hash/CA2/_0158_ ;
 wire \hash/CA2/_0159_ ;
 wire \hash/CA2/_0160_ ;
 wire \hash/CA2/_0161_ ;
 wire \hash/CA2/_0162_ ;
 wire \hash/CA2/_0163_ ;
 wire \hash/CA2/_0164_ ;
 wire \hash/CA2/_0165_ ;
 wire \hash/CA2/_0166_ ;
 wire \hash/CA2/_0167_ ;
 wire \hash/CA2/_0168_ ;
 wire \hash/CA2/_0169_ ;
 wire \hash/CA2/_0170_ ;
 wire \hash/CA2/_0171_ ;
 wire \hash/CA2/_0172_ ;
 wire \hash/CA2/_0173_ ;
 wire \hash/CA2/_0174_ ;
 wire \hash/CA2/_0175_ ;
 wire \hash/CA2/_0176_ ;
 wire \hash/CA2/_0177_ ;
 wire \hash/CA2/_0178_ ;
 wire \hash/CA2/_0179_ ;
 wire \hash/CA2/_0180_ ;
 wire \hash/CA2/_0181_ ;
 wire \hash/CA2/_0182_ ;
 wire \hash/CA2/_0183_ ;
 wire \hash/CA2/_0184_ ;
 wire \hash/CA2/_0185_ ;
 wire \hash/CA2/_0186_ ;
 wire \hash/CA2/_0187_ ;
 wire \hash/CA2/_0188_ ;
 wire \hash/CA2/_0189_ ;
 wire \hash/CA2/_0190_ ;
 wire \hash/CA2/_0191_ ;
 wire \hash/CA2/_0192_ ;
 wire \hash/CA2/_0193_ ;
 wire \hash/CA2/_0194_ ;
 wire \hash/CA2/_0195_ ;
 wire \hash/CA2/_0196_ ;
 wire \hash/CA2/_0197_ ;
 wire \hash/CA2/_0198_ ;
 wire \hash/CA2/_0199_ ;
 wire \hash/CA2/_0200_ ;
 wire \hash/CA2/_0201_ ;
 wire \hash/CA2/_0202_ ;
 wire \hash/CA2/_0203_ ;
 wire \hash/CA2/_0204_ ;
 wire \hash/CA2/_0205_ ;
 wire \hash/CA2/_0206_ ;
 wire \hash/CA2/_0207_ ;
 wire \hash/CA2/_0208_ ;
 wire \hash/CA2/_0209_ ;
 wire \hash/CA2/_0210_ ;
 wire \hash/CA2/_0211_ ;
 wire \hash/CA2/_0212_ ;
 wire \hash/CA2/_0213_ ;
 wire \hash/CA2/_0214_ ;
 wire \hash/CA2/_0215_ ;
 wire \hash/CA2/_0216_ ;
 wire \hash/CA2/_0217_ ;
 wire \hash/CA2/_0218_ ;
 wire \hash/CA2/_0219_ ;
 wire \hash/CA2/_0220_ ;
 wire \hash/CA2/_0221_ ;
 wire \hash/CA2/_0222_ ;
 wire \hash/CA2/_0223_ ;
 wire \hash/CA2/_0224_ ;
 wire \hash/CA2/_0225_ ;
 wire \hash/CA2/_0226_ ;
 wire \hash/CA2/_0227_ ;
 wire \hash/CA2/_0228_ ;
 wire \hash/CA2/_0229_ ;
 wire \hash/CA2/_0230_ ;
 wire \hash/CA2/_0231_ ;
 wire \hash/CA2/_0232_ ;
 wire \hash/CA2/_0233_ ;
 wire \hash/CA2/_0234_ ;
 wire \hash/CA2/_0235_ ;
 wire \hash/CA2/_0236_ ;
 wire \hash/CA2/_0237_ ;
 wire \hash/CA2/_0238_ ;
 wire \hash/CA2/_0239_ ;
 wire \hash/CA2/_0240_ ;
 wire \hash/CA2/_0241_ ;
 wire \hash/CA2/_0242_ ;
 wire \hash/CA2/_0243_ ;
 wire \hash/CA2/_0244_ ;
 wire \hash/CA2/_0245_ ;
 wire \hash/CA2/_0246_ ;
 wire \hash/CA2/_0247_ ;
 wire \hash/CA2/_0248_ ;
 wire \hash/CA2/_0249_ ;
 wire \hash/CA2/_0250_ ;
 wire \hash/CA2/_0251_ ;
 wire \hash/CA2/_0252_ ;
 wire \hash/CA2/_0253_ ;
 wire \hash/CA2/_0254_ ;
 wire \hash/CA2/_0255_ ;
 wire \hash/CA2/_0256_ ;
 wire \hash/CA2/_0257_ ;
 wire \hash/CA2/_0258_ ;
 wire \hash/CA2/_0259_ ;
 wire \hash/CA2/_0260_ ;
 wire \hash/CA2/_0261_ ;
 wire \hash/CA2/_0262_ ;
 wire \hash/CA2/_0263_ ;
 wire \hash/CA2/_0264_ ;
 wire \hash/CA2/_0265_ ;
 wire \hash/CA2/_0266_ ;
 wire \hash/CA2/_0267_ ;
 wire \hash/CA2/_0268_ ;
 wire \hash/CA2/_0269_ ;
 wire \hash/CA2/_0270_ ;
 wire \hash/CA2/_0271_ ;
 wire \hash/CA2/_0272_ ;
 wire \hash/CA2/_0273_ ;
 wire \hash/CA2/_0274_ ;
 wire \hash/CA2/_0275_ ;
 wire \hash/CA2/_0276_ ;
 wire \hash/CA2/_0277_ ;
 wire \hash/CA2/_0278_ ;
 wire \hash/CA2/_0279_ ;
 wire \hash/CA2/_0280_ ;
 wire \hash/CA2/_0281_ ;
 wire \hash/CA2/_0282_ ;
 wire \hash/CA2/_0283_ ;
 wire \hash/CA2/_0284_ ;
 wire \hash/CA2/_0285_ ;
 wire \hash/CA2/_0286_ ;
 wire \hash/CA2/_0287_ ;
 wire \hash/CA2/_0288_ ;
 wire \hash/CA2/_0289_ ;
 wire \hash/CA2/_0290_ ;
 wire \hash/CA2/_0291_ ;
 wire \hash/CA2/_0292_ ;
 wire \hash/CA2/_0293_ ;
 wire \hash/CA2/_0294_ ;
 wire \hash/CA2/_0295_ ;
 wire \hash/CA2/_0296_ ;
 wire \hash/CA2/_0297_ ;
 wire \hash/CA2/_0298_ ;
 wire \hash/CA2/_0299_ ;
 wire \hash/CA2/_0300_ ;
 wire \hash/CA2/_0301_ ;
 wire \hash/CA2/_0302_ ;
 wire \hash/CA2/_0303_ ;
 wire \hash/CA2/_0304_ ;
 wire \hash/CA2/_0305_ ;
 wire \hash/CA2/_0306_ ;
 wire \hash/CA2/_0307_ ;
 wire \hash/CA2/_0308_ ;
 wire \hash/CA2/_0309_ ;
 wire \hash/CA2/_0310_ ;
 wire \hash/CA2/_0311_ ;
 wire \hash/CA2/_0312_ ;
 wire \hash/CA2/_0313_ ;
 wire \hash/CA2/_0314_ ;
 wire \hash/CA2/_0315_ ;
 wire \hash/CA2/_0316_ ;
 wire \hash/CA2/_0317_ ;
 wire \hash/CA2/_0318_ ;
 wire \hash/CA2/_0319_ ;
 wire \hash/CA2/_0320_ ;
 wire \hash/CA2/_0321_ ;
 wire \hash/CA2/_0322_ ;
 wire \hash/CA2/_0323_ ;
 wire \hash/CA2/_0324_ ;
 wire \hash/CA2/_0325_ ;
 wire \hash/CA2/_0326_ ;
 wire \hash/CA2/_0327_ ;
 wire \hash/CA2/_0328_ ;
 wire \hash/CA2/_0329_ ;
 wire \hash/CA2/_0330_ ;
 wire \hash/CA2/_0331_ ;
 wire \hash/CA2/_0332_ ;
 wire \hash/CA2/_0333_ ;
 wire \hash/CA2/_0334_ ;
 wire \hash/CA2/_0335_ ;
 wire \hash/CA2/_0336_ ;
 wire \hash/CA2/_0337_ ;
 wire \hash/CA2/_0338_ ;
 wire \hash/CA2/_0339_ ;
 wire \hash/CA2/_0340_ ;
 wire \hash/CA2/_0341_ ;
 wire \hash/CA2/_0342_ ;
 wire \hash/CA2/_0343_ ;
 wire \hash/CA2/_0344_ ;
 wire \hash/CA2/_0345_ ;
 wire \hash/CA2/_0346_ ;
 wire \hash/CA2/_0347_ ;
 wire \hash/CA2/_0348_ ;
 wire \hash/CA2/_0349_ ;
 wire \hash/CA2/_0350_ ;
 wire \hash/CA2/_0351_ ;
 wire \hash/CA2/_0352_ ;
 wire \hash/CA2/_0353_ ;
 wire \hash/CA2/_0354_ ;
 wire \hash/CA2/_0355_ ;
 wire \hash/CA2/_0356_ ;
 wire \hash/CA2/_0357_ ;
 wire \hash/CA2/_0358_ ;
 wire \hash/CA2/_0359_ ;
 wire \hash/CA2/_0360_ ;
 wire \hash/CA2/_0361_ ;
 wire \hash/CA2/_0362_ ;
 wire \hash/CA2/_0363_ ;
 wire \hash/CA2/_0364_ ;
 wire \hash/CA2/_0365_ ;
 wire \hash/CA2/_0366_ ;
 wire \hash/CA2/_0367_ ;
 wire \hash/CA2/_0368_ ;
 wire \hash/CA2/_0369_ ;
 wire \hash/CA2/_0370_ ;
 wire \hash/CA2/_0371_ ;
 wire \hash/CA2/_0372_ ;
 wire \hash/CA2/_0373_ ;
 wire \hash/CA2/_0374_ ;
 wire \hash/CA2/_0375_ ;
 wire \hash/CA2/_0376_ ;
 wire \hash/CA2/_0377_ ;
 wire \hash/CA2/_0378_ ;
 wire \hash/CA2/_0379_ ;
 wire \hash/CA2/_0380_ ;
 wire \hash/CA2/_0381_ ;
 wire \hash/CA2/_0382_ ;
 wire \hash/CA2/_0383_ ;
 wire \hash/CA2/_0384_ ;
 wire \hash/CA2/_0385_ ;
 wire \hash/CA2/_0386_ ;
 wire \hash/CA2/_0387_ ;
 wire \hash/CA2/_0388_ ;
 wire \hash/CA2/_0389_ ;
 wire \hash/CA2/_0390_ ;
 wire \hash/CA2/_0391_ ;
 wire \hash/CA2/_0392_ ;
 wire \hash/CA2/_0393_ ;
 wire \hash/CA2/_0394_ ;
 wire \hash/CA2/_0395_ ;
 wire \hash/CA2/_0396_ ;
 wire \hash/CA2/_0397_ ;
 wire \hash/CA2/_0398_ ;
 wire \hash/CA2/_0399_ ;
 wire \hash/CA2/_0400_ ;
 wire \hash/CA2/_0401_ ;
 wire \hash/CA2/_0402_ ;
 wire \hash/CA2/_0403_ ;
 wire \hash/CA2/_0404_ ;
 wire \hash/CA2/_0405_ ;
 wire \hash/CA2/_0406_ ;
 wire \hash/CA2/_0407_ ;
 wire \hash/CA2/_0408_ ;
 wire \hash/CA2/_0409_ ;
 wire \hash/CA2/_0410_ ;
 wire \hash/CA2/_0411_ ;
 wire \hash/CA2/_0412_ ;
 wire \hash/CA2/_0413_ ;
 wire \hash/CA2/_0414_ ;
 wire \hash/CA2/_0415_ ;
 wire \hash/CA2/_0416_ ;
 wire \hash/CA2/_0417_ ;
 wire \hash/CA2/_0418_ ;
 wire \hash/CA2/_0419_ ;
 wire \hash/CA2/_0420_ ;
 wire \hash/CA2/_0421_ ;
 wire \hash/CA2/_0422_ ;
 wire \hash/CA2/_0423_ ;
 wire \hash/CA2/_0424_ ;
 wire \hash/CA2/_0425_ ;
 wire \hash/CA2/_0426_ ;
 wire \hash/CA2/_0427_ ;
 wire \hash/CA2/_0428_ ;
 wire \hash/CA2/_0429_ ;
 wire \hash/CA2/_0430_ ;
 wire \hash/CA2/_0431_ ;
 wire \hash/CA2/_0432_ ;
 wire \hash/CA2/_0433_ ;
 wire \hash/CA2/_0434_ ;
 wire \hash/CA2/_0435_ ;
 wire \hash/CA2/_0436_ ;
 wire \hash/CA2/_0437_ ;
 wire \hash/CA2/_0438_ ;
 wire \hash/CA2/_0439_ ;
 wire \hash/CA2/_0440_ ;
 wire \hash/CA2/_0441_ ;
 wire \hash/CA2/_0442_ ;
 wire \hash/CA2/_0443_ ;
 wire \hash/CA2/_0444_ ;
 wire \hash/CA2/_0445_ ;
 wire \hash/CA2/_0446_ ;
 wire \hash/CA2/_0447_ ;
 wire \hash/CA2/_0448_ ;
 wire \hash/CA2/_0449_ ;
 wire \hash/CA2/_0450_ ;
 wire \hash/CA2/_0451_ ;
 wire \hash/CA2/_0452_ ;
 wire \hash/CA2/_0453_ ;
 wire \hash/CA2/_0454_ ;
 wire \hash/CA2/_0455_ ;
 wire \hash/CA2/_0456_ ;
 wire \hash/CA2/_0457_ ;
 wire \hash/CA2/_0458_ ;
 wire \hash/CA2/_0459_ ;
 wire \hash/CA2/_0460_ ;
 wire \hash/CA2/_0461_ ;
 wire \hash/CA2/_0462_ ;
 wire \hash/CA2/_0463_ ;
 wire \hash/CA2/_0464_ ;
 wire \hash/CA2/_0465_ ;
 wire \hash/CA2/_0466_ ;
 wire \hash/CA2/_0467_ ;
 wire \hash/CA2/_0468_ ;
 wire \hash/CA2/_0469_ ;
 wire \hash/CA2/_0470_ ;
 wire \hash/CA2/_0471_ ;
 wire \hash/CA2/_0472_ ;
 wire \hash/CA2/_0473_ ;
 wire \hash/CA2/_0474_ ;
 wire \hash/CA2/_0475_ ;
 wire \hash/CA2/_0476_ ;
 wire \hash/CA2/_0477_ ;
 wire \hash/CA2/_0478_ ;
 wire \hash/CA2/_0479_ ;
 wire \hash/CA2/_0480_ ;
 wire \hash/CA2/_0481_ ;
 wire \hash/CA2/_0482_ ;
 wire \hash/CA2/_0483_ ;
 wire \hash/CA2/_0484_ ;
 wire \hash/CA2/_0485_ ;
 wire \hash/CA2/_0487_ ;
 wire \hash/CA2/_0488_ ;
 wire \hash/CA2/_0489_ ;
 wire \hash/CA2/_0490_ ;
 wire \hash/CA2/_0491_ ;
 wire \hash/CA2/_0492_ ;
 wire \hash/CA2/_0493_ ;
 wire \hash/CA2/_0494_ ;
 wire \hash/CA2/_0495_ ;
 wire \hash/CA2/_0496_ ;
 wire \hash/CA2/_0497_ ;
 wire \hash/CA2/_0498_ ;
 wire \hash/CA2/_0499_ ;
 wire \hash/CA2/_0500_ ;
 wire \hash/CA2/_0501_ ;
 wire \hash/CA2/_0502_ ;
 wire \hash/CA2/_0503_ ;
 wire \hash/CA2/_0504_ ;
 wire \hash/CA2/_0505_ ;
 wire \hash/CA2/_0506_ ;
 wire \hash/CA2/_0507_ ;
 wire \hash/CA2/_0508_ ;
 wire \hash/CA2/_0509_ ;
 wire \hash/CA2/_0510_ ;
 wire \hash/CA2/_0511_ ;
 wire \hash/CA2/_0512_ ;
 wire \hash/CA2/_0513_ ;
 wire \hash/CA2/_0514_ ;
 wire \hash/CA2/_0515_ ;
 wire \hash/CA2/_0516_ ;
 wire \hash/CA2/_0517_ ;
 wire \hash/CA2/_0518_ ;
 wire \hash/CA2/_0519_ ;
 wire \hash/CA2/_0520_ ;
 wire \hash/CA2/_0521_ ;
 wire \hash/CA2/_0522_ ;
 wire \hash/CA2/_0523_ ;
 wire \hash/CA2/_0524_ ;
 wire \hash/CA2/_0525_ ;
 wire \hash/CA2/_0526_ ;
 wire \hash/CA2/_0527_ ;
 wire \hash/CA2/_0528_ ;
 wire \hash/CA2/_0529_ ;
 wire \hash/CA2/_0530_ ;
 wire \hash/CA2/_0531_ ;
 wire \hash/CA2/_0532_ ;
 wire \hash/CA2/_0533_ ;
 wire \hash/CA2/_0534_ ;
 wire \hash/CA2/_0535_ ;
 wire \hash/CA2/_0536_ ;
 wire \hash/CA2/_0537_ ;
 wire \hash/CA2/_0538_ ;
 wire \hash/CA2/_0539_ ;
 wire \hash/CA2/_0540_ ;
 wire \hash/CA2/_0541_ ;
 wire \hash/CA2/_0542_ ;
 wire \hash/CA2/_0543_ ;
 wire \hash/CA2/_0544_ ;
 wire \hash/CA2/_0545_ ;
 wire \hash/CA2/_0546_ ;
 wire \hash/CA2/_0547_ ;
 wire \hash/CA2/_0548_ ;
 wire \hash/CA2/_0549_ ;
 wire \hash/CA2/_0550_ ;
 wire \hash/CA2/_0551_ ;
 wire \hash/CA2/_0552_ ;
 wire \hash/CA2/_0553_ ;
 wire \hash/CA2/_0554_ ;
 wire \hash/CA2/_0555_ ;
 wire \hash/CA2/_0556_ ;
 wire \hash/CA2/_0557_ ;
 wire \hash/CA2/_0558_ ;
 wire \hash/CA2/_0559_ ;
 wire \hash/CA2/_0560_ ;
 wire \hash/CA2/_0561_ ;
 wire \hash/CA2/_0562_ ;
 wire \hash/CA2/_0563_ ;
 wire \hash/CA2/_0564_ ;
 wire \hash/CA2/_0565_ ;
 wire \hash/CA2/_0566_ ;
 wire \hash/CA2/_0567_ ;
 wire \hash/CA2/_0568_ ;
 wire \hash/CA2/_0569_ ;
 wire \hash/CA2/_0570_ ;
 wire \hash/CA2/_0571_ ;
 wire \hash/CA2/_0572_ ;
 wire \hash/CA2/_0573_ ;
 wire \hash/CA2/_0574_ ;
 wire \hash/CA2/_0575_ ;
 wire \hash/CA2/_0576_ ;
 wire \hash/CA2/_0577_ ;
 wire \hash/CA2/_0578_ ;
 wire \hash/CA2/_0579_ ;
 wire \hash/CA2/_0580_ ;
 wire \hash/CA2/_0581_ ;
 wire \hash/CA2/_0582_ ;
 wire \hash/CA2/_0583_ ;
 wire \hash/CA2/_0584_ ;
 wire \hash/CA2/_0585_ ;
 wire \hash/CA2/_0586_ ;
 wire \hash/CA2/_0587_ ;
 wire \hash/CA2/_0588_ ;
 wire \hash/CA2/_0589_ ;
 wire \hash/CA2/_0590_ ;
 wire \hash/CA2/_0591_ ;
 wire \hash/CA2/_0592_ ;
 wire \hash/CA2/_0593_ ;
 wire \hash/CA2/_0594_ ;
 wire \hash/CA2/_0595_ ;
 wire \hash/CA2/_0596_ ;
 wire \hash/CA2/_0597_ ;
 wire \hash/CA2/_0598_ ;
 wire \hash/CA2/_0599_ ;
 wire \hash/CA2/_0600_ ;
 wire \hash/CA2/_0601_ ;
 wire \hash/CA2/_0602_ ;
 wire \hash/CA2/_0603_ ;
 wire \hash/CA2/_0604_ ;
 wire \hash/CA2/_0605_ ;
 wire \hash/CA2/_0606_ ;
 wire \hash/CA2/_0607_ ;
 wire \hash/CA2/_0608_ ;
 wire \hash/CA2/_0609_ ;
 wire \hash/CA2/_0610_ ;
 wire \hash/CA2/_0611_ ;
 wire \hash/CA2/_0612_ ;
 wire \hash/CA2/_0613_ ;
 wire \hash/CA2/_0614_ ;
 wire \hash/CA2/_0615_ ;
 wire \hash/CA2/_0616_ ;
 wire \hash/CA2/_0617_ ;
 wire \hash/CA2/_0618_ ;
 wire \hash/CA2/_0619_ ;
 wire \hash/CA2/_0620_ ;
 wire \hash/CA2/_0621_ ;
 wire \hash/CA2/_0622_ ;
 wire \hash/CA2/_0623_ ;
 wire \hash/CA2/_0624_ ;
 wire \hash/CA2/_0625_ ;
 wire \hash/CA2/_0626_ ;
 wire \hash/CA2/_0627_ ;
 wire \hash/CA2/_0628_ ;
 wire \hash/CA2/_0629_ ;
 wire \hash/CA2/_0630_ ;
 wire \hash/CA2/_0631_ ;
 wire \hash/CA2/_0632_ ;
 wire \hash/CA2/_0633_ ;
 wire \hash/CA2/_0634_ ;
 wire \hash/CA2/_0635_ ;
 wire \hash/CA2/_0636_ ;
 wire \hash/CA2/_0637_ ;
 wire \hash/CA2/_0638_ ;
 wire \hash/CA2/_0639_ ;
 wire \hash/CA2/_0640_ ;
 wire \hash/CA2/_0641_ ;
 wire \hash/CA2/_0642_ ;
 wire \hash/CA2/_0643_ ;
 wire \hash/CA2/_0644_ ;
 wire \hash/CA2/_0645_ ;
 wire \hash/CA2/_0646_ ;
 wire \hash/CA2/_0647_ ;
 wire \hash/CA2/_0648_ ;
 wire \hash/CA2/_0649_ ;
 wire \hash/CA2/_0650_ ;
 wire \hash/CA2/_0651_ ;
 wire \hash/CA2/_0652_ ;
 wire \hash/CA2/_0653_ ;
 wire \hash/CA2/_0654_ ;
 wire \hash/CA2/_0655_ ;
 wire \hash/CA2/_0656_ ;
 wire \hash/CA2/_0657_ ;
 wire \hash/CA2/_0658_ ;
 wire \hash/CA2/_0659_ ;
 wire \hash/CA2/_0660_ ;
 wire \hash/CA2/_0661_ ;
 wire \hash/CA2/_0662_ ;
 wire \hash/CA2/_0663_ ;
 wire \hash/CA2/_0664_ ;
 wire \hash/CA2/_0665_ ;
 wire \hash/CA2/_0666_ ;
 wire \hash/CA2/_0667_ ;
 wire \hash/CA2/_0668_ ;
 wire \hash/CA2/_0669_ ;
 wire \hash/CA2/_0670_ ;
 wire \hash/CA2/_0671_ ;
 wire \hash/CA2/_0672_ ;
 wire \hash/CA2/_0673_ ;
 wire \hash/CA2/_0674_ ;
 wire \hash/CA2/_0675_ ;
 wire \hash/CA2/_0676_ ;
 wire \hash/CA2/_0677_ ;
 wire \hash/CA2/_0678_ ;
 wire \hash/CA2/_0679_ ;
 wire \hash/CA2/_0680_ ;
 wire \hash/CA2/_0681_ ;
 wire \hash/CA2/_0682_ ;
 wire \hash/CA2/_0683_ ;
 wire \hash/CA2/_0684_ ;
 wire \hash/CA2/_0685_ ;
 wire \hash/CA2/_0686_ ;
 wire \hash/CA2/_0687_ ;
 wire \hash/CA2/_0688_ ;
 wire \hash/CA2/_0689_ ;
 wire \hash/CA2/_0690_ ;
 wire \hash/CA2/_0691_ ;
 wire \hash/CA2/_0692_ ;
 wire \hash/CA2/_0693_ ;
 wire \hash/CA2/_0694_ ;
 wire \hash/CA2/_0695_ ;
 wire \hash/CA2/_0696_ ;
 wire \hash/CA2/_0697_ ;
 wire \hash/CA2/_0698_ ;
 wire \hash/CA2/_0699_ ;
 wire \hash/CA2/_0700_ ;
 wire \hash/CA2/_0701_ ;
 wire \hash/CA2/_0702_ ;
 wire \hash/CA2/_0703_ ;
 wire \hash/CA2/_0704_ ;
 wire \hash/CA2/_0705_ ;
 wire \hash/CA2/_0706_ ;
 wire \hash/CA2/_0707_ ;
 wire \hash/CA2/_0708_ ;
 wire \hash/CA2/_0709_ ;
 wire \hash/CA2/_0710_ ;
 wire \hash/CA2/_0711_ ;
 wire \hash/CA2/_0712_ ;
 wire \hash/CA2/_0713_ ;
 wire \hash/CA2/_0714_ ;
 wire \hash/CA2/_0715_ ;
 wire \hash/CA2/_0716_ ;
 wire \hash/CA2/_0717_ ;
 wire \hash/CA2/_0718_ ;
 wire \hash/CA2/_0719_ ;
 wire \hash/CA2/_0720_ ;
 wire \hash/CA2/_0721_ ;
 wire \hash/CA2/_0722_ ;
 wire \hash/CA2/_0723_ ;
 wire \hash/CA2/_0724_ ;
 wire \hash/CA2/_0725_ ;
 wire \hash/CA2/_0726_ ;
 wire \hash/CA2/_0727_ ;
 wire \hash/CA2/_0728_ ;
 wire \hash/CA2/_0729_ ;
 wire \hash/CA2/_0730_ ;
 wire \hash/CA2/_0731_ ;
 wire \hash/CA2/_0732_ ;
 wire \hash/CA2/_0733_ ;
 wire \hash/CA2/_0734_ ;
 wire \hash/CA2/_0735_ ;
 wire \hash/CA2/_0736_ ;
 wire \hash/CA2/_0737_ ;
 wire \hash/CA2/_0738_ ;
 wire \hash/CA2/_0739_ ;
 wire \hash/CA2/_0740_ ;
 wire \hash/CA2/_0741_ ;
 wire \hash/CA2/_0742_ ;
 wire \hash/CA2/_0743_ ;
 wire \hash/CA2/_0744_ ;
 wire \hash/CA2/_0745_ ;
 wire \hash/CA2/_0746_ ;
 wire \hash/CA2/_0747_ ;
 wire \hash/CA2/_0748_ ;
 wire \hash/CA2/_0749_ ;
 wire \hash/CA2/_0750_ ;
 wire \hash/CA2/_0751_ ;
 wire \hash/CA2/_0752_ ;
 wire \hash/CA2/_0753_ ;
 wire \hash/CA2/_0754_ ;
 wire \hash/CA2/_0755_ ;
 wire \hash/CA2/_0756_ ;
 wire \hash/CA2/_0757_ ;
 wire \hash/CA2/_0758_ ;
 wire \hash/CA2/_0759_ ;
 wire \hash/CA2/_0760_ ;
 wire \hash/CA2/_0761_ ;
 wire \hash/CA2/_0762_ ;
 wire \hash/CA2/_0763_ ;
 wire \hash/CA2/_0764_ ;
 wire \hash/CA2/_0765_ ;
 wire \hash/CA2/_0766_ ;
 wire \hash/CA2/_0767_ ;
 wire \hash/CA2/_0768_ ;
 wire \hash/CA2/_0769_ ;
 wire \hash/CA2/_0770_ ;
 wire \hash/CA2/_0771_ ;
 wire \hash/CA2/_0772_ ;
 wire \hash/CA2/_0773_ ;
 wire \hash/CA2/_0774_ ;
 wire \hash/CA2/_0775_ ;
 wire \hash/CA2/_0776_ ;
 wire \hash/CA2/_0777_ ;
 wire \hash/CA2/_0778_ ;
 wire \hash/CA2/_0779_ ;
 wire \hash/CA2/_0780_ ;
 wire \hash/CA2/_0781_ ;
 wire \hash/CA2/_0782_ ;
 wire \hash/CA2/_0783_ ;
 wire \hash/CA2/_0784_ ;
 wire \hash/CA2/_0785_ ;
 wire \hash/CA2/_0786_ ;
 wire \hash/CA2/_0787_ ;
 wire \hash/CA2/_0788_ ;
 wire \hash/CA2/_0789_ ;
 wire \hash/CA2/_0790_ ;
 wire \hash/CA2/_0791_ ;
 wire \hash/CA2/_0792_ ;
 wire \hash/CA2/_0793_ ;
 wire \hash/CA2/_0794_ ;
 wire \hash/CA2/_0795_ ;
 wire \hash/CA2/_0796_ ;
 wire \hash/CA2/_0797_ ;
 wire \hash/CA2/_0798_ ;
 wire \hash/CA2/_0799_ ;
 wire \hash/CA2/_0800_ ;
 wire \hash/CA2/_0801_ ;
 wire \hash/CA2/_0802_ ;
 wire \hash/CA2/_0803_ ;
 wire \hash/CA2/_0804_ ;
 wire \hash/CA2/_0805_ ;
 wire \hash/CA2/_0806_ ;
 wire \hash/CA2/_0807_ ;
 wire \hash/CA2/_0808_ ;
 wire \hash/CA2/_0809_ ;
 wire \hash/CA2/_0810_ ;
 wire \hash/CA2/_0811_ ;
 wire \hash/CA2/_0812_ ;
 wire \hash/CA2/_0813_ ;
 wire \hash/CA2/_0814_ ;
 wire \hash/CA2/_0815_ ;
 wire \hash/CA2/_0816_ ;
 wire \hash/CA2/_0817_ ;
 wire \hash/CA2/_0818_ ;
 wire \hash/CA2/_0819_ ;
 wire \hash/CA2/_0820_ ;
 wire \hash/CA2/_0821_ ;
 wire \hash/CA2/_0822_ ;
 wire \hash/CA2/_0823_ ;
 wire \hash/CA2/_0824_ ;
 wire \hash/CA2/_0825_ ;
 wire \hash/CA2/_0826_ ;
 wire \hash/CA2/_0827_ ;
 wire \hash/CA2/_0828_ ;
 wire \hash/CA2/_0829_ ;
 wire \hash/CA2/_0830_ ;
 wire \hash/CA2/_0831_ ;
 wire \hash/CA2/_0832_ ;
 wire \hash/CA2/_0833_ ;
 wire \hash/CA2/_0834_ ;
 wire \hash/CA2/_0835_ ;
 wire \hash/CA2/_0836_ ;
 wire \hash/CA2/_0837_ ;
 wire \hash/CA2/_0838_ ;
 wire \hash/CA2/_0839_ ;
 wire \hash/CA2/_0840_ ;
 wire \hash/CA2/_0841_ ;
 wire \hash/CA2/_0842_ ;
 wire \hash/CA2/_0843_ ;
 wire \hash/CA2/_0844_ ;
 wire \hash/CA2/_0845_ ;
 wire \hash/CA2/_0846_ ;
 wire \hash/CA2/_0847_ ;
 wire \hash/CA2/_0848_ ;
 wire \hash/CA2/_0849_ ;
 wire \hash/CA2/_0850_ ;
 wire \hash/CA2/_0851_ ;
 wire \hash/CA2/_0852_ ;
 wire \hash/CA2/_0853_ ;
 wire \hash/CA2/_0854_ ;
 wire \hash/CA2/_0855_ ;
 wire \hash/CA2/_0856_ ;
 wire \hash/CA2/_0857_ ;
 wire \hash/CA2/_0858_ ;
 wire \hash/CA2/_0859_ ;
 wire \hash/CA2/_0860_ ;
 wire \hash/CA2/_0861_ ;
 wire \hash/CA2/_0862_ ;
 wire \hash/CA2/_0863_ ;
 wire \hash/CA2/_0864_ ;
 wire \hash/CA2/_0865_ ;
 wire \hash/CA2/_0866_ ;
 wire \hash/CA2/_0867_ ;
 wire \hash/CA2/_0868_ ;
 wire \hash/CA2/_0869_ ;
 wire \hash/CA2/_0870_ ;
 wire \hash/CA2/_0871_ ;
 wire \hash/CA2/_0872_ ;
 wire \hash/CA2/_0873_ ;
 wire \hash/CA2/_0874_ ;
 wire \hash/CA2/_0875_ ;
 wire \hash/CA2/_0876_ ;
 wire \hash/CA2/_0877_ ;
 wire \hash/CA2/_0878_ ;
 wire \hash/CA2/_0879_ ;
 wire \hash/CA2/_0880_ ;
 wire \hash/CA2/_0881_ ;
 wire \hash/CA2/_0882_ ;
 wire \hash/CA2/_0883_ ;
 wire \hash/CA2/_0884_ ;
 wire \hash/CA2/_0885_ ;
 wire \hash/CA2/_0886_ ;
 wire \hash/CA2/_0887_ ;
 wire \hash/CA2/_0888_ ;
 wire \hash/CA2/_0889_ ;
 wire \hash/CA2/_0890_ ;
 wire \hash/CA2/_0891_ ;
 wire \hash/CA2/_0892_ ;
 wire \hash/CA2/_0893_ ;
 wire \hash/CA2/_0894_ ;
 wire \hash/CA2/_0895_ ;
 wire \hash/CA2/_0896_ ;
 wire \hash/CA2/_0897_ ;
 wire \hash/CA2/_0898_ ;
 wire \hash/CA2/_0899_ ;
 wire \hash/CA2/_0900_ ;
 wire \hash/CA2/_0901_ ;
 wire \hash/CA2/_0902_ ;
 wire \hash/CA2/_0903_ ;
 wire \hash/CA2/_0904_ ;
 wire \hash/CA2/_0905_ ;
 wire \hash/CA2/_0906_ ;
 wire \hash/CA2/_0907_ ;
 wire \hash/CA2/_0908_ ;
 wire \hash/CA2/_0909_ ;
 wire \hash/CA2/_0910_ ;
 wire \hash/CA2/_0911_ ;
 wire \hash/CA2/_0912_ ;
 wire \hash/CA2/_0913_ ;
 wire \hash/CA2/_0914_ ;
 wire \hash/CA2/_0915_ ;
 wire \hash/CA2/_0916_ ;
 wire \hash/CA2/_0917_ ;
 wire \hash/CA2/_0918_ ;
 wire \hash/CA2/_0919_ ;
 wire \hash/CA2/_0920_ ;
 wire \hash/CA2/_0921_ ;
 wire \hash/CA2/_0922_ ;
 wire \hash/CA2/_0923_ ;
 wire \hash/CA2/_0924_ ;
 wire \hash/CA2/_0925_ ;
 wire \hash/CA2/_0926_ ;
 wire \hash/CA2/_0927_ ;
 wire \hash/CA2/_0928_ ;
 wire \hash/CA2/_0929_ ;
 wire \hash/CA2/_0930_ ;
 wire \hash/CA2/_0931_ ;
 wire \hash/CA2/_0932_ ;
 wire \hash/CA2/_0933_ ;
 wire \hash/CA2/_0934_ ;
 wire \hash/CA2/_0935_ ;
 wire \hash/CA2/_0936_ ;
 wire \hash/CA2/_0937_ ;
 wire \hash/CA2/_0938_ ;
 wire \hash/CA2/_0939_ ;
 wire \hash/CA2/_0940_ ;
 wire \hash/CA2/_0941_ ;
 wire \hash/CA2/_0942_ ;
 wire \hash/CA2/_0943_ ;
 wire \hash/CA2/_0944_ ;
 wire \hash/CA2/_0945_ ;
 wire \hash/CA2/_0946_ ;
 wire \hash/CA2/_0947_ ;
 wire \hash/CA2/_0948_ ;
 wire \hash/CA2/_0949_ ;
 wire \hash/CA2/_0950_ ;
 wire \hash/CA2/_0951_ ;
 wire \hash/CA2/_0952_ ;
 wire \hash/CA2/_0953_ ;
 wire \hash/CA2/_0954_ ;
 wire \hash/CA2/_0955_ ;
 wire \hash/CA2/_0956_ ;
 wire \hash/CA2/_0957_ ;
 wire \hash/CA2/_0958_ ;
 wire \hash/CA2/_0959_ ;
 wire \hash/CA2/_0960_ ;
 wire \hash/CA2/_0961_ ;
 wire \hash/CA2/_0962_ ;
 wire \hash/CA2/_0963_ ;
 wire \hash/CA2/_0964_ ;
 wire \hash/CA2/_0965_ ;
 wire \hash/CA2/_0966_ ;
 wire \hash/CA2/_0967_ ;
 wire \hash/CA2/_0968_ ;
 wire \hash/CA2/_0969_ ;
 wire \hash/CA2/_0970_ ;
 wire \hash/CA2/_0971_ ;
 wire \hash/CA2/_0972_ ;
 wire \hash/CA2/_0973_ ;
 wire \hash/CA2/_0974_ ;
 wire \hash/CA2/_0975_ ;
 wire \hash/CA2/_0976_ ;
 wire \hash/CA2/_0977_ ;
 wire \hash/CA2/_0978_ ;
 wire \hash/CA2/_0979_ ;
 wire \hash/CA2/_0980_ ;
 wire \hash/CA2/_0981_ ;
 wire \hash/CA2/_0982_ ;
 wire \hash/CA2/_0983_ ;
 wire \hash/CA2/_0984_ ;
 wire \hash/CA2/_0985_ ;
 wire \hash/CA2/_0986_ ;
 wire \hash/CA2/_0987_ ;
 wire \hash/CA2/_0988_ ;
 wire \hash/CA2/_0989_ ;
 wire \hash/CA2/_0990_ ;
 wire \hash/CA2/_0991_ ;
 wire \hash/CA2/_0992_ ;
 wire \hash/CA2/_0993_ ;
 wire \hash/CA2/_0994_ ;
 wire \hash/CA2/_0995_ ;
 wire \hash/CA2/_0996_ ;
 wire \hash/CA2/_0997_ ;
 wire \hash/CA2/_0998_ ;
 wire \hash/CA2/_0999_ ;
 wire \hash/CA2/_1000_ ;
 wire \hash/CA2/_1001_ ;
 wire \hash/CA2/_1002_ ;
 wire \hash/CA2/_1003_ ;
 wire \hash/CA2/_1004_ ;
 wire \hash/CA2/_1005_ ;
 wire \hash/CA2/_1006_ ;
 wire \hash/CA2/_1007_ ;
 wire \hash/CA2/_1008_ ;
 wire \hash/CA2/_1009_ ;
 wire \hash/CA2/_1010_ ;
 wire \hash/CA2/_1011_ ;
 wire \hash/CA2/_1012_ ;
 wire \hash/CA2/_1013_ ;
 wire \hash/CA2/_1014_ ;
 wire \hash/CA2/_1015_ ;
 wire \hash/CA2/_1016_ ;
 wire \hash/CA2/_1017_ ;
 wire \hash/CA2/_1018_ ;
 wire \hash/CA2/_1019_ ;
 wire \hash/CA2/_1020_ ;
 wire \hash/CA2/_1021_ ;
 wire \hash/CA2/_1022_ ;
 wire \hash/CA2/_1023_ ;
 wire \hash/CA2/_1024_ ;
 wire \hash/CA2/_1025_ ;
 wire \hash/CA2/_1026_ ;
 wire \hash/CA2/_1027_ ;
 wire \hash/CA2/_1028_ ;
 wire \hash/CA2/_1029_ ;
 wire \hash/CA2/_1030_ ;
 wire \hash/CA2/_1031_ ;
 wire \hash/CA2/_1032_ ;
 wire \hash/CA2/_1033_ ;
 wire \hash/CA2/_1034_ ;
 wire \hash/CA2/_1035_ ;
 wire \hash/CA2/_1036_ ;
 wire \hash/CA2/_1037_ ;
 wire \hash/CA2/_1038_ ;
 wire \hash/CA2/_1039_ ;
 wire \hash/CA2/_1040_ ;
 wire \hash/CA2/_1041_ ;
 wire \hash/CA2/_1042_ ;
 wire \hash/CA2/_1043_ ;
 wire \hash/CA2/_1044_ ;
 wire \hash/CA2/_1045_ ;
 wire \hash/CA2/_1046_ ;
 wire \hash/CA2/_1047_ ;
 wire \hash/CA2/_1048_ ;
 wire \hash/CA2/_1049_ ;
 wire \hash/CA2/_1050_ ;
 wire \hash/CA2/_1051_ ;
 wire \hash/CA2/_1052_ ;
 wire \hash/CA2/_1053_ ;
 wire \hash/CA2/_1054_ ;
 wire \hash/CA2/_1055_ ;
 wire \hash/CA2/_1056_ ;
 wire \hash/CA2/_1057_ ;
 wire \hash/CA2/_1058_ ;
 wire \hash/CA2/_1059_ ;
 wire \hash/CA2/_1060_ ;
 wire \hash/CA2/_1061_ ;
 wire \hash/CA2/_1062_ ;
 wire \hash/CA2/_1063_ ;
 wire \hash/CA2/_1064_ ;
 wire \hash/CA2/_1065_ ;
 wire \hash/CA2/_1066_ ;
 wire \hash/CA2/_1067_ ;
 wire \hash/CA2/_1068_ ;
 wire \hash/CA2/_1069_ ;
 wire \hash/CA2/_1070_ ;
 wire \hash/CA2/_1071_ ;
 wire \hash/CA2/_1072_ ;
 wire \hash/CA2/_1073_ ;
 wire \hash/CA2/_1074_ ;
 wire \hash/CA2/_1075_ ;
 wire \hash/CA2/_1076_ ;
 wire \hash/CA2/_1077_ ;
 wire \hash/CA2/_1078_ ;
 wire \hash/CA2/_1079_ ;
 wire \hash/CA2/_1080_ ;
 wire \hash/CA2/_1081_ ;
 wire \hash/CA2/_1082_ ;
 wire \hash/CA2/_1083_ ;
 wire \hash/CA2/_1084_ ;
 wire \hash/CA2/_1085_ ;
 wire \hash/CA2/_1086_ ;
 wire \hash/CA2/_1087_ ;
 wire \hash/CA2/_1088_ ;
 wire \hash/CA2/_1089_ ;
 wire \hash/CA2/_1090_ ;
 wire \hash/CA2/_1091_ ;
 wire \hash/CA2/_1092_ ;
 wire \hash/CA2/_1093_ ;
 wire \hash/CA2/_1094_ ;
 wire \hash/CA2/_1095_ ;
 wire \hash/CA2/_1096_ ;
 wire \hash/CA2/_1097_ ;
 wire \hash/CA2/_1098_ ;
 wire \hash/CA2/_1099_ ;
 wire \hash/CA2/_1100_ ;
 wire \hash/CA2/_1101_ ;
 wire \hash/CA2/_1102_ ;
 wire \hash/CA2/_1103_ ;
 wire \hash/CA2/_1104_ ;
 wire \hash/CA2/_1105_ ;
 wire \hash/CA2/_1106_ ;
 wire \hash/CA2/_1107_ ;
 wire \hash/CA2/_1108_ ;
 wire \hash/CA2/_1109_ ;
 wire \hash/CA2/_1110_ ;
 wire \hash/CA2/_1111_ ;
 wire \hash/CA2/_1112_ ;
 wire \hash/CA2/_1113_ ;
 wire \hash/CA2/_1114_ ;
 wire \hash/CA2/_1115_ ;
 wire \hash/CA2/_1116_ ;
 wire \hash/CA2/_1117_ ;
 wire \hash/CA2/_1118_ ;
 wire \hash/CA2/_1119_ ;
 wire \hash/CA2/_1120_ ;
 wire \hash/CA2/_1121_ ;
 wire \hash/CA2/_1122_ ;
 wire \hash/CA2/_1123_ ;
 wire \hash/CA2/_1124_ ;
 wire \hash/CA2/_1125_ ;
 wire \hash/CA2/_1126_ ;
 wire \hash/CA2/_1127_ ;
 wire \hash/CA2/_1128_ ;
 wire \hash/CA2/_1129_ ;
 wire \hash/CA2/_1130_ ;
 wire \hash/CA2/_1131_ ;
 wire \hash/CA2/_1132_ ;
 wire \hash/CA2/_1133_ ;
 wire \hash/CA2/_1134_ ;
 wire \hash/CA2/_1135_ ;
 wire \hash/CA2/_1136_ ;
 wire \hash/CA2/_1137_ ;
 wire \hash/CA2/_1138_ ;
 wire \hash/CA2/_1139_ ;
 wire \hash/CA2/_1140_ ;
 wire \hash/CA2/_1141_ ;
 wire \hash/CA2/_1142_ ;
 wire \hash/CA2/_1143_ ;
 wire \hash/CA2/_1144_ ;
 wire \hash/CA2/_1145_ ;
 wire \hash/CA2/_1146_ ;
 wire \hash/CA2/_1147_ ;
 wire \hash/CA2/_1148_ ;
 wire \hash/CA2/_1149_ ;
 wire \hash/CA2/_1150_ ;
 wire \hash/CA2/_1151_ ;
 wire \hash/CA2/_1152_ ;
 wire \hash/CA2/_1153_ ;
 wire \hash/CA2/_1154_ ;
 wire \hash/CA2/_1155_ ;
 wire \hash/CA2/_1156_ ;
 wire \hash/CA2/_1157_ ;
 wire \hash/CA2/_1158_ ;
 wire \hash/CA2/_1159_ ;
 wire \hash/CA2/_1160_ ;
 wire \hash/CA2/_1161_ ;
 wire \hash/CA2/_1162_ ;
 wire \hash/CA2/_1163_ ;
 wire \hash/CA2/_1164_ ;
 wire \hash/CA2/_1165_ ;
 wire \hash/CA2/_1166_ ;
 wire \hash/CA2/_1167_ ;
 wire \hash/CA2/_1168_ ;
 wire \hash/CA2/_1169_ ;
 wire \hash/CA2/_1170_ ;
 wire \hash/CA2/_1171_ ;
 wire \hash/CA2/_1172_ ;
 wire \hash/CA2/_1173_ ;
 wire \hash/CA2/_1174_ ;
 wire \hash/CA2/_1175_ ;
 wire \hash/CA2/_1176_ ;
 wire \hash/CA2/_1177_ ;
 wire \hash/CA2/_1178_ ;
 wire \hash/CA2/_1179_ ;
 wire \hash/CA2/_1180_ ;
 wire \hash/CA2/_1181_ ;
 wire \hash/CA2/_1182_ ;
 wire \hash/CA2/_1183_ ;
 wire \hash/CA2/_1184_ ;
 wire \hash/CA2/_1185_ ;
 wire \hash/CA2/_1186_ ;
 wire \hash/CA2/_1187_ ;
 wire \hash/CA2/_1188_ ;
 wire \hash/CA2/_1189_ ;
 wire \hash/CA2/_1190_ ;
 wire \hash/CA2/_1191_ ;
 wire \hash/CA2/_1192_ ;
 wire \hash/CA2/_1193_ ;
 wire \hash/CA2/_1194_ ;
 wire \hash/CA2/_1195_ ;
 wire \hash/CA2/_1196_ ;
 wire \hash/CA2/_1197_ ;
 wire \hash/CA2/_1198_ ;
 wire \hash/CA2/_1199_ ;
 wire \hash/CA2/_1200_ ;
 wire \hash/CA2/_1201_ ;
 wire \hash/CA2/_1202_ ;
 wire \hash/CA2/_1203_ ;
 wire \hash/CA2/_1204_ ;
 wire \hash/CA2/_1205_ ;
 wire \hash/CA2/_1206_ ;
 wire \hash/CA2/_1207_ ;
 wire \hash/CA2/_1208_ ;
 wire \hash/CA2/_1209_ ;
 wire \hash/CA2/_1210_ ;
 wire \hash/CA2/_1211_ ;
 wire \hash/CA2/_1212_ ;
 wire \hash/CA2/_1213_ ;
 wire \hash/CA2/s0[0] ;
 wire \hash/CA2/s0[10] ;
 wire \hash/CA2/s0[11] ;
 wire \hash/CA2/s0[12] ;
 wire \hash/CA2/s0[13] ;
 wire \hash/CA2/s0[14] ;
 wire \hash/CA2/s0[15] ;
 wire \hash/CA2/s0[16] ;
 wire \hash/CA2/s0[17] ;
 wire \hash/CA2/s0[18] ;
 wire \hash/CA2/s0[19] ;
 wire \hash/CA2/s0[1] ;
 wire \hash/CA2/s0[20] ;
 wire \hash/CA2/s0[21] ;
 wire \hash/CA2/s0[22] ;
 wire \hash/CA2/s0[23] ;
 wire \hash/CA2/s0[24] ;
 wire \hash/CA2/s0[25] ;
 wire \hash/CA2/s0[26] ;
 wire \hash/CA2/s0[27] ;
 wire \hash/CA2/s0[28] ;
 wire \hash/CA2/s0[29] ;
 wire \hash/CA2/s0[2] ;
 wire \hash/CA2/s0[30] ;
 wire \hash/CA2/s0[31] ;
 wire \hash/CA2/s0[3] ;
 wire \hash/CA2/s0[4] ;
 wire \hash/CA2/s0[5] ;
 wire \hash/CA2/s0[6] ;
 wire \hash/CA2/s0[7] ;
 wire \hash/CA2/s0[8] ;
 wire \hash/CA2/s0[9] ;
 wire \hash/CA2/s1[0] ;
 wire \hash/CA2/s1[10] ;
 wire \hash/CA2/s1[11] ;
 wire \hash/CA2/s1[12] ;
 wire \hash/CA2/s1[13] ;
 wire \hash/CA2/s1[14] ;
 wire \hash/CA2/s1[15] ;
 wire \hash/CA2/s1[16] ;
 wire \hash/CA2/s1[17] ;
 wire \hash/CA2/s1[18] ;
 wire \hash/CA2/s1[19] ;
 wire \hash/CA2/s1[1] ;
 wire \hash/CA2/s1[20] ;
 wire \hash/CA2/s1[21] ;
 wire \hash/CA2/s1[22] ;
 wire \hash/CA2/s1[23] ;
 wire \hash/CA2/s1[24] ;
 wire \hash/CA2/s1[25] ;
 wire \hash/CA2/s1[26] ;
 wire \hash/CA2/s1[27] ;
 wire \hash/CA2/s1[28] ;
 wire \hash/CA2/s1[29] ;
 wire \hash/CA2/s1[2] ;
 wire \hash/CA2/s1[30] ;
 wire \hash/CA2/s1[31] ;
 wire \hash/CA2/s1[3] ;
 wire \hash/CA2/s1[4] ;
 wire \hash/CA2/s1[5] ;
 wire \hash/CA2/s1[6] ;
 wire \hash/CA2/s1[7] ;
 wire \hash/CA2/s1[8] ;
 wire \hash/CA2/s1[9] ;

 sky130_fd_sc_hd__nand4_1 _09580_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_09567_),
    .D(\count_2[5] ),
    .Y(_05330_));
 sky130_fd_sc_hd__or2_2 _09581_ (.A(\count_2[6] ),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__inv_1 _09583_ (.A(_05331_),
    .Y(_00128_));
 sky130_fd_sc_hd__inv_2 _09585_ (.A(reset),
    .Y(_05334_));
 sky130_fd_sc_hd__nor3_1 _09590_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _09592_ (.A(_09554_),
    .B(_05338_),
    .Y(_05340_));
 sky130_fd_sc_hd__nand2_1 _09593_ (.A(_05334_),
    .B(_05340_),
    .Y(_00127_));
 sky130_fd_sc_hd__nor3b_1 _09596_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C_N(\count_1[3] ),
    .Y(_05343_));
 sky130_fd_sc_hd__nand2_1 _09598_ (.A(_09557_),
    .B(_05343_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_1 _09599_ (.A(_05334_),
    .B(_05345_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _09601_ (.A(_09555_),
    .B(_05343_),
    .Y(_05347_));
 sky130_fd_sc_hd__nand2_1 _09602_ (.A(_05334_),
    .B(_05347_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _09604_ (.A(_09559_),
    .B(_05343_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _09605_ (.A(_05334_),
    .B(_05349_),
    .Y(_00124_));
 sky130_fd_sc_hd__nor3b_1 _09606_ (.A(\count_1[5] ),
    .B(\count_1[3] ),
    .C_N(\count_1[4] ),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2_1 _09607_ (.A(_09554_),
    .B(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__nand2_1 _09608_ (.A(_05334_),
    .B(_05351_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _09609_ (.A(_09557_),
    .B(_05350_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_1 _09610_ (.A(_05334_),
    .B(_05352_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_1 _09611_ (.A(_09555_),
    .B(_05350_),
    .Y(_05353_));
 sky130_fd_sc_hd__nand2_1 _09612_ (.A(_05334_),
    .B(_05353_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_1 _09613_ (.A(_09559_),
    .B(_05350_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_1 _09614_ (.A(_05334_),
    .B(_05354_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _09615_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .Y(_05355_));
 sky130_fd_sc_hd__nor2_1 _09616_ (.A(\count_1[5] ),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_1 _09617_ (.A(_09554_),
    .B(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__nand2_1 _09618_ (.A(_05334_),
    .B(_05357_),
    .Y(_00119_));
 sky130_fd_sc_hd__nand2_1 _09621_ (.A(_09557_),
    .B(_05356_),
    .Y(_05360_));
 sky130_fd_sc_hd__nand2_1 _09622_ (.A(_05334_),
    .B(_05360_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_1 _09623_ (.A(_09555_),
    .B(_05356_),
    .Y(_05361_));
 sky130_fd_sc_hd__nand2_1 _09624_ (.A(_05334_),
    .B(_05361_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_1 _09625_ (.A(_09557_),
    .B(_05338_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_1 _09626_ (.A(_05334_),
    .B(_05362_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(_09559_),
    .B(_05356_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(_05334_),
    .B(_05363_),
    .Y(_00115_));
 sky130_fd_sc_hd__nor3b_1 _09629_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C_N(\count_1[5] ),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_1 _09630_ (.A(_09554_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__nand2_1 _09631_ (.A(_05334_),
    .B(_05365_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _09632_ (.A(_09557_),
    .B(_05364_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _09633_ (.A(_05334_),
    .B(_05366_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_1 _09634_ (.A(_09555_),
    .B(_05364_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_05334_),
    .B(_05367_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _09636_ (.A(_09559_),
    .B(_05364_),
    .Y(_05368_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_05334_),
    .B(_05368_),
    .Y(_00111_));
 sky130_fd_sc_hd__and3b_1 _09638_ (.A_N(\count_1[4] ),
    .B(\count_1[3] ),
    .C(\count_1[5] ),
    .X(_05369_));
 sky130_fd_sc_hd__nand2_1 _09640_ (.A(_09554_),
    .B(_05369_),
    .Y(_05371_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(_05334_),
    .B(_05371_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_1 _09642_ (.A(_09557_),
    .B(_05369_),
    .Y(_05372_));
 sky130_fd_sc_hd__nand2_1 _09643_ (.A(_05334_),
    .B(_05372_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand2_1 _09645_ (.A(_09555_),
    .B(_05369_),
    .Y(_05374_));
 sky130_fd_sc_hd__nand2_1 _09646_ (.A(_05334_),
    .B(_05374_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_1 _09647_ (.A(_09559_),
    .B(_05369_),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_1 _09648_ (.A(_05334_),
    .B(_05375_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3b_1 _09649_ (.A_N(\count_1[3] ),
    .B(\count_1[4] ),
    .C(\count_1[5] ),
    .X(_05376_));
 sky130_fd_sc_hd__nand2_1 _09651_ (.A(_09554_),
    .B(_05376_),
    .Y(_05378_));
 sky130_fd_sc_hd__nand2_1 _09652_ (.A(_05334_),
    .B(_05378_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_1 _09653_ (.A(_09555_),
    .B(_05338_),
    .Y(_05379_));
 sky130_fd_sc_hd__nand2_1 _09654_ (.A(_05334_),
    .B(_05379_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_1 _09655_ (.A(_09557_),
    .B(_05376_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand2_1 _09656_ (.A(_05334_),
    .B(_05380_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_1 _09657_ (.A(_09555_),
    .B(_05376_),
    .Y(_05381_));
 sky130_fd_sc_hd__nand2_1 _09658_ (.A(_05334_),
    .B(_05381_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_1 _09659_ (.A(_09559_),
    .B(_05376_),
    .Y(_05382_));
 sky130_fd_sc_hd__nand2_1 _09660_ (.A(_05334_),
    .B(_05382_),
    .Y(_00102_));
 sky130_fd_sc_hd__and3_1 _09661_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .X(_05383_));
 sky130_fd_sc_hd__nand2_1 _09663_ (.A(_09554_),
    .B(_05383_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand2_1 _09664_ (.A(_05334_),
    .B(_05385_),
    .Y(_00101_));
 sky130_fd_sc_hd__nor3b_1 _09668_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .C_N(\count_2[3] ),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(_09565_),
    .B(_05389_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _09671_ (.A(_05334_),
    .B(_05391_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_1 _09672_ (.A(_09557_),
    .B(_05383_),
    .Y(_05392_));
 sky130_fd_sc_hd__nand2_1 _09673_ (.A(_05334_),
    .B(_05392_),
    .Y(_00100_));
 sky130_fd_sc_hd__nand2_1 _09676_ (.A(_09563_),
    .B(_05389_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_1 _09677_ (.A(_05334_),
    .B(_05395_),
    .Y(_00094_));
 sky130_fd_sc_hd__nand2_1 _09679_ (.A(_09567_),
    .B(_05389_),
    .Y(_05397_));
 sky130_fd_sc_hd__nand2_1 _09680_ (.A(_05334_),
    .B(_05397_),
    .Y(_00093_));
 sky130_fd_sc_hd__nand2b_1 _09682_ (.A_N(\count_2[3] ),
    .B(\count_2[4] ),
    .Y(_05399_));
 sky130_fd_sc_hd__nor2_1 _09683_ (.A(\count_2[5] ),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_1 _09684_ (.A(_09562_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__nand2_1 _09685_ (.A(_05334_),
    .B(_05401_),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_1 _09686_ (.A(_09565_),
    .B(_05400_),
    .Y(_05402_));
 sky130_fd_sc_hd__nand2_1 _09687_ (.A(_05334_),
    .B(_05402_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor3_1 _09688_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(\count_2[5] ),
    .Y(_05403_));
 sky130_fd_sc_hd__nand2_1 _09690_ (.A(_09562_),
    .B(_05403_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_1 _09691_ (.A(_05334_),
    .B(_05405_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_1 _09692_ (.A(_09563_),
    .B(_05400_),
    .Y(_05406_));
 sky130_fd_sc_hd__nand2_1 _09693_ (.A(_05334_),
    .B(_05406_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_1 _09694_ (.A(_09555_),
    .B(_05383_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_1 _09695_ (.A(_05334_),
    .B(_05407_),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_1 _09696_ (.A(\count_2[5] ),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_1 _09697_ (.A(_09567_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__o21ai_2 _09698_ (.A1(_05399_),
    .A2(_05409_),
    .B1(_05334_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_1 _09699_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .Y(_05410_));
 sky130_fd_sc_hd__nor2_1 _09700_ (.A(\count_2[5] ),
    .B(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_1 _09701_ (.A(_09562_),
    .B(_05411_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _09702_ (.A(_05334_),
    .B(_05412_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand2_1 _09703_ (.A(_09565_),
    .B(_05411_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_05334_),
    .B(_05413_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_1 _09705_ (.A(_09563_),
    .B(_05411_),
    .Y(_05414_));
 sky130_fd_sc_hd__nand2_1 _09706_ (.A(_05334_),
    .B(_05414_),
    .Y(_00085_));
 sky130_fd_sc_hd__nand2_1 _09708_ (.A(_09567_),
    .B(_05411_),
    .Y(_05416_));
 sky130_fd_sc_hd__nand2_1 _09709_ (.A(_05334_),
    .B(_05416_),
    .Y(_00084_));
 sky130_fd_sc_hd__nor3_1 _09710_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_05408_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_1 _09711_ (.A(_09562_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__nand2_1 _09712_ (.A(_05334_),
    .B(_05418_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_1 _09713_ (.A(_09559_),
    .B(_05383_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_1 _09714_ (.A(_05334_),
    .B(_05419_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(_09565_),
    .B(_05417_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand2_1 _09716_ (.A(_05334_),
    .B(_05420_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand2_1 _09717_ (.A(_09563_),
    .B(_05417_),
    .Y(_05421_));
 sky130_fd_sc_hd__nand2_1 _09718_ (.A(_05334_),
    .B(_05421_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _09719_ (.A(_09567_),
    .B(\count_2[5] ),
    .Y(_05422_));
 sky130_fd_sc_hd__o31ai_4 _09720_ (.A1(\count_2[4] ),
    .A2(\count_2[3] ),
    .A3(_05422_),
    .B1(_05334_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_1 _09721_ (.A(_09565_),
    .B(_05403_),
    .Y(_05423_));
 sky130_fd_sc_hd__nand2_1 _09722_ (.A(_05334_),
    .B(_05423_),
    .Y(_00079_));
 sky130_fd_sc_hd__nor3b_1 _09723_ (.A(_05408_),
    .B(\count_2[4] ),
    .C_N(\count_2[3] ),
    .Y(_05424_));
 sky130_fd_sc_hd__nand2_1 _09724_ (.A(_09562_),
    .B(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _09725_ (.A(_05334_),
    .B(_05425_),
    .Y(_00078_));
 sky130_fd_sc_hd__nand2_1 _09726_ (.A(_09565_),
    .B(_05424_),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_1 _09727_ (.A(_05334_),
    .B(_05426_),
    .Y(_00077_));
 sky130_fd_sc_hd__nand2_1 _09728_ (.A(_09559_),
    .B(_05338_),
    .Y(_05427_));
 sky130_fd_sc_hd__nand2_1 _09729_ (.A(_05334_),
    .B(_05427_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_1 _09730_ (.A(_09563_),
    .B(_05424_),
    .Y(_05428_));
 sky130_fd_sc_hd__nand2_1 _09731_ (.A(_05334_),
    .B(_05428_),
    .Y(_00076_));
 sky130_fd_sc_hd__nand2_1 _09733_ (.A(_09567_),
    .B(_05424_),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _09734_ (.A(_05334_),
    .B(_05430_),
    .Y(_00075_));
 sky130_fd_sc_hd__nor2_1 _09735_ (.A(_05408_),
    .B(_05399_),
    .Y(_05431_));
 sky130_fd_sc_hd__nand2_1 _09736_ (.A(_09562_),
    .B(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand2_1 _09737_ (.A(_05334_),
    .B(_05432_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_1 _09738_ (.A(_09565_),
    .B(_05431_),
    .Y(_05433_));
 sky130_fd_sc_hd__nand2_1 _09739_ (.A(_05334_),
    .B(_05433_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_1 _09740_ (.A(_09563_),
    .B(_05431_),
    .Y(_05434_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_05334_),
    .B(_05434_),
    .Y(_00072_));
 sky130_fd_sc_hd__o21ai_2 _09742_ (.A1(_05422_),
    .A2(_05399_),
    .B1(_05334_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand2_1 _09743_ (.A(_09554_),
    .B(_05343_),
    .Y(_05435_));
 sky130_fd_sc_hd__nand2_1 _09744_ (.A(_05334_),
    .B(_05435_),
    .Y(_00096_));
 sky130_fd_sc_hd__nor2_1 _09745_ (.A(_05408_),
    .B(_05410_),
    .Y(_05436_));
 sky130_fd_sc_hd__nand2_1 _09746_ (.A(_09562_),
    .B(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__nand2_1 _09747_ (.A(_05334_),
    .B(_05437_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_1 _09748_ (.A(_09565_),
    .B(_05436_),
    .Y(_05438_));
 sky130_fd_sc_hd__nand2_1 _09749_ (.A(_05334_),
    .B(_05438_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_1 _09750_ (.A(_09563_),
    .B(_05403_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_1 _09751_ (.A(_05334_),
    .B(_05439_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_1 _09752_ (.A(_09563_),
    .B(_05436_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_1 _09753_ (.A(_05334_),
    .B(_05440_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_1 _09754_ (.A(_05334_),
    .B(_05330_),
    .Y(_00066_));
 sky130_fd_sc_hd__o31ai_4 _09755_ (.A1(\count_2[4] ),
    .A2(\count_2[3] ),
    .A3(_05409_),
    .B1(_05334_),
    .Y(_00065_));
 sky130_fd_sc_hd__nand2_1 _09757_ (.A(_09562_),
    .B(_05389_),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_1 _09758_ (.A(_05334_),
    .B(_05442_),
    .Y(_00064_));
 sky130_fd_sc_hd__mux4_2 _09764_ (.A0(\w[19][0] ),
    .A1(\w[23][0] ),
    .A2(\w[17][0] ),
    .A3(\w[21][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05448_));
 sky130_fd_sc_hd__mux4_2 _09767_ (.A0(\w[27][0] ),
    .A1(\w[31][0] ),
    .A2(\w[25][0] ),
    .A3(\w[29][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05451_));
 sky130_fd_sc_hd__mux4_2 _09768_ (.A0(\w[3][0] ),
    .A1(\w[7][0] ),
    .A2(\w[1][0] ),
    .A3(\w[5][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05452_));
 sky130_fd_sc_hd__mux4_2 _09772_ (.A0(\w[11][0] ),
    .A1(\w[15][0] ),
    .A2(\w[9][0] ),
    .A3(\w[13][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05456_));
 sky130_fd_sc_hd__xor2_4 _09774_ (.A(\count_hash2[3] ),
    .B(_09354_),
    .X(_05458_));
 sky130_fd_sc_hd__nand3_1 _09776_ (.A(\count_hash2[3] ),
    .B(\count_hash2[2] ),
    .C(\count_hash2[1] ),
    .Y(_05460_));
 sky130_fd_sc_hd__xor2_4 _09777_ (.A(\count_hash2[4] ),
    .B(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__mux4_2 _09780_ (.A0(_05448_),
    .A1(_05451_),
    .A2(_05452_),
    .A3(_05456_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05464_));
 sky130_fd_sc_hd__mux4_2 _09781_ (.A0(\w[51][0] ),
    .A1(\w[55][0] ),
    .A2(\w[49][0] ),
    .A3(\w[53][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05465_));
 sky130_fd_sc_hd__mux4_2 _09782_ (.A0(\w[59][0] ),
    .A1(\w[63][0] ),
    .A2(\w[57][0] ),
    .A3(\w[61][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05466_));
 sky130_fd_sc_hd__mux4_2 _09783_ (.A0(\w[35][0] ),
    .A1(\w[39][0] ),
    .A2(\w[33][0] ),
    .A3(\w[37][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05467_));
 sky130_fd_sc_hd__mux4_2 _09785_ (.A0(\w[43][0] ),
    .A1(\w[47][0] ),
    .A2(\w[41][0] ),
    .A3(\w[45][0] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05469_));
 sky130_fd_sc_hd__mux4_2 _09786_ (.A0(_05465_),
    .A1(_05466_),
    .A2(_05467_),
    .A3(_05469_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05470_));
 sky130_fd_sc_hd__nand3_1 _09787_ (.A(\count_hash2[4] ),
    .B(\count_hash2[3] ),
    .C(_09354_),
    .Y(_05471_));
 sky130_fd_sc_hd__xnor2_2 _09788_ (.A(\count_hash2[5] ),
    .B(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__mux2i_1 _09791_ (.A0(_05464_),
    .A1(_05470_),
    .S(_05472_),
    .Y(_05475_));
 sky130_fd_sc_hd__inv_1 _09792_ (.A(reset_hash),
    .Y(_05476_));
 sky130_fd_sc_hd__inv_1 _09793_ (.A(\count_hash1[2] ),
    .Y(_09356_));
 sky130_fd_sc_hd__nand3_1 _09796_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(\count_hash1[5] ),
    .Y(_05479_));
 sky130_fd_sc_hd__nor3_1 _09797_ (.A(_09356_),
    .B(_09360_),
    .C(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__nor2_1 _09798_ (.A(\count_hash1[6] ),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(_05476_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand2_1 _09803_ (.A(reset_hash),
    .B(\w[1][0] ),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_0 _09804_ (.A1(_05475_),
    .A2(_05482_),
    .B1(_05486_),
    .Y(_00032_));
 sky130_fd_sc_hd__mux4_2 _09809_ (.A0(\w[19][1] ),
    .A1(\w[23][1] ),
    .A2(\w[17][1] ),
    .A3(\w[21][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05491_));
 sky130_fd_sc_hd__mux4_2 _09812_ (.A0(\w[27][1] ),
    .A1(\w[31][1] ),
    .A2(\w[25][1] ),
    .A3(\w[29][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05494_));
 sky130_fd_sc_hd__mux4_2 _09815_ (.A0(\w[3][1] ),
    .A1(\w[7][1] ),
    .A2(\w[1][1] ),
    .A3(\w[5][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05497_));
 sky130_fd_sc_hd__mux4_2 _09818_ (.A0(\w[11][1] ),
    .A1(\w[15][1] ),
    .A2(\w[9][1] ),
    .A3(\w[13][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05500_));
 sky130_fd_sc_hd__mux4_2 _09822_ (.A0(_05491_),
    .A1(_05494_),
    .A2(_05497_),
    .A3(_05500_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05504_));
 sky130_fd_sc_hd__mux4_2 _09825_ (.A0(\w[51][1] ),
    .A1(\w[55][1] ),
    .A2(\w[49][1] ),
    .A3(\w[53][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05507_));
 sky130_fd_sc_hd__mux4_2 _09826_ (.A0(\w[59][1] ),
    .A1(\w[63][1] ),
    .A2(\w[57][1] ),
    .A3(\w[61][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05508_));
 sky130_fd_sc_hd__mux4_2 _09827_ (.A0(\w[35][1] ),
    .A1(\w[39][1] ),
    .A2(\w[33][1] ),
    .A3(\w[37][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05509_));
 sky130_fd_sc_hd__mux4_2 _09830_ (.A0(\w[43][1] ),
    .A1(\w[47][1] ),
    .A2(\w[41][1] ),
    .A3(\w[45][1] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05512_));
 sky130_fd_sc_hd__mux4_2 _09833_ (.A0(_05507_),
    .A1(_05508_),
    .A2(_05509_),
    .A3(_05512_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05515_));
 sky130_fd_sc_hd__mux2i_1 _09836_ (.A0(_05504_),
    .A1(_05515_),
    .S(_05472_),
    .Y(_05518_));
 sky130_fd_sc_hd__nand2_1 _09837_ (.A(reset_hash),
    .B(\w[1][1] ),
    .Y(_05519_));
 sky130_fd_sc_hd__o21ai_0 _09838_ (.A1(_05482_),
    .A2(_05518_),
    .B1(_05519_),
    .Y(_00043_));
 sky130_fd_sc_hd__mux4_2 _09840_ (.A0(\w[19][2] ),
    .A1(\w[23][2] ),
    .A2(\w[17][2] ),
    .A3(\w[21][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05521_));
 sky130_fd_sc_hd__mux4_2 _09842_ (.A0(\w[27][2] ),
    .A1(\w[31][2] ),
    .A2(\w[25][2] ),
    .A3(\w[29][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05523_));
 sky130_fd_sc_hd__mux4_2 _09843_ (.A0(\w[3][2] ),
    .A1(\w[7][2] ),
    .A2(\w[1][2] ),
    .A3(\w[5][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05524_));
 sky130_fd_sc_hd__mux4_2 _09844_ (.A0(\w[11][2] ),
    .A1(\w[15][2] ),
    .A2(\w[9][2] ),
    .A3(\w[13][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05525_));
 sky130_fd_sc_hd__mux4_2 _09845_ (.A0(_05521_),
    .A1(_05523_),
    .A2(_05524_),
    .A3(_05525_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05526_));
 sky130_fd_sc_hd__mux4_2 _09846_ (.A0(\w[51][2] ),
    .A1(\w[55][2] ),
    .A2(\w[49][2] ),
    .A3(\w[53][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05527_));
 sky130_fd_sc_hd__mux4_2 _09847_ (.A0(\w[59][2] ),
    .A1(\w[63][2] ),
    .A2(\w[57][2] ),
    .A3(\w[61][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05528_));
 sky130_fd_sc_hd__mux4_2 _09848_ (.A0(\w[35][2] ),
    .A1(\w[39][2] ),
    .A2(\w[33][2] ),
    .A3(\w[37][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05529_));
 sky130_fd_sc_hd__mux4_2 _09849_ (.A0(\w[43][2] ),
    .A1(\w[47][2] ),
    .A2(\w[41][2] ),
    .A3(\w[45][2] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05530_));
 sky130_fd_sc_hd__mux4_2 _09851_ (.A0(_05527_),
    .A1(_05528_),
    .A2(_05529_),
    .A3(_05530_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05532_));
 sky130_fd_sc_hd__mux2i_1 _09852_ (.A0(_05526_),
    .A1(_05532_),
    .S(_05472_),
    .Y(_05533_));
 sky130_fd_sc_hd__nand2_1 _09853_ (.A(reset_hash),
    .B(\w[1][2] ),
    .Y(_05534_));
 sky130_fd_sc_hd__o21ai_0 _09854_ (.A1(_05482_),
    .A2(_05533_),
    .B1(_05534_),
    .Y(_00054_));
 sky130_fd_sc_hd__mux4_2 _09855_ (.A0(\w[19][3] ),
    .A1(\w[23][3] ),
    .A2(\w[17][3] ),
    .A3(\w[21][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05535_));
 sky130_fd_sc_hd__mux4_2 _09857_ (.A0(\w[27][3] ),
    .A1(\w[31][3] ),
    .A2(\w[25][3] ),
    .A3(\w[29][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05537_));
 sky130_fd_sc_hd__mux4_2 _09858_ (.A0(\w[3][3] ),
    .A1(\w[7][3] ),
    .A2(\w[1][3] ),
    .A3(\w[5][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05538_));
 sky130_fd_sc_hd__mux4_2 _09859_ (.A0(\w[11][3] ),
    .A1(\w[15][3] ),
    .A2(\w[9][3] ),
    .A3(\w[13][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05539_));
 sky130_fd_sc_hd__mux4_2 _09860_ (.A0(_05535_),
    .A1(_05537_),
    .A2(_05538_),
    .A3(_05539_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05540_));
 sky130_fd_sc_hd__mux4_2 _09861_ (.A0(\w[51][3] ),
    .A1(\w[55][3] ),
    .A2(\w[49][3] ),
    .A3(\w[53][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05541_));
 sky130_fd_sc_hd__mux4_2 _09862_ (.A0(\w[59][3] ),
    .A1(\w[63][3] ),
    .A2(\w[57][3] ),
    .A3(\w[61][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05542_));
 sky130_fd_sc_hd__mux4_2 _09864_ (.A0(\w[35][3] ),
    .A1(\w[39][3] ),
    .A2(\w[33][3] ),
    .A3(\w[37][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05544_));
 sky130_fd_sc_hd__mux4_2 _09865_ (.A0(\w[43][3] ),
    .A1(\w[47][3] ),
    .A2(\w[41][3] ),
    .A3(\w[45][3] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05545_));
 sky130_fd_sc_hd__mux4_2 _09866_ (.A0(_05541_),
    .A1(_05542_),
    .A2(_05544_),
    .A3(_05545_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05546_));
 sky130_fd_sc_hd__mux2i_1 _09867_ (.A0(_05540_),
    .A1(_05546_),
    .S(_05472_),
    .Y(_05547_));
 sky130_fd_sc_hd__nand2_1 _09868_ (.A(reset_hash),
    .B(\w[1][3] ),
    .Y(_05548_));
 sky130_fd_sc_hd__o21ai_0 _09869_ (.A1(_05482_),
    .A2(_05547_),
    .B1(_05548_),
    .Y(_00057_));
 sky130_fd_sc_hd__mux4_2 _09870_ (.A0(\w[19][4] ),
    .A1(\w[23][4] ),
    .A2(\w[17][4] ),
    .A3(\w[21][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05549_));
 sky130_fd_sc_hd__mux4_2 _09871_ (.A0(\w[27][4] ),
    .A1(\w[31][4] ),
    .A2(\w[25][4] ),
    .A3(\w[29][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05550_));
 sky130_fd_sc_hd__mux4_2 _09872_ (.A0(\w[3][4] ),
    .A1(\w[7][4] ),
    .A2(\w[1][4] ),
    .A3(\w[5][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05551_));
 sky130_fd_sc_hd__mux4_2 _09873_ (.A0(\w[11][4] ),
    .A1(\w[15][4] ),
    .A2(\w[9][4] ),
    .A3(\w[13][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05552_));
 sky130_fd_sc_hd__mux4_2 _09875_ (.A0(_05549_),
    .A1(_05550_),
    .A2(_05551_),
    .A3(_05552_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05554_));
 sky130_fd_sc_hd__mux4_2 _09876_ (.A0(\w[51][4] ),
    .A1(\w[55][4] ),
    .A2(\w[49][4] ),
    .A3(\w[53][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05555_));
 sky130_fd_sc_hd__mux4_2 _09877_ (.A0(\w[59][4] ),
    .A1(\w[63][4] ),
    .A2(\w[57][4] ),
    .A3(\w[61][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05556_));
 sky130_fd_sc_hd__mux4_2 _09879_ (.A0(\w[35][4] ),
    .A1(\w[39][4] ),
    .A2(\w[33][4] ),
    .A3(\w[37][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05558_));
 sky130_fd_sc_hd__mux4_2 _09880_ (.A0(\w[43][4] ),
    .A1(\w[47][4] ),
    .A2(\w[41][4] ),
    .A3(\w[45][4] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05559_));
 sky130_fd_sc_hd__mux4_2 _09881_ (.A0(_05555_),
    .A1(_05556_),
    .A2(_05558_),
    .A3(_05559_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05560_));
 sky130_fd_sc_hd__mux2i_1 _09882_ (.A0(_05554_),
    .A1(_05560_),
    .S(_05472_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(reset_hash),
    .B(\w[1][4] ),
    .Y(_05563_));
 sky130_fd_sc_hd__o21ai_0 _09885_ (.A1(_05482_),
    .A2(_05561_),
    .B1(_05563_),
    .Y(_00058_));
 sky130_fd_sc_hd__mux4_2 _09886_ (.A0(\w[19][5] ),
    .A1(\w[23][5] ),
    .A2(\w[17][5] ),
    .A3(\w[21][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05564_));
 sky130_fd_sc_hd__mux4_2 _09887_ (.A0(\w[27][5] ),
    .A1(\w[31][5] ),
    .A2(\w[25][5] ),
    .A3(\w[29][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05565_));
 sky130_fd_sc_hd__mux4_2 _09888_ (.A0(\w[3][5] ),
    .A1(\w[7][5] ),
    .A2(\w[1][5] ),
    .A3(\w[5][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05566_));
 sky130_fd_sc_hd__mux4_2 _09889_ (.A0(\w[11][5] ),
    .A1(\w[15][5] ),
    .A2(\w[9][5] ),
    .A3(\w[13][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05567_));
 sky130_fd_sc_hd__mux4_2 _09890_ (.A0(_05564_),
    .A1(_05565_),
    .A2(_05566_),
    .A3(_05567_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05568_));
 sky130_fd_sc_hd__mux4_2 _09892_ (.A0(\w[51][5] ),
    .A1(\w[55][5] ),
    .A2(\w[49][5] ),
    .A3(\w[53][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05570_));
 sky130_fd_sc_hd__mux4_2 _09893_ (.A0(\w[59][5] ),
    .A1(\w[63][5] ),
    .A2(\w[57][5] ),
    .A3(\w[61][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05571_));
 sky130_fd_sc_hd__mux4_2 _09894_ (.A0(\w[35][5] ),
    .A1(\w[39][5] ),
    .A2(\w[33][5] ),
    .A3(\w[37][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05572_));
 sky130_fd_sc_hd__mux4_2 _09895_ (.A0(\w[43][5] ),
    .A1(\w[47][5] ),
    .A2(\w[41][5] ),
    .A3(\w[45][5] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05573_));
 sky130_fd_sc_hd__mux4_2 _09897_ (.A0(_05570_),
    .A1(_05571_),
    .A2(_05572_),
    .A3(_05573_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05575_));
 sky130_fd_sc_hd__mux2i_1 _09898_ (.A0(_05568_),
    .A1(_05575_),
    .S(_05472_),
    .Y(_05576_));
 sky130_fd_sc_hd__nand2_1 _09899_ (.A(reset_hash),
    .B(\w[1][5] ),
    .Y(_05577_));
 sky130_fd_sc_hd__o21ai_0 _09900_ (.A1(_05482_),
    .A2(_05576_),
    .B1(_05577_),
    .Y(_00059_));
 sky130_fd_sc_hd__mux4_2 _09901_ (.A0(\w[19][6] ),
    .A1(\w[23][6] ),
    .A2(\w[17][6] ),
    .A3(\w[21][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05578_));
 sky130_fd_sc_hd__mux4_2 _09902_ (.A0(\w[27][6] ),
    .A1(\w[31][6] ),
    .A2(\w[25][6] ),
    .A3(\w[29][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05579_));
 sky130_fd_sc_hd__mux4_2 _09904_ (.A0(\w[3][6] ),
    .A1(\w[7][6] ),
    .A2(\w[1][6] ),
    .A3(\w[5][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05581_));
 sky130_fd_sc_hd__mux4_2 _09905_ (.A0(\w[11][6] ),
    .A1(\w[15][6] ),
    .A2(\w[9][6] ),
    .A3(\w[13][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05582_));
 sky130_fd_sc_hd__mux4_2 _09907_ (.A0(_05578_),
    .A1(_05579_),
    .A2(_05581_),
    .A3(_05582_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05584_));
 sky130_fd_sc_hd__mux4_2 _09909_ (.A0(\w[51][6] ),
    .A1(\w[55][6] ),
    .A2(\w[49][6] ),
    .A3(\w[53][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05586_));
 sky130_fd_sc_hd__mux4_2 _09910_ (.A0(\w[59][6] ),
    .A1(\w[63][6] ),
    .A2(\w[57][6] ),
    .A3(\w[61][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05587_));
 sky130_fd_sc_hd__mux4_2 _09911_ (.A0(\w[35][6] ),
    .A1(\w[39][6] ),
    .A2(\w[33][6] ),
    .A3(\w[37][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05588_));
 sky130_fd_sc_hd__mux4_2 _09912_ (.A0(\w[43][6] ),
    .A1(\w[47][6] ),
    .A2(\w[41][6] ),
    .A3(\w[45][6] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05589_));
 sky130_fd_sc_hd__mux4_2 _09913_ (.A0(_05586_),
    .A1(_05587_),
    .A2(_05588_),
    .A3(_05589_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05590_));
 sky130_fd_sc_hd__mux2i_1 _09914_ (.A0(_05584_),
    .A1(_05590_),
    .S(_05472_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand2_1 _09915_ (.A(reset_hash),
    .B(\w[1][6] ),
    .Y(_05592_));
 sky130_fd_sc_hd__o21ai_0 _09916_ (.A1(_05482_),
    .A2(_05591_),
    .B1(_05592_),
    .Y(_00060_));
 sky130_fd_sc_hd__mux4_2 _09918_ (.A0(\w[19][7] ),
    .A1(\w[23][7] ),
    .A2(\w[17][7] ),
    .A3(\w[21][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05594_));
 sky130_fd_sc_hd__mux4_2 _09919_ (.A0(\w[27][7] ),
    .A1(\w[31][7] ),
    .A2(\w[25][7] ),
    .A3(\w[29][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05595_));
 sky130_fd_sc_hd__mux4_2 _09921_ (.A0(\w[3][7] ),
    .A1(\w[7][7] ),
    .A2(\w[1][7] ),
    .A3(\w[5][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05597_));
 sky130_fd_sc_hd__mux4_2 _09922_ (.A0(\w[11][7] ),
    .A1(\w[15][7] ),
    .A2(\w[9][7] ),
    .A3(\w[13][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05598_));
 sky130_fd_sc_hd__mux4_2 _09923_ (.A0(_05594_),
    .A1(_05595_),
    .A2(_05597_),
    .A3(_05598_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05599_));
 sky130_fd_sc_hd__mux4_2 _09924_ (.A0(\w[51][7] ),
    .A1(\w[55][7] ),
    .A2(\w[49][7] ),
    .A3(\w[53][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05600_));
 sky130_fd_sc_hd__mux4_2 _09925_ (.A0(\w[59][7] ),
    .A1(\w[63][7] ),
    .A2(\w[57][7] ),
    .A3(\w[61][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05601_));
 sky130_fd_sc_hd__mux4_2 _09926_ (.A0(\w[35][7] ),
    .A1(\w[39][7] ),
    .A2(\w[33][7] ),
    .A3(\w[37][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05602_));
 sky130_fd_sc_hd__mux4_2 _09927_ (.A0(\w[43][7] ),
    .A1(\w[47][7] ),
    .A2(\w[41][7] ),
    .A3(\w[45][7] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05603_));
 sky130_fd_sc_hd__mux4_2 _09928_ (.A0(_05600_),
    .A1(_05601_),
    .A2(_05602_),
    .A3(_05603_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05604_));
 sky130_fd_sc_hd__mux2i_1 _09929_ (.A0(_05599_),
    .A1(_05604_),
    .S(_05472_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(reset_hash),
    .B(\w[1][7] ),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_0 _09931_ (.A1(_05482_),
    .A2(_05605_),
    .B1(_05606_),
    .Y(_00061_));
 sky130_fd_sc_hd__mux4_2 _09933_ (.A0(\w[19][8] ),
    .A1(\w[23][8] ),
    .A2(\w[17][8] ),
    .A3(\w[21][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05608_));
 sky130_fd_sc_hd__mux4_2 _09934_ (.A0(\w[27][8] ),
    .A1(\w[31][8] ),
    .A2(\w[25][8] ),
    .A3(\w[29][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05609_));
 sky130_fd_sc_hd__mux4_2 _09935_ (.A0(\w[3][8] ),
    .A1(\w[7][8] ),
    .A2(\w[1][8] ),
    .A3(\w[5][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05610_));
 sky130_fd_sc_hd__mux4_2 _09936_ (.A0(\w[11][8] ),
    .A1(\w[15][8] ),
    .A2(\w[9][8] ),
    .A3(\w[13][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05611_));
 sky130_fd_sc_hd__mux4_2 _09937_ (.A0(_05608_),
    .A1(_05609_),
    .A2(_05610_),
    .A3(_05611_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05612_));
 sky130_fd_sc_hd__mux4_2 _09938_ (.A0(\w[51][8] ),
    .A1(\w[55][8] ),
    .A2(\w[49][8] ),
    .A3(\w[53][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05613_));
 sky130_fd_sc_hd__mux4_2 _09939_ (.A0(\w[59][8] ),
    .A1(\w[63][8] ),
    .A2(\w[57][8] ),
    .A3(\w[61][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05614_));
 sky130_fd_sc_hd__mux4_2 _09940_ (.A0(\w[35][8] ),
    .A1(\w[39][8] ),
    .A2(\w[33][8] ),
    .A3(\w[37][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05615_));
 sky130_fd_sc_hd__mux4_2 _09942_ (.A0(\w[43][8] ),
    .A1(\w[47][8] ),
    .A2(\w[41][8] ),
    .A3(\w[45][8] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05617_));
 sky130_fd_sc_hd__mux4_2 _09943_ (.A0(_05613_),
    .A1(_05614_),
    .A2(_05615_),
    .A3(_05617_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05618_));
 sky130_fd_sc_hd__mux2i_1 _09945_ (.A0(_05612_),
    .A1(_05618_),
    .S(_05472_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _09946_ (.A(reset_hash),
    .B(\w[1][8] ),
    .Y(_05621_));
 sky130_fd_sc_hd__o21ai_0 _09947_ (.A1(_05482_),
    .A2(_05620_),
    .B1(_05621_),
    .Y(_00062_));
 sky130_fd_sc_hd__mux4_2 _09948_ (.A0(\w[19][9] ),
    .A1(\w[23][9] ),
    .A2(\w[17][9] ),
    .A3(\w[21][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05622_));
 sky130_fd_sc_hd__mux4_2 _09949_ (.A0(\w[27][9] ),
    .A1(\w[31][9] ),
    .A2(\w[25][9] ),
    .A3(\w[29][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05623_));
 sky130_fd_sc_hd__mux4_2 _09950_ (.A0(\w[3][9] ),
    .A1(\w[7][9] ),
    .A2(\w[1][9] ),
    .A3(\w[5][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05624_));
 sky130_fd_sc_hd__mux4_2 _09952_ (.A0(\w[11][9] ),
    .A1(\w[15][9] ),
    .A2(\w[9][9] ),
    .A3(\w[13][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05626_));
 sky130_fd_sc_hd__mux4_2 _09953_ (.A0(_05622_),
    .A1(_05623_),
    .A2(_05624_),
    .A3(_05626_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05627_));
 sky130_fd_sc_hd__mux4_2 _09954_ (.A0(\w[51][9] ),
    .A1(\w[55][9] ),
    .A2(\w[49][9] ),
    .A3(\w[53][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05628_));
 sky130_fd_sc_hd__mux4_2 _09956_ (.A0(\w[59][9] ),
    .A1(\w[63][9] ),
    .A2(\w[57][9] ),
    .A3(\w[61][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05630_));
 sky130_fd_sc_hd__mux4_2 _09957_ (.A0(\w[35][9] ),
    .A1(\w[39][9] ),
    .A2(\w[33][9] ),
    .A3(\w[37][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05631_));
 sky130_fd_sc_hd__mux4_2 _09959_ (.A0(\w[43][9] ),
    .A1(\w[47][9] ),
    .A2(\w[41][9] ),
    .A3(\w[45][9] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05633_));
 sky130_fd_sc_hd__mux4_2 _09960_ (.A0(_05628_),
    .A1(_05630_),
    .A2(_05631_),
    .A3(_05633_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05634_));
 sky130_fd_sc_hd__mux2i_1 _09961_ (.A0(_05627_),
    .A1(_05634_),
    .S(_05472_),
    .Y(_05635_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(reset_hash),
    .B(\w[1][9] ),
    .Y(_05636_));
 sky130_fd_sc_hd__o21ai_0 _09963_ (.A1(_05482_),
    .A2(_05635_),
    .B1(_05636_),
    .Y(_00063_));
 sky130_fd_sc_hd__mux4_2 _09964_ (.A0(\w[19][10] ),
    .A1(\w[23][10] ),
    .A2(\w[17][10] ),
    .A3(\w[21][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05637_));
 sky130_fd_sc_hd__mux4_2 _09965_ (.A0(\w[27][10] ),
    .A1(\w[31][10] ),
    .A2(\w[25][10] ),
    .A3(\w[29][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05638_));
 sky130_fd_sc_hd__mux4_2 _09966_ (.A0(\w[3][10] ),
    .A1(\w[7][10] ),
    .A2(\w[1][10] ),
    .A3(\w[5][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05639_));
 sky130_fd_sc_hd__mux4_2 _09968_ (.A0(\w[11][10] ),
    .A1(\w[15][10] ),
    .A2(\w[9][10] ),
    .A3(\w[13][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05641_));
 sky130_fd_sc_hd__mux4_2 _09969_ (.A0(_05637_),
    .A1(_05638_),
    .A2(_05639_),
    .A3(_05641_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05642_));
 sky130_fd_sc_hd__mux4_2 _09970_ (.A0(\w[51][10] ),
    .A1(\w[55][10] ),
    .A2(\w[49][10] ),
    .A3(\w[53][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05643_));
 sky130_fd_sc_hd__mux4_2 _09972_ (.A0(\w[59][10] ),
    .A1(\w[63][10] ),
    .A2(\w[57][10] ),
    .A3(\w[61][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05645_));
 sky130_fd_sc_hd__mux4_2 _09973_ (.A0(\w[35][10] ),
    .A1(\w[39][10] ),
    .A2(\w[33][10] ),
    .A3(\w[37][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05646_));
 sky130_fd_sc_hd__mux4_2 _09974_ (.A0(\w[43][10] ),
    .A1(\w[47][10] ),
    .A2(\w[41][10] ),
    .A3(\w[45][10] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05647_));
 sky130_fd_sc_hd__mux4_2 _09975_ (.A0(_05643_),
    .A1(_05645_),
    .A2(_05646_),
    .A3(_05647_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05648_));
 sky130_fd_sc_hd__mux2i_1 _09976_ (.A0(_05642_),
    .A1(_05648_),
    .S(_05472_),
    .Y(_05649_));
 sky130_fd_sc_hd__nand2_1 _09977_ (.A(reset_hash),
    .B(\w[1][10] ),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_0 _09978_ (.A1(_05482_),
    .A2(_05649_),
    .B1(_05650_),
    .Y(_00033_));
 sky130_fd_sc_hd__mux4_2 _09979_ (.A0(\w[19][11] ),
    .A1(\w[23][11] ),
    .A2(\w[17][11] ),
    .A3(\w[21][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05651_));
 sky130_fd_sc_hd__mux4_2 _09980_ (.A0(\w[27][11] ),
    .A1(\w[31][11] ),
    .A2(\w[25][11] ),
    .A3(\w[29][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05652_));
 sky130_fd_sc_hd__mux4_2 _09981_ (.A0(\w[3][11] ),
    .A1(\w[7][11] ),
    .A2(\w[1][11] ),
    .A3(\w[5][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05653_));
 sky130_fd_sc_hd__mux4_2 _09982_ (.A0(\w[11][11] ),
    .A1(\w[15][11] ),
    .A2(\w[9][11] ),
    .A3(\w[13][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05654_));
 sky130_fd_sc_hd__mux4_2 _09983_ (.A0(_05651_),
    .A1(_05652_),
    .A2(_05653_),
    .A3(_05654_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05655_));
 sky130_fd_sc_hd__mux4_2 _09984_ (.A0(\w[51][11] ),
    .A1(\w[55][11] ),
    .A2(\w[49][11] ),
    .A3(\w[53][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05656_));
 sky130_fd_sc_hd__mux4_2 _09985_ (.A0(\w[59][11] ),
    .A1(\w[63][11] ),
    .A2(\w[57][11] ),
    .A3(\w[61][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05657_));
 sky130_fd_sc_hd__mux4_2 _09986_ (.A0(\w[35][11] ),
    .A1(\w[39][11] ),
    .A2(\w[33][11] ),
    .A3(\w[37][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05658_));
 sky130_fd_sc_hd__mux4_2 _09987_ (.A0(\w[43][11] ),
    .A1(\w[47][11] ),
    .A2(\w[41][11] ),
    .A3(\w[45][11] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05659_));
 sky130_fd_sc_hd__mux4_2 _09988_ (.A0(_05656_),
    .A1(_05657_),
    .A2(_05658_),
    .A3(_05659_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05660_));
 sky130_fd_sc_hd__mux2i_1 _09989_ (.A0(_05655_),
    .A1(_05660_),
    .S(_05472_),
    .Y(_05661_));
 sky130_fd_sc_hd__nand2_1 _09990_ (.A(reset_hash),
    .B(\w[1][11] ),
    .Y(_05662_));
 sky130_fd_sc_hd__o21ai_0 _09991_ (.A1(_05482_),
    .A2(_05661_),
    .B1(_05662_),
    .Y(_00034_));
 sky130_fd_sc_hd__mux4_2 _09993_ (.A0(\w[19][12] ),
    .A1(\w[23][12] ),
    .A2(\w[17][12] ),
    .A3(\w[21][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05664_));
 sky130_fd_sc_hd__mux4_2 _09995_ (.A0(\w[27][12] ),
    .A1(\w[31][12] ),
    .A2(\w[25][12] ),
    .A3(\w[29][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05666_));
 sky130_fd_sc_hd__mux4_2 _09996_ (.A0(\w[3][12] ),
    .A1(\w[7][12] ),
    .A2(\w[1][12] ),
    .A3(\w[5][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05667_));
 sky130_fd_sc_hd__mux4_2 _09997_ (.A0(\w[11][12] ),
    .A1(\w[15][12] ),
    .A2(\w[9][12] ),
    .A3(\w[13][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05668_));
 sky130_fd_sc_hd__mux4_2 _09998_ (.A0(_05664_),
    .A1(_05666_),
    .A2(_05667_),
    .A3(_05668_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05669_));
 sky130_fd_sc_hd__mux4_2 _09999_ (.A0(\w[51][12] ),
    .A1(\w[55][12] ),
    .A2(\w[49][12] ),
    .A3(\w[53][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05670_));
 sky130_fd_sc_hd__mux4_2 _10000_ (.A0(\w[59][12] ),
    .A1(\w[63][12] ),
    .A2(\w[57][12] ),
    .A3(\w[61][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05671_));
 sky130_fd_sc_hd__mux4_2 _10001_ (.A0(\w[35][12] ),
    .A1(\w[39][12] ),
    .A2(\w[33][12] ),
    .A3(\w[37][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05672_));
 sky130_fd_sc_hd__mux4_2 _10002_ (.A0(\w[43][12] ),
    .A1(\w[47][12] ),
    .A2(\w[41][12] ),
    .A3(\w[45][12] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05673_));
 sky130_fd_sc_hd__mux4_2 _10004_ (.A0(_05670_),
    .A1(_05671_),
    .A2(_05672_),
    .A3(_05673_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05675_));
 sky130_fd_sc_hd__mux2i_1 _10005_ (.A0(_05669_),
    .A1(_05675_),
    .S(_05472_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand2_1 _10006_ (.A(reset_hash),
    .B(\w[1][12] ),
    .Y(_05677_));
 sky130_fd_sc_hd__o21ai_0 _10007_ (.A1(_05482_),
    .A2(_05676_),
    .B1(_05677_),
    .Y(_00035_));
 sky130_fd_sc_hd__mux4_2 _10008_ (.A0(\w[19][13] ),
    .A1(\w[23][13] ),
    .A2(\w[17][13] ),
    .A3(\w[21][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05678_));
 sky130_fd_sc_hd__mux4_2 _10010_ (.A0(\w[27][13] ),
    .A1(\w[31][13] ),
    .A2(\w[25][13] ),
    .A3(\w[29][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05680_));
 sky130_fd_sc_hd__mux4_2 _10011_ (.A0(\w[3][13] ),
    .A1(\w[7][13] ),
    .A2(\w[1][13] ),
    .A3(\w[5][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05681_));
 sky130_fd_sc_hd__mux4_2 _10012_ (.A0(\w[11][13] ),
    .A1(\w[15][13] ),
    .A2(\w[9][13] ),
    .A3(\w[13][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05682_));
 sky130_fd_sc_hd__mux4_2 _10013_ (.A0(_05678_),
    .A1(_05680_),
    .A2(_05681_),
    .A3(_05682_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05683_));
 sky130_fd_sc_hd__mux4_2 _10014_ (.A0(\w[51][13] ),
    .A1(\w[55][13] ),
    .A2(\w[49][13] ),
    .A3(\w[53][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05684_));
 sky130_fd_sc_hd__mux4_2 _10015_ (.A0(\w[59][13] ),
    .A1(\w[63][13] ),
    .A2(\w[57][13] ),
    .A3(\w[61][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05685_));
 sky130_fd_sc_hd__mux4_2 _10017_ (.A0(\w[35][13] ),
    .A1(\w[39][13] ),
    .A2(\w[33][13] ),
    .A3(\w[37][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05687_));
 sky130_fd_sc_hd__mux4_2 _10018_ (.A0(\w[43][13] ),
    .A1(\w[47][13] ),
    .A2(\w[41][13] ),
    .A3(\w[45][13] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05688_));
 sky130_fd_sc_hd__mux4_2 _10019_ (.A0(_05684_),
    .A1(_05685_),
    .A2(_05687_),
    .A3(_05688_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05689_));
 sky130_fd_sc_hd__mux2i_1 _10020_ (.A0(_05683_),
    .A1(_05689_),
    .S(_05472_),
    .Y(_05690_));
 sky130_fd_sc_hd__nand2_1 _10021_ (.A(reset_hash),
    .B(\w[1][13] ),
    .Y(_05691_));
 sky130_fd_sc_hd__o21ai_0 _10022_ (.A1(_05482_),
    .A2(_05690_),
    .B1(_05691_),
    .Y(_00036_));
 sky130_fd_sc_hd__mux4_2 _10023_ (.A0(\w[19][14] ),
    .A1(\w[23][14] ),
    .A2(\w[17][14] ),
    .A3(\w[21][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05692_));
 sky130_fd_sc_hd__mux4_2 _10024_ (.A0(\w[27][14] ),
    .A1(\w[31][14] ),
    .A2(\w[25][14] ),
    .A3(\w[29][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05693_));
 sky130_fd_sc_hd__mux4_2 _10025_ (.A0(\w[3][14] ),
    .A1(\w[7][14] ),
    .A2(\w[1][14] ),
    .A3(\w[5][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05694_));
 sky130_fd_sc_hd__mux4_2 _10026_ (.A0(\w[11][14] ),
    .A1(\w[15][14] ),
    .A2(\w[9][14] ),
    .A3(\w[13][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05695_));
 sky130_fd_sc_hd__mux4_2 _10028_ (.A0(_05692_),
    .A1(_05693_),
    .A2(_05694_),
    .A3(_05695_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05697_));
 sky130_fd_sc_hd__mux4_2 _10029_ (.A0(\w[51][14] ),
    .A1(\w[55][14] ),
    .A2(\w[49][14] ),
    .A3(\w[53][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05698_));
 sky130_fd_sc_hd__mux4_2 _10030_ (.A0(\w[59][14] ),
    .A1(\w[63][14] ),
    .A2(\w[57][14] ),
    .A3(\w[61][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05699_));
 sky130_fd_sc_hd__mux4_2 _10032_ (.A0(\w[35][14] ),
    .A1(\w[39][14] ),
    .A2(\w[33][14] ),
    .A3(\w[37][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05701_));
 sky130_fd_sc_hd__mux4_2 _10033_ (.A0(\w[43][14] ),
    .A1(\w[47][14] ),
    .A2(\w[41][14] ),
    .A3(\w[45][14] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05702_));
 sky130_fd_sc_hd__mux4_2 _10034_ (.A0(_05698_),
    .A1(_05699_),
    .A2(_05701_),
    .A3(_05702_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05703_));
 sky130_fd_sc_hd__mux2i_1 _10035_ (.A0(_05697_),
    .A1(_05703_),
    .S(_05472_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(reset_hash),
    .B(\w[1][14] ),
    .Y(_05706_));
 sky130_fd_sc_hd__o21ai_0 _10038_ (.A1(_05482_),
    .A2(_05704_),
    .B1(_05706_),
    .Y(_00037_));
 sky130_fd_sc_hd__mux4_2 _10039_ (.A0(\w[19][15] ),
    .A1(\w[23][15] ),
    .A2(\w[17][15] ),
    .A3(\w[21][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05707_));
 sky130_fd_sc_hd__mux4_2 _10040_ (.A0(\w[27][15] ),
    .A1(\w[31][15] ),
    .A2(\w[25][15] ),
    .A3(\w[29][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05708_));
 sky130_fd_sc_hd__mux4_2 _10041_ (.A0(\w[3][15] ),
    .A1(\w[7][15] ),
    .A2(\w[1][15] ),
    .A3(\w[5][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05709_));
 sky130_fd_sc_hd__mux4_2 _10042_ (.A0(\w[11][15] ),
    .A1(\w[15][15] ),
    .A2(\w[9][15] ),
    .A3(\w[13][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05710_));
 sky130_fd_sc_hd__mux4_2 _10043_ (.A0(_05707_),
    .A1(_05708_),
    .A2(_05709_),
    .A3(_05710_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05711_));
 sky130_fd_sc_hd__mux4_2 _10045_ (.A0(\w[51][15] ),
    .A1(\w[55][15] ),
    .A2(\w[49][15] ),
    .A3(\w[53][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05713_));
 sky130_fd_sc_hd__mux4_2 _10046_ (.A0(\w[59][15] ),
    .A1(\w[63][15] ),
    .A2(\w[57][15] ),
    .A3(\w[61][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05714_));
 sky130_fd_sc_hd__mux4_2 _10047_ (.A0(\w[35][15] ),
    .A1(\w[39][15] ),
    .A2(\w[33][15] ),
    .A3(\w[37][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05715_));
 sky130_fd_sc_hd__mux4_2 _10048_ (.A0(\w[43][15] ),
    .A1(\w[47][15] ),
    .A2(\w[41][15] ),
    .A3(\w[45][15] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05716_));
 sky130_fd_sc_hd__mux4_2 _10050_ (.A0(_05713_),
    .A1(_05714_),
    .A2(_05715_),
    .A3(_05716_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05718_));
 sky130_fd_sc_hd__mux2i_1 _10051_ (.A0(_05711_),
    .A1(_05718_),
    .S(_05472_),
    .Y(_05719_));
 sky130_fd_sc_hd__nand2_1 _10052_ (.A(reset_hash),
    .B(\w[1][15] ),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ai_0 _10053_ (.A1(_05482_),
    .A2(_05719_),
    .B1(_05720_),
    .Y(_00038_));
 sky130_fd_sc_hd__mux4_2 _10054_ (.A0(\w[19][16] ),
    .A1(\w[23][16] ),
    .A2(\w[17][16] ),
    .A3(\w[21][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05721_));
 sky130_fd_sc_hd__mux4_2 _10055_ (.A0(\w[27][16] ),
    .A1(\w[31][16] ),
    .A2(\w[25][16] ),
    .A3(\w[29][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05722_));
 sky130_fd_sc_hd__mux4_2 _10057_ (.A0(\w[3][16] ),
    .A1(\w[7][16] ),
    .A2(\w[1][16] ),
    .A3(\w[5][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05724_));
 sky130_fd_sc_hd__mux4_2 _10058_ (.A0(\w[11][16] ),
    .A1(\w[15][16] ),
    .A2(\w[9][16] ),
    .A3(\w[13][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05725_));
 sky130_fd_sc_hd__mux4_2 _10060_ (.A0(_05721_),
    .A1(_05722_),
    .A2(_05724_),
    .A3(_05725_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05727_));
 sky130_fd_sc_hd__mux4_2 _10062_ (.A0(\w[51][16] ),
    .A1(\w[55][16] ),
    .A2(\w[49][16] ),
    .A3(\w[53][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05729_));
 sky130_fd_sc_hd__mux4_2 _10063_ (.A0(\w[59][16] ),
    .A1(\w[63][16] ),
    .A2(\w[57][16] ),
    .A3(\w[61][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05730_));
 sky130_fd_sc_hd__mux4_2 _10064_ (.A0(\w[35][16] ),
    .A1(\w[39][16] ),
    .A2(\w[33][16] ),
    .A3(\w[37][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05731_));
 sky130_fd_sc_hd__mux4_2 _10065_ (.A0(\w[43][16] ),
    .A1(\w[47][16] ),
    .A2(\w[41][16] ),
    .A3(\w[45][16] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05732_));
 sky130_fd_sc_hd__mux4_2 _10066_ (.A0(_05729_),
    .A1(_05730_),
    .A2(_05731_),
    .A3(_05732_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05733_));
 sky130_fd_sc_hd__mux2i_1 _10067_ (.A0(_05727_),
    .A1(_05733_),
    .S(_05472_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand2_1 _10068_ (.A(reset_hash),
    .B(\w[1][16] ),
    .Y(_05735_));
 sky130_fd_sc_hd__o21ai_0 _10069_ (.A1(_05482_),
    .A2(_05734_),
    .B1(_05735_),
    .Y(_00039_));
 sky130_fd_sc_hd__mux4_2 _10071_ (.A0(\w[19][17] ),
    .A1(\w[23][17] ),
    .A2(\w[17][17] ),
    .A3(\w[21][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05737_));
 sky130_fd_sc_hd__mux4_2 _10072_ (.A0(\w[27][17] ),
    .A1(\w[31][17] ),
    .A2(\w[25][17] ),
    .A3(\w[29][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05738_));
 sky130_fd_sc_hd__mux4_2 _10074_ (.A0(\w[3][17] ),
    .A1(\w[7][17] ),
    .A2(\w[1][17] ),
    .A3(\w[5][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05740_));
 sky130_fd_sc_hd__mux4_2 _10075_ (.A0(\w[11][17] ),
    .A1(\w[15][17] ),
    .A2(\w[9][17] ),
    .A3(\w[13][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05741_));
 sky130_fd_sc_hd__mux4_2 _10076_ (.A0(_05737_),
    .A1(_05738_),
    .A2(_05740_),
    .A3(_05741_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05742_));
 sky130_fd_sc_hd__mux4_2 _10077_ (.A0(\w[51][17] ),
    .A1(\w[55][17] ),
    .A2(\w[49][17] ),
    .A3(\w[53][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05743_));
 sky130_fd_sc_hd__mux4_2 _10078_ (.A0(\w[59][17] ),
    .A1(\w[63][17] ),
    .A2(\w[57][17] ),
    .A3(\w[61][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05744_));
 sky130_fd_sc_hd__mux4_2 _10079_ (.A0(\w[35][17] ),
    .A1(\w[39][17] ),
    .A2(\w[33][17] ),
    .A3(\w[37][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05745_));
 sky130_fd_sc_hd__mux4_2 _10080_ (.A0(\w[43][17] ),
    .A1(\w[47][17] ),
    .A2(\w[41][17] ),
    .A3(\w[45][17] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05746_));
 sky130_fd_sc_hd__mux4_2 _10081_ (.A0(_05743_),
    .A1(_05744_),
    .A2(_05745_),
    .A3(_05746_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05747_));
 sky130_fd_sc_hd__mux2i_1 _10082_ (.A0(_05742_),
    .A1(_05747_),
    .S(_05472_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand2_1 _10083_ (.A(reset_hash),
    .B(\w[1][17] ),
    .Y(_05749_));
 sky130_fd_sc_hd__o21ai_0 _10084_ (.A1(_05482_),
    .A2(_05748_),
    .B1(_05749_),
    .Y(_00040_));
 sky130_fd_sc_hd__mux4_2 _10086_ (.A0(\w[19][18] ),
    .A1(\w[23][18] ),
    .A2(\w[17][18] ),
    .A3(\w[21][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05751_));
 sky130_fd_sc_hd__mux4_2 _10087_ (.A0(\w[27][18] ),
    .A1(\w[31][18] ),
    .A2(\w[25][18] ),
    .A3(\w[29][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05752_));
 sky130_fd_sc_hd__mux4_2 _10088_ (.A0(\w[3][18] ),
    .A1(\w[7][18] ),
    .A2(\w[1][18] ),
    .A3(\w[5][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05753_));
 sky130_fd_sc_hd__mux4_2 _10089_ (.A0(\w[11][18] ),
    .A1(\w[15][18] ),
    .A2(\w[9][18] ),
    .A3(\w[13][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05754_));
 sky130_fd_sc_hd__mux4_2 _10090_ (.A0(_05751_),
    .A1(_05752_),
    .A2(_05753_),
    .A3(_05754_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05755_));
 sky130_fd_sc_hd__mux4_2 _10091_ (.A0(\w[51][18] ),
    .A1(\w[55][18] ),
    .A2(\w[49][18] ),
    .A3(\w[53][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05756_));
 sky130_fd_sc_hd__mux4_2 _10092_ (.A0(\w[59][18] ),
    .A1(\w[63][18] ),
    .A2(\w[57][18] ),
    .A3(\w[61][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05757_));
 sky130_fd_sc_hd__mux4_2 _10093_ (.A0(\w[35][18] ),
    .A1(\w[39][18] ),
    .A2(\w[33][18] ),
    .A3(\w[37][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05758_));
 sky130_fd_sc_hd__mux4_2 _10095_ (.A0(\w[43][18] ),
    .A1(\w[47][18] ),
    .A2(\w[41][18] ),
    .A3(\w[45][18] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05760_));
 sky130_fd_sc_hd__mux4_2 _10096_ (.A0(_05756_),
    .A1(_05757_),
    .A2(_05758_),
    .A3(_05760_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05761_));
 sky130_fd_sc_hd__mux2i_1 _10098_ (.A0(_05755_),
    .A1(_05761_),
    .S(_05472_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2_1 _10099_ (.A(reset_hash),
    .B(\w[1][18] ),
    .Y(_05764_));
 sky130_fd_sc_hd__o21ai_0 _10100_ (.A1(_05482_),
    .A2(_05763_),
    .B1(_05764_),
    .Y(_00041_));
 sky130_fd_sc_hd__mux4_2 _10101_ (.A0(\w[19][19] ),
    .A1(\w[23][19] ),
    .A2(\w[17][19] ),
    .A3(\w[21][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05765_));
 sky130_fd_sc_hd__mux4_2 _10102_ (.A0(\w[27][19] ),
    .A1(\w[31][19] ),
    .A2(\w[25][19] ),
    .A3(\w[29][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05766_));
 sky130_fd_sc_hd__mux4_2 _10103_ (.A0(\w[3][19] ),
    .A1(\w[7][19] ),
    .A2(\w[1][19] ),
    .A3(\w[5][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05767_));
 sky130_fd_sc_hd__mux4_2 _10105_ (.A0(\w[11][19] ),
    .A1(\w[15][19] ),
    .A2(\w[9][19] ),
    .A3(\w[13][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05769_));
 sky130_fd_sc_hd__mux4_2 _10106_ (.A0(_05765_),
    .A1(_05766_),
    .A2(_05767_),
    .A3(_05769_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05770_));
 sky130_fd_sc_hd__mux4_2 _10107_ (.A0(\w[51][19] ),
    .A1(\w[55][19] ),
    .A2(\w[49][19] ),
    .A3(\w[53][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05771_));
 sky130_fd_sc_hd__mux4_2 _10109_ (.A0(\w[59][19] ),
    .A1(\w[63][19] ),
    .A2(\w[57][19] ),
    .A3(\w[61][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05773_));
 sky130_fd_sc_hd__mux4_2 _10110_ (.A0(\w[35][19] ),
    .A1(\w[39][19] ),
    .A2(\w[33][19] ),
    .A3(\w[37][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05774_));
 sky130_fd_sc_hd__mux4_2 _10112_ (.A0(\w[43][19] ),
    .A1(\w[47][19] ),
    .A2(\w[41][19] ),
    .A3(\w[45][19] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05776_));
 sky130_fd_sc_hd__mux4_2 _10113_ (.A0(_05771_),
    .A1(_05773_),
    .A2(_05774_),
    .A3(_05776_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05777_));
 sky130_fd_sc_hd__mux2i_1 _10114_ (.A0(_05770_),
    .A1(_05777_),
    .S(_05472_),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_1 _10115_ (.A(reset_hash),
    .B(\w[1][19] ),
    .Y(_05779_));
 sky130_fd_sc_hd__o21ai_0 _10116_ (.A1(_05482_),
    .A2(_05778_),
    .B1(_05779_),
    .Y(_00042_));
 sky130_fd_sc_hd__mux4_2 _10117_ (.A0(\w[19][20] ),
    .A1(\w[23][20] ),
    .A2(\w[17][20] ),
    .A3(\w[21][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05780_));
 sky130_fd_sc_hd__mux4_2 _10118_ (.A0(\w[27][20] ),
    .A1(\w[31][20] ),
    .A2(\w[25][20] ),
    .A3(\w[29][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05781_));
 sky130_fd_sc_hd__mux4_2 _10119_ (.A0(\w[3][20] ),
    .A1(\w[7][20] ),
    .A2(\w[1][20] ),
    .A3(\w[5][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05782_));
 sky130_fd_sc_hd__mux4_2 _10121_ (.A0(\w[11][20] ),
    .A1(\w[15][20] ),
    .A2(\w[9][20] ),
    .A3(\w[13][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05784_));
 sky130_fd_sc_hd__mux4_2 _10122_ (.A0(_05780_),
    .A1(_05781_),
    .A2(_05782_),
    .A3(_05784_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05785_));
 sky130_fd_sc_hd__mux4_2 _10123_ (.A0(\w[51][20] ),
    .A1(\w[55][20] ),
    .A2(\w[49][20] ),
    .A3(\w[53][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05786_));
 sky130_fd_sc_hd__mux4_2 _10125_ (.A0(\w[59][20] ),
    .A1(\w[63][20] ),
    .A2(\w[57][20] ),
    .A3(\w[61][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05788_));
 sky130_fd_sc_hd__mux4_2 _10126_ (.A0(\w[35][20] ),
    .A1(\w[39][20] ),
    .A2(\w[33][20] ),
    .A3(\w[37][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05789_));
 sky130_fd_sc_hd__mux4_2 _10127_ (.A0(\w[43][20] ),
    .A1(\w[47][20] ),
    .A2(\w[41][20] ),
    .A3(\w[45][20] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05790_));
 sky130_fd_sc_hd__mux4_2 _10128_ (.A0(_05786_),
    .A1(_05788_),
    .A2(_05789_),
    .A3(_05790_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05791_));
 sky130_fd_sc_hd__mux2i_1 _10129_ (.A0(_05785_),
    .A1(_05791_),
    .S(_05472_),
    .Y(_05792_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(reset_hash),
    .B(\w[1][20] ),
    .Y(_05793_));
 sky130_fd_sc_hd__o21ai_0 _10131_ (.A1(_05482_),
    .A2(_05792_),
    .B1(_05793_),
    .Y(_00044_));
 sky130_fd_sc_hd__mux4_2 _10132_ (.A0(\w[19][21] ),
    .A1(\w[23][21] ),
    .A2(\w[17][21] ),
    .A3(\w[21][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05794_));
 sky130_fd_sc_hd__mux4_2 _10133_ (.A0(\w[27][21] ),
    .A1(\w[31][21] ),
    .A2(\w[25][21] ),
    .A3(\w[29][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05795_));
 sky130_fd_sc_hd__mux4_2 _10134_ (.A0(\w[3][21] ),
    .A1(\w[7][21] ),
    .A2(\w[1][21] ),
    .A3(\w[5][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05796_));
 sky130_fd_sc_hd__mux4_2 _10135_ (.A0(\w[11][21] ),
    .A1(\w[15][21] ),
    .A2(\w[9][21] ),
    .A3(\w[13][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05797_));
 sky130_fd_sc_hd__mux4_2 _10136_ (.A0(_05794_),
    .A1(_05795_),
    .A2(_05796_),
    .A3(_05797_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05798_));
 sky130_fd_sc_hd__mux4_2 _10137_ (.A0(\w[51][21] ),
    .A1(\w[55][21] ),
    .A2(\w[49][21] ),
    .A3(\w[53][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05799_));
 sky130_fd_sc_hd__mux4_2 _10138_ (.A0(\w[59][21] ),
    .A1(\w[63][21] ),
    .A2(\w[57][21] ),
    .A3(\w[61][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05800_));
 sky130_fd_sc_hd__mux4_2 _10139_ (.A0(\w[35][21] ),
    .A1(\w[39][21] ),
    .A2(\w[33][21] ),
    .A3(\w[37][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05801_));
 sky130_fd_sc_hd__mux4_2 _10140_ (.A0(\w[43][21] ),
    .A1(\w[47][21] ),
    .A2(\w[41][21] ),
    .A3(\w[45][21] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05802_));
 sky130_fd_sc_hd__mux4_2 _10141_ (.A0(_05799_),
    .A1(_05800_),
    .A2(_05801_),
    .A3(_05802_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05803_));
 sky130_fd_sc_hd__mux2i_1 _10142_ (.A0(_05798_),
    .A1(_05803_),
    .S(_05472_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_1 _10143_ (.A(reset_hash),
    .B(\w[1][21] ),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_0 _10144_ (.A1(_05482_),
    .A2(_05804_),
    .B1(_05805_),
    .Y(_00045_));
 sky130_fd_sc_hd__mux4_2 _10146_ (.A0(\w[19][22] ),
    .A1(\w[23][22] ),
    .A2(\w[17][22] ),
    .A3(\w[21][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05807_));
 sky130_fd_sc_hd__mux4_2 _10148_ (.A0(\w[27][22] ),
    .A1(\w[31][22] ),
    .A2(\w[25][22] ),
    .A3(\w[29][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05809_));
 sky130_fd_sc_hd__mux4_2 _10149_ (.A0(\w[3][22] ),
    .A1(\w[7][22] ),
    .A2(\w[1][22] ),
    .A3(\w[5][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05810_));
 sky130_fd_sc_hd__mux4_2 _10150_ (.A0(\w[11][22] ),
    .A1(\w[15][22] ),
    .A2(\w[9][22] ),
    .A3(\w[13][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05811_));
 sky130_fd_sc_hd__mux4_2 _10151_ (.A0(_05807_),
    .A1(_05809_),
    .A2(_05810_),
    .A3(_05811_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05812_));
 sky130_fd_sc_hd__mux4_2 _10152_ (.A0(\w[51][22] ),
    .A1(\w[55][22] ),
    .A2(\w[49][22] ),
    .A3(\w[53][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05813_));
 sky130_fd_sc_hd__mux4_2 _10153_ (.A0(\w[59][22] ),
    .A1(\w[63][22] ),
    .A2(\w[57][22] ),
    .A3(\w[61][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05814_));
 sky130_fd_sc_hd__mux4_2 _10154_ (.A0(\w[35][22] ),
    .A1(\w[39][22] ),
    .A2(\w[33][22] ),
    .A3(\w[37][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05815_));
 sky130_fd_sc_hd__mux4_2 _10155_ (.A0(\w[43][22] ),
    .A1(\w[47][22] ),
    .A2(\w[41][22] ),
    .A3(\w[45][22] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05816_));
 sky130_fd_sc_hd__mux4_2 _10157_ (.A0(_05813_),
    .A1(_05814_),
    .A2(_05815_),
    .A3(_05816_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05818_));
 sky130_fd_sc_hd__mux2i_1 _10158_ (.A0(_05812_),
    .A1(_05818_),
    .S(_05472_),
    .Y(_05819_));
 sky130_fd_sc_hd__nand2_1 _10159_ (.A(reset_hash),
    .B(\w[1][22] ),
    .Y(_05820_));
 sky130_fd_sc_hd__o21ai_0 _10160_ (.A1(_05482_),
    .A2(_05819_),
    .B1(_05820_),
    .Y(_00046_));
 sky130_fd_sc_hd__mux4_2 _10161_ (.A0(\w[19][23] ),
    .A1(\w[23][23] ),
    .A2(\w[17][23] ),
    .A3(\w[21][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05821_));
 sky130_fd_sc_hd__mux4_2 _10162_ (.A0(\w[27][23] ),
    .A1(\w[31][23] ),
    .A2(\w[25][23] ),
    .A3(\w[29][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05822_));
 sky130_fd_sc_hd__mux4_2 _10163_ (.A0(\w[3][23] ),
    .A1(\w[7][23] ),
    .A2(\w[1][23] ),
    .A3(\w[5][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05823_));
 sky130_fd_sc_hd__mux4_2 _10164_ (.A0(\w[11][23] ),
    .A1(\w[15][23] ),
    .A2(\w[9][23] ),
    .A3(\w[13][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05824_));
 sky130_fd_sc_hd__mux4_2 _10165_ (.A0(_05821_),
    .A1(_05822_),
    .A2(_05823_),
    .A3(_05824_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05825_));
 sky130_fd_sc_hd__mux4_2 _10166_ (.A0(\w[51][23] ),
    .A1(\w[55][23] ),
    .A2(\w[49][23] ),
    .A3(\w[53][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05826_));
 sky130_fd_sc_hd__mux4_2 _10167_ (.A0(\w[59][23] ),
    .A1(\w[63][23] ),
    .A2(\w[57][23] ),
    .A3(\w[61][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05827_));
 sky130_fd_sc_hd__mux4_2 _10168_ (.A0(\w[35][23] ),
    .A1(\w[39][23] ),
    .A2(\w[33][23] ),
    .A3(\w[37][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05828_));
 sky130_fd_sc_hd__mux4_2 _10169_ (.A0(\w[43][23] ),
    .A1(\w[47][23] ),
    .A2(\w[41][23] ),
    .A3(\w[45][23] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05829_));
 sky130_fd_sc_hd__mux4_2 _10170_ (.A0(_05826_),
    .A1(_05827_),
    .A2(_05828_),
    .A3(_05829_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05830_));
 sky130_fd_sc_hd__mux2i_1 _10171_ (.A0(_05825_),
    .A1(_05830_),
    .S(_05472_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand2_1 _10172_ (.A(reset_hash),
    .B(\w[1][23] ),
    .Y(_05832_));
 sky130_fd_sc_hd__o21ai_0 _10173_ (.A1(_05482_),
    .A2(_05831_),
    .B1(_05832_),
    .Y(_00047_));
 sky130_fd_sc_hd__mux4_2 _10174_ (.A0(\w[19][24] ),
    .A1(\w[23][24] ),
    .A2(\w[17][24] ),
    .A3(\w[21][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05833_));
 sky130_fd_sc_hd__mux4_2 _10175_ (.A0(\w[27][24] ),
    .A1(\w[31][24] ),
    .A2(\w[25][24] ),
    .A3(\w[29][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05834_));
 sky130_fd_sc_hd__mux4_2 _10176_ (.A0(\w[3][24] ),
    .A1(\w[7][24] ),
    .A2(\w[1][24] ),
    .A3(\w[5][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05835_));
 sky130_fd_sc_hd__mux4_2 _10177_ (.A0(\w[11][24] ),
    .A1(\w[15][24] ),
    .A2(\w[9][24] ),
    .A3(\w[13][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05836_));
 sky130_fd_sc_hd__mux4_2 _10178_ (.A0(_05833_),
    .A1(_05834_),
    .A2(_05835_),
    .A3(_05836_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05837_));
 sky130_fd_sc_hd__mux4_2 _10179_ (.A0(\w[51][24] ),
    .A1(\w[55][24] ),
    .A2(\w[49][24] ),
    .A3(\w[53][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05838_));
 sky130_fd_sc_hd__mux4_2 _10180_ (.A0(\w[59][24] ),
    .A1(\w[63][24] ),
    .A2(\w[57][24] ),
    .A3(\w[61][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05839_));
 sky130_fd_sc_hd__mux4_2 _10181_ (.A0(\w[35][24] ),
    .A1(\w[39][24] ),
    .A2(\w[33][24] ),
    .A3(\w[37][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05840_));
 sky130_fd_sc_hd__mux4_2 _10182_ (.A0(\w[43][24] ),
    .A1(\w[47][24] ),
    .A2(\w[41][24] ),
    .A3(\w[45][24] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05841_));
 sky130_fd_sc_hd__mux4_2 _10183_ (.A0(_05838_),
    .A1(_05839_),
    .A2(_05840_),
    .A3(_05841_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05842_));
 sky130_fd_sc_hd__mux2i_1 _10184_ (.A0(_05837_),
    .A1(_05842_),
    .S(_05472_),
    .Y(_05843_));
 sky130_fd_sc_hd__nand2_1 _10186_ (.A(reset_hash),
    .B(\w[1][24] ),
    .Y(_05845_));
 sky130_fd_sc_hd__o21ai_0 _10187_ (.A1(_05482_),
    .A2(_05843_),
    .B1(_05845_),
    .Y(_00048_));
 sky130_fd_sc_hd__mux4_2 _10188_ (.A0(\w[19][25] ),
    .A1(\w[23][25] ),
    .A2(\w[17][25] ),
    .A3(\w[21][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05846_));
 sky130_fd_sc_hd__mux4_2 _10189_ (.A0(\w[27][25] ),
    .A1(\w[31][25] ),
    .A2(\w[25][25] ),
    .A3(\w[29][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05847_));
 sky130_fd_sc_hd__mux4_2 _10190_ (.A0(\w[3][25] ),
    .A1(\w[7][25] ),
    .A2(\w[1][25] ),
    .A3(\w[5][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05848_));
 sky130_fd_sc_hd__mux4_2 _10191_ (.A0(\w[11][25] ),
    .A1(\w[15][25] ),
    .A2(\w[9][25] ),
    .A3(\w[13][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05849_));
 sky130_fd_sc_hd__mux4_2 _10192_ (.A0(_05846_),
    .A1(_05847_),
    .A2(_05848_),
    .A3(_05849_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05850_));
 sky130_fd_sc_hd__mux4_2 _10193_ (.A0(\w[51][25] ),
    .A1(\w[55][25] ),
    .A2(\w[49][25] ),
    .A3(\w[53][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05851_));
 sky130_fd_sc_hd__mux4_2 _10194_ (.A0(\w[59][25] ),
    .A1(\w[63][25] ),
    .A2(\w[57][25] ),
    .A3(\w[61][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05852_));
 sky130_fd_sc_hd__mux4_2 _10195_ (.A0(\w[35][25] ),
    .A1(\w[39][25] ),
    .A2(\w[33][25] ),
    .A3(\w[37][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05853_));
 sky130_fd_sc_hd__mux4_2 _10196_ (.A0(\w[43][25] ),
    .A1(\w[47][25] ),
    .A2(\w[41][25] ),
    .A3(\w[45][25] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05854_));
 sky130_fd_sc_hd__mux4_2 _10197_ (.A0(_05851_),
    .A1(_05852_),
    .A2(_05853_),
    .A3(_05854_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05855_));
 sky130_fd_sc_hd__mux2i_1 _10198_ (.A0(_05850_),
    .A1(_05855_),
    .S(_05472_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _10199_ (.A(reset_hash),
    .B(\w[1][25] ),
    .Y(_05857_));
 sky130_fd_sc_hd__o21ai_0 _10200_ (.A1(_05482_),
    .A2(_05856_),
    .B1(_05857_),
    .Y(_00049_));
 sky130_fd_sc_hd__mux4_2 _10201_ (.A0(\w[19][26] ),
    .A1(\w[23][26] ),
    .A2(\w[17][26] ),
    .A3(\w[21][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05858_));
 sky130_fd_sc_hd__mux4_2 _10202_ (.A0(\w[27][26] ),
    .A1(\w[31][26] ),
    .A2(\w[25][26] ),
    .A3(\w[29][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05859_));
 sky130_fd_sc_hd__mux4_2 _10203_ (.A0(\w[3][26] ),
    .A1(\w[7][26] ),
    .A2(\w[1][26] ),
    .A3(\w[5][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05860_));
 sky130_fd_sc_hd__mux4_2 _10204_ (.A0(\w[11][26] ),
    .A1(\w[15][26] ),
    .A2(\w[9][26] ),
    .A3(\w[13][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05861_));
 sky130_fd_sc_hd__mux4_2 _10205_ (.A0(_05858_),
    .A1(_05859_),
    .A2(_05860_),
    .A3(_05861_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05862_));
 sky130_fd_sc_hd__mux4_2 _10206_ (.A0(\w[51][26] ),
    .A1(\w[55][26] ),
    .A2(\w[49][26] ),
    .A3(\w[53][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05863_));
 sky130_fd_sc_hd__mux4_2 _10207_ (.A0(\w[59][26] ),
    .A1(\w[63][26] ),
    .A2(\w[57][26] ),
    .A3(\w[61][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05864_));
 sky130_fd_sc_hd__mux4_2 _10208_ (.A0(\w[35][26] ),
    .A1(\w[39][26] ),
    .A2(\w[33][26] ),
    .A3(\w[37][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05865_));
 sky130_fd_sc_hd__mux4_2 _10209_ (.A0(\w[43][26] ),
    .A1(\w[47][26] ),
    .A2(\w[41][26] ),
    .A3(\w[45][26] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05866_));
 sky130_fd_sc_hd__mux4_2 _10210_ (.A0(_05863_),
    .A1(_05864_),
    .A2(_05865_),
    .A3(_05866_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05867_));
 sky130_fd_sc_hd__mux2i_1 _10211_ (.A0(_05862_),
    .A1(_05867_),
    .S(_05472_),
    .Y(_05868_));
 sky130_fd_sc_hd__nand2_1 _10212_ (.A(reset_hash),
    .B(\w[1][26] ),
    .Y(_05869_));
 sky130_fd_sc_hd__o21ai_0 _10213_ (.A1(_05482_),
    .A2(_05868_),
    .B1(_05869_),
    .Y(_00050_));
 sky130_fd_sc_hd__mux4_2 _10214_ (.A0(\w[19][27] ),
    .A1(\w[23][27] ),
    .A2(\w[17][27] ),
    .A3(\w[21][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05870_));
 sky130_fd_sc_hd__mux4_2 _10215_ (.A0(\w[27][27] ),
    .A1(\w[31][27] ),
    .A2(\w[25][27] ),
    .A3(\w[29][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05871_));
 sky130_fd_sc_hd__mux4_2 _10216_ (.A0(\w[3][27] ),
    .A1(\w[7][27] ),
    .A2(\w[1][27] ),
    .A3(\w[5][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05872_));
 sky130_fd_sc_hd__mux4_2 _10217_ (.A0(\w[11][27] ),
    .A1(\w[15][27] ),
    .A2(\w[9][27] ),
    .A3(\w[13][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05873_));
 sky130_fd_sc_hd__mux4_2 _10218_ (.A0(_05870_),
    .A1(_05871_),
    .A2(_05872_),
    .A3(_05873_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05874_));
 sky130_fd_sc_hd__mux4_2 _10219_ (.A0(\w[51][27] ),
    .A1(\w[55][27] ),
    .A2(\w[49][27] ),
    .A3(\w[53][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05875_));
 sky130_fd_sc_hd__mux4_2 _10220_ (.A0(\w[59][27] ),
    .A1(\w[63][27] ),
    .A2(\w[57][27] ),
    .A3(\w[61][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05876_));
 sky130_fd_sc_hd__mux4_2 _10221_ (.A0(\w[35][27] ),
    .A1(\w[39][27] ),
    .A2(\w[33][27] ),
    .A3(\w[37][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05877_));
 sky130_fd_sc_hd__mux4_2 _10222_ (.A0(\w[43][27] ),
    .A1(\w[47][27] ),
    .A2(\w[41][27] ),
    .A3(\w[45][27] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05878_));
 sky130_fd_sc_hd__mux4_2 _10223_ (.A0(_05875_),
    .A1(_05876_),
    .A2(_05877_),
    .A3(_05878_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05879_));
 sky130_fd_sc_hd__mux2i_1 _10224_ (.A0(_05874_),
    .A1(_05879_),
    .S(_05472_),
    .Y(_05880_));
 sky130_fd_sc_hd__nand2_1 _10225_ (.A(reset_hash),
    .B(\w[1][27] ),
    .Y(_05881_));
 sky130_fd_sc_hd__o21ai_0 _10226_ (.A1(_05482_),
    .A2(_05880_),
    .B1(_05881_),
    .Y(_00051_));
 sky130_fd_sc_hd__mux4_2 _10227_ (.A0(\w[19][28] ),
    .A1(\w[23][28] ),
    .A2(\w[17][28] ),
    .A3(\w[21][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05882_));
 sky130_fd_sc_hd__mux4_2 _10228_ (.A0(\w[27][28] ),
    .A1(\w[31][28] ),
    .A2(\w[25][28] ),
    .A3(\w[29][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05883_));
 sky130_fd_sc_hd__mux4_2 _10229_ (.A0(\w[3][28] ),
    .A1(\w[7][28] ),
    .A2(\w[1][28] ),
    .A3(\w[5][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05884_));
 sky130_fd_sc_hd__mux4_2 _10230_ (.A0(\w[11][28] ),
    .A1(\w[15][28] ),
    .A2(\w[9][28] ),
    .A3(\w[13][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05885_));
 sky130_fd_sc_hd__mux4_2 _10231_ (.A0(_05882_),
    .A1(_05883_),
    .A2(_05884_),
    .A3(_05885_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05886_));
 sky130_fd_sc_hd__mux4_2 _10232_ (.A0(\w[51][28] ),
    .A1(\w[55][28] ),
    .A2(\w[49][28] ),
    .A3(\w[53][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05887_));
 sky130_fd_sc_hd__mux4_2 _10233_ (.A0(\w[59][28] ),
    .A1(\w[63][28] ),
    .A2(\w[57][28] ),
    .A3(\w[61][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05888_));
 sky130_fd_sc_hd__mux4_2 _10234_ (.A0(\w[35][28] ),
    .A1(\w[39][28] ),
    .A2(\w[33][28] ),
    .A3(\w[37][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05889_));
 sky130_fd_sc_hd__mux4_2 _10235_ (.A0(\w[43][28] ),
    .A1(\w[47][28] ),
    .A2(\w[41][28] ),
    .A3(\w[45][28] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05890_));
 sky130_fd_sc_hd__mux4_2 _10236_ (.A0(_05887_),
    .A1(_05888_),
    .A2(_05889_),
    .A3(_05890_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05891_));
 sky130_fd_sc_hd__mux2i_1 _10237_ (.A0(_05886_),
    .A1(_05891_),
    .S(_05472_),
    .Y(_05892_));
 sky130_fd_sc_hd__nand2_1 _10238_ (.A(reset_hash),
    .B(\w[1][28] ),
    .Y(_05893_));
 sky130_fd_sc_hd__o21ai_0 _10239_ (.A1(_05482_),
    .A2(_05892_),
    .B1(_05893_),
    .Y(_00052_));
 sky130_fd_sc_hd__mux4_2 _10240_ (.A0(\w[19][29] ),
    .A1(\w[23][29] ),
    .A2(\w[17][29] ),
    .A3(\w[21][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05894_));
 sky130_fd_sc_hd__mux4_2 _10241_ (.A0(\w[27][29] ),
    .A1(\w[31][29] ),
    .A2(\w[25][29] ),
    .A3(\w[29][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05895_));
 sky130_fd_sc_hd__mux4_2 _10242_ (.A0(\w[3][29] ),
    .A1(\w[7][29] ),
    .A2(\w[1][29] ),
    .A3(\w[5][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05896_));
 sky130_fd_sc_hd__mux4_2 _10243_ (.A0(\w[11][29] ),
    .A1(\w[15][29] ),
    .A2(\w[9][29] ),
    .A3(\w[13][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05897_));
 sky130_fd_sc_hd__mux4_2 _10244_ (.A0(_05894_),
    .A1(_05895_),
    .A2(_05896_),
    .A3(_05897_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05898_));
 sky130_fd_sc_hd__mux4_2 _10245_ (.A0(\w[51][29] ),
    .A1(\w[55][29] ),
    .A2(\w[49][29] ),
    .A3(\w[53][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05899_));
 sky130_fd_sc_hd__mux4_2 _10246_ (.A0(\w[59][29] ),
    .A1(\w[63][29] ),
    .A2(\w[57][29] ),
    .A3(\w[61][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05900_));
 sky130_fd_sc_hd__mux4_2 _10247_ (.A0(\w[35][29] ),
    .A1(\w[39][29] ),
    .A2(\w[33][29] ),
    .A3(\w[37][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05901_));
 sky130_fd_sc_hd__mux4_2 _10248_ (.A0(\w[43][29] ),
    .A1(\w[47][29] ),
    .A2(\w[41][29] ),
    .A3(\w[45][29] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05902_));
 sky130_fd_sc_hd__mux4_2 _10249_ (.A0(_05899_),
    .A1(_05900_),
    .A2(_05901_),
    .A3(_05902_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05903_));
 sky130_fd_sc_hd__mux2i_1 _10250_ (.A0(_05898_),
    .A1(_05903_),
    .S(_05472_),
    .Y(_05904_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(reset_hash),
    .B(\w[1][29] ),
    .Y(_05905_));
 sky130_fd_sc_hd__o21ai_0 _10252_ (.A1(_05482_),
    .A2(_05904_),
    .B1(_05905_),
    .Y(_00053_));
 sky130_fd_sc_hd__mux4_2 _10253_ (.A0(\w[19][30] ),
    .A1(\w[23][30] ),
    .A2(\w[17][30] ),
    .A3(\w[21][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05906_));
 sky130_fd_sc_hd__mux4_2 _10254_ (.A0(\w[27][30] ),
    .A1(\w[31][30] ),
    .A2(\w[25][30] ),
    .A3(\w[29][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05907_));
 sky130_fd_sc_hd__mux4_2 _10255_ (.A0(\w[3][30] ),
    .A1(\w[7][30] ),
    .A2(\w[1][30] ),
    .A3(\w[5][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05908_));
 sky130_fd_sc_hd__mux4_2 _10256_ (.A0(\w[11][30] ),
    .A1(\w[15][30] ),
    .A2(\w[9][30] ),
    .A3(\w[13][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05909_));
 sky130_fd_sc_hd__mux4_2 _10257_ (.A0(_05906_),
    .A1(_05907_),
    .A2(_05908_),
    .A3(_05909_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05910_));
 sky130_fd_sc_hd__mux4_2 _10258_ (.A0(\w[51][30] ),
    .A1(\w[55][30] ),
    .A2(\w[49][30] ),
    .A3(\w[53][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05911_));
 sky130_fd_sc_hd__mux4_2 _10259_ (.A0(\w[59][30] ),
    .A1(\w[63][30] ),
    .A2(\w[57][30] ),
    .A3(\w[61][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05912_));
 sky130_fd_sc_hd__mux4_2 _10260_ (.A0(\w[35][30] ),
    .A1(\w[39][30] ),
    .A2(\w[33][30] ),
    .A3(\w[37][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05913_));
 sky130_fd_sc_hd__mux4_2 _10261_ (.A0(\w[43][30] ),
    .A1(\w[47][30] ),
    .A2(\w[41][30] ),
    .A3(\w[45][30] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05914_));
 sky130_fd_sc_hd__mux4_2 _10262_ (.A0(_05911_),
    .A1(_05912_),
    .A2(_05913_),
    .A3(_05914_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05915_));
 sky130_fd_sc_hd__mux2i_1 _10263_ (.A0(_05910_),
    .A1(_05915_),
    .S(_05472_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_1 _10264_ (.A(reset_hash),
    .B(\w[1][30] ),
    .Y(_05917_));
 sky130_fd_sc_hd__o21ai_0 _10265_ (.A1(_05482_),
    .A2(_05916_),
    .B1(_05917_),
    .Y(_00055_));
 sky130_fd_sc_hd__mux4_2 _10266_ (.A0(\w[19][31] ),
    .A1(\w[23][31] ),
    .A2(\w[17][31] ),
    .A3(\w[21][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05918_));
 sky130_fd_sc_hd__mux4_2 _10267_ (.A0(\w[27][31] ),
    .A1(\w[31][31] ),
    .A2(\w[25][31] ),
    .A3(\w[29][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05919_));
 sky130_fd_sc_hd__mux4_2 _10268_ (.A0(\w[3][31] ),
    .A1(\w[7][31] ),
    .A2(\w[1][31] ),
    .A3(\w[5][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05920_));
 sky130_fd_sc_hd__mux4_2 _10269_ (.A0(\w[11][31] ),
    .A1(\w[15][31] ),
    .A2(\w[9][31] ),
    .A3(\w[13][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05921_));
 sky130_fd_sc_hd__mux4_2 _10270_ (.A0(_05918_),
    .A1(_05919_),
    .A2(_05920_),
    .A3(_05921_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05922_));
 sky130_fd_sc_hd__mux4_2 _10271_ (.A0(\w[51][31] ),
    .A1(\w[55][31] ),
    .A2(\w[49][31] ),
    .A3(\w[53][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05923_));
 sky130_fd_sc_hd__mux4_2 _10272_ (.A0(\w[59][31] ),
    .A1(\w[63][31] ),
    .A2(\w[57][31] ),
    .A3(\w[61][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05924_));
 sky130_fd_sc_hd__mux4_2 _10273_ (.A0(\w[35][31] ),
    .A1(\w[39][31] ),
    .A2(\w[33][31] ),
    .A3(\w[37][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05925_));
 sky130_fd_sc_hd__mux4_2 _10274_ (.A0(\w[43][31] ),
    .A1(\w[47][31] ),
    .A2(\w[41][31] ),
    .A3(\w[45][31] ),
    .S0(_00657_),
    .S1(\count_hash2[1] ),
    .X(_05926_));
 sky130_fd_sc_hd__mux4_2 _10275_ (.A0(_05923_),
    .A1(_05924_),
    .A2(_05925_),
    .A3(_05926_),
    .S0(_05458_),
    .S1(_05461_),
    .X(_05927_));
 sky130_fd_sc_hd__mux2i_1 _10276_ (.A0(_05922_),
    .A1(_05927_),
    .S(_05472_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _10277_ (.A(reset_hash),
    .B(\w[1][31] ),
    .Y(_05929_));
 sky130_fd_sc_hd__o21ai_0 _10278_ (.A1(_05482_),
    .A2(_05928_),
    .B1(_05929_),
    .Y(_00056_));
 sky130_fd_sc_hd__mux4_2 _10286_ (.A0(\w[18][0] ),
    .A1(\w[16][0] ),
    .A2(\w[22][0] ),
    .A3(\w[20][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05937_));
 sky130_fd_sc_hd__mux4_2 _10291_ (.A0(\w[26][0] ),
    .A1(\w[24][0] ),
    .A2(\w[30][0] ),
    .A3(\w[28][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05942_));
 sky130_fd_sc_hd__mux4_2 _10294_ (.A0(\w[2][0] ),
    .A1(\w[0][0] ),
    .A2(\w[6][0] ),
    .A3(\w[4][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05945_));
 sky130_fd_sc_hd__mux4_2 _10299_ (.A0(\w[10][0] ),
    .A1(\w[8][0] ),
    .A2(\w[14][0] ),
    .A3(\w[12][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05950_));
 sky130_fd_sc_hd__nor2b_1 _10300_ (.A(_09366_),
    .B_N(\count_hash1[3] ),
    .Y(_05951_));
 sky130_fd_sc_hd__nor2b_1 _10301_ (.A(\count_hash1[3] ),
    .B_N(_09366_),
    .Y(_05952_));
 sky130_fd_sc_hd__or2_4 _10302_ (.A(_05951_),
    .B(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__inv_1 _10305_ (.A(\count_hash1[4] ),
    .Y(_05956_));
 sky130_fd_sc_hd__nand3_2 _10306_ (.A(\count_hash1[3] ),
    .B(\count_hash1[2] ),
    .C(\count_hash1[1] ),
    .Y(_05957_));
 sky130_fd_sc_hd__xnor2_2 _10307_ (.A(_05956_),
    .B(_05957_),
    .Y(_05958_));
 sky130_fd_sc_hd__mux4_2 _10310_ (.A0(_05937_),
    .A1(_05942_),
    .A2(_05945_),
    .A3(_05950_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_05961_));
 sky130_fd_sc_hd__mux4_2 _10313_ (.A0(\w[50][0] ),
    .A1(\w[48][0] ),
    .A2(\w[54][0] ),
    .A3(\w[52][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05964_));
 sky130_fd_sc_hd__mux4_2 _10316_ (.A0(\w[58][0] ),
    .A1(\w[56][0] ),
    .A2(\w[62][0] ),
    .A3(\w[60][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05967_));
 sky130_fd_sc_hd__mux4_2 _10319_ (.A0(\w[34][0] ),
    .A1(\w[32][0] ),
    .A2(\w[38][0] ),
    .A3(\w[36][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05970_));
 sky130_fd_sc_hd__mux4_2 _10322_ (.A0(\w[42][0] ),
    .A1(\w[40][0] ),
    .A2(\w[46][0] ),
    .A3(\w[44][0] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05973_));
 sky130_fd_sc_hd__mux4_2 _10325_ (.A0(_05964_),
    .A1(_05967_),
    .A2(_05970_),
    .A3(_05973_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_05976_));
 sky130_fd_sc_hd__nand3_1 _10326_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(_09366_),
    .Y(_05977_));
 sky130_fd_sc_hd__xnor2_2 _10327_ (.A(\count_hash1[5] ),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__mux2i_1 _10331_ (.A0(_05961_),
    .A1(_05976_),
    .S(_05978_),
    .Y(_05982_));
 sky130_fd_sc_hd__nand2_1 _10332_ (.A(reset_hash),
    .B(\w[0][0] ),
    .Y(_05983_));
 sky130_fd_sc_hd__o21ai_0 _10333_ (.A1(_05482_),
    .A2(_05982_),
    .B1(_05983_),
    .Y(_00000_));
 sky130_fd_sc_hd__mux4_2 _10334_ (.A0(\w[18][1] ),
    .A1(\w[16][1] ),
    .A2(\w[22][1] ),
    .A3(\w[20][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05984_));
 sky130_fd_sc_hd__mux4_2 _10335_ (.A0(\w[26][1] ),
    .A1(\w[24][1] ),
    .A2(\w[30][1] ),
    .A3(\w[28][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05985_));
 sky130_fd_sc_hd__mux4_2 _10336_ (.A0(\w[2][1] ),
    .A1(\w[0][1] ),
    .A2(\w[6][1] ),
    .A3(\w[4][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05986_));
 sky130_fd_sc_hd__mux4_2 _10337_ (.A0(\w[10][1] ),
    .A1(\w[8][1] ),
    .A2(\w[14][1] ),
    .A3(\w[12][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05987_));
 sky130_fd_sc_hd__mux4_2 _10338_ (.A0(_05984_),
    .A1(_05985_),
    .A2(_05986_),
    .A3(_05987_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_05988_));
 sky130_fd_sc_hd__mux4_2 _10340_ (.A0(\w[50][1] ),
    .A1(\w[48][1] ),
    .A2(\w[54][1] ),
    .A3(\w[52][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05990_));
 sky130_fd_sc_hd__mux4_2 _10341_ (.A0(\w[58][1] ),
    .A1(\w[56][1] ),
    .A2(\w[62][1] ),
    .A3(\w[60][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05991_));
 sky130_fd_sc_hd__mux4_2 _10342_ (.A0(\w[34][1] ),
    .A1(\w[32][1] ),
    .A2(\w[38][1] ),
    .A3(\w[36][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05992_));
 sky130_fd_sc_hd__mux4_2 _10343_ (.A0(\w[42][1] ),
    .A1(\w[40][1] ),
    .A2(\w[46][1] ),
    .A3(\w[44][1] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05993_));
 sky130_fd_sc_hd__mux4_2 _10344_ (.A0(_05990_),
    .A1(_05991_),
    .A2(_05992_),
    .A3(_05993_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_05994_));
 sky130_fd_sc_hd__mux2i_1 _10345_ (.A0(_05988_),
    .A1(_05994_),
    .S(_05978_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2_1 _10346_ (.A(reset_hash),
    .B(\w[0][1] ),
    .Y(_05996_));
 sky130_fd_sc_hd__o21ai_0 _10347_ (.A1(_05482_),
    .A2(_05995_),
    .B1(_05996_),
    .Y(_00011_));
 sky130_fd_sc_hd__mux4_2 _10348_ (.A0(\w[18][2] ),
    .A1(\w[16][2] ),
    .A2(\w[22][2] ),
    .A3(\w[20][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05997_));
 sky130_fd_sc_hd__mux4_2 _10349_ (.A0(\w[26][2] ),
    .A1(\w[24][2] ),
    .A2(\w[30][2] ),
    .A3(\w[28][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_05998_));
 sky130_fd_sc_hd__mux4_2 _10351_ (.A0(\w[2][2] ),
    .A1(\w[0][2] ),
    .A2(\w[6][2] ),
    .A3(\w[4][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06000_));
 sky130_fd_sc_hd__mux4_2 _10352_ (.A0(\w[10][2] ),
    .A1(\w[8][2] ),
    .A2(\w[14][2] ),
    .A3(\w[12][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06001_));
 sky130_fd_sc_hd__mux4_2 _10353_ (.A0(_05997_),
    .A1(_05998_),
    .A2(_06000_),
    .A3(_06001_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06002_));
 sky130_fd_sc_hd__mux4_2 _10354_ (.A0(\w[50][2] ),
    .A1(\w[48][2] ),
    .A2(\w[54][2] ),
    .A3(\w[52][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06003_));
 sky130_fd_sc_hd__mux4_2 _10355_ (.A0(\w[58][2] ),
    .A1(\w[56][2] ),
    .A2(\w[62][2] ),
    .A3(\w[60][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06004_));
 sky130_fd_sc_hd__mux4_2 _10356_ (.A0(\w[34][2] ),
    .A1(\w[32][2] ),
    .A2(\w[38][2] ),
    .A3(\w[36][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06005_));
 sky130_fd_sc_hd__mux4_2 _10357_ (.A0(\w[42][2] ),
    .A1(\w[40][2] ),
    .A2(\w[46][2] ),
    .A3(\w[44][2] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06006_));
 sky130_fd_sc_hd__mux4_2 _10358_ (.A0(_06003_),
    .A1(_06004_),
    .A2(_06005_),
    .A3(_06006_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06007_));
 sky130_fd_sc_hd__mux2i_1 _10359_ (.A0(_06002_),
    .A1(_06007_),
    .S(_05978_),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_1 _10361_ (.A(reset_hash),
    .B(\w[0][2] ),
    .Y(_06010_));
 sky130_fd_sc_hd__o21ai_0 _10362_ (.A1(_05482_),
    .A2(_06008_),
    .B1(_06010_),
    .Y(_00022_));
 sky130_fd_sc_hd__mux4_2 _10363_ (.A0(\w[18][3] ),
    .A1(\w[16][3] ),
    .A2(\w[22][3] ),
    .A3(\w[20][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06011_));
 sky130_fd_sc_hd__mux4_2 _10364_ (.A0(\w[26][3] ),
    .A1(\w[24][3] ),
    .A2(\w[30][3] ),
    .A3(\w[28][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06012_));
 sky130_fd_sc_hd__mux4_2 _10366_ (.A0(\w[2][3] ),
    .A1(\w[0][3] ),
    .A2(\w[6][3] ),
    .A3(\w[4][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06014_));
 sky130_fd_sc_hd__mux4_2 _10367_ (.A0(\w[10][3] ),
    .A1(\w[8][3] ),
    .A2(\w[14][3] ),
    .A3(\w[12][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06015_));
 sky130_fd_sc_hd__mux4_2 _10368_ (.A0(_06011_),
    .A1(_06012_),
    .A2(_06014_),
    .A3(_06015_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06016_));
 sky130_fd_sc_hd__mux4_2 _10369_ (.A0(\w[50][3] ),
    .A1(\w[48][3] ),
    .A2(\w[54][3] ),
    .A3(\w[52][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06017_));
 sky130_fd_sc_hd__mux4_2 _10370_ (.A0(\w[58][3] ),
    .A1(\w[56][3] ),
    .A2(\w[62][3] ),
    .A3(\w[60][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06018_));
 sky130_fd_sc_hd__mux4_2 _10371_ (.A0(\w[34][3] ),
    .A1(\w[32][3] ),
    .A2(\w[38][3] ),
    .A3(\w[36][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06019_));
 sky130_fd_sc_hd__mux4_2 _10372_ (.A0(\w[42][3] ),
    .A1(\w[40][3] ),
    .A2(\w[46][3] ),
    .A3(\w[44][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06020_));
 sky130_fd_sc_hd__mux4_2 _10373_ (.A0(_06017_),
    .A1(_06018_),
    .A2(_06019_),
    .A3(_06020_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06021_));
 sky130_fd_sc_hd__mux2i_1 _10374_ (.A0(_06016_),
    .A1(_06021_),
    .S(_05978_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand2_1 _10375_ (.A(reset_hash),
    .B(\w[0][3] ),
    .Y(_06023_));
 sky130_fd_sc_hd__o21ai_0 _10376_ (.A1(_05482_),
    .A2(_06022_),
    .B1(_06023_),
    .Y(_00025_));
 sky130_fd_sc_hd__mux4_2 _10378_ (.A0(\w[18][4] ),
    .A1(\w[16][4] ),
    .A2(\w[22][4] ),
    .A3(\w[20][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06025_));
 sky130_fd_sc_hd__mux4_2 _10379_ (.A0(\w[26][4] ),
    .A1(\w[24][4] ),
    .A2(\w[30][4] ),
    .A3(\w[28][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06026_));
 sky130_fd_sc_hd__mux4_2 _10380_ (.A0(\w[2][4] ),
    .A1(\w[0][4] ),
    .A2(\w[6][4] ),
    .A3(\w[4][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06027_));
 sky130_fd_sc_hd__mux4_2 _10381_ (.A0(\w[10][4] ),
    .A1(\w[8][4] ),
    .A2(\w[14][4] ),
    .A3(\w[12][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06028_));
 sky130_fd_sc_hd__mux4_2 _10382_ (.A0(_06025_),
    .A1(_06026_),
    .A2(_06027_),
    .A3(_06028_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06029_));
 sky130_fd_sc_hd__mux4_2 _10383_ (.A0(\w[50][4] ),
    .A1(\w[48][4] ),
    .A2(\w[54][4] ),
    .A3(\w[52][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06030_));
 sky130_fd_sc_hd__mux4_2 _10385_ (.A0(\w[58][4] ),
    .A1(\w[56][4] ),
    .A2(\w[62][4] ),
    .A3(\w[60][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06032_));
 sky130_fd_sc_hd__mux4_2 _10386_ (.A0(\w[34][4] ),
    .A1(\w[32][4] ),
    .A2(\w[38][4] ),
    .A3(\w[36][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06033_));
 sky130_fd_sc_hd__mux4_2 _10387_ (.A0(\w[42][4] ),
    .A1(\w[40][4] ),
    .A2(\w[46][4] ),
    .A3(\w[44][4] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06034_));
 sky130_fd_sc_hd__mux4_2 _10389_ (.A0(_06030_),
    .A1(_06032_),
    .A2(_06033_),
    .A3(_06034_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06036_));
 sky130_fd_sc_hd__mux2i_1 _10390_ (.A0(_06029_),
    .A1(_06036_),
    .S(_05978_),
    .Y(_06037_));
 sky130_fd_sc_hd__nand2_1 _10391_ (.A(reset_hash),
    .B(\w[0][4] ),
    .Y(_06038_));
 sky130_fd_sc_hd__o21ai_0 _10392_ (.A1(_05482_),
    .A2(_06037_),
    .B1(_06038_),
    .Y(_00026_));
 sky130_fd_sc_hd__mux4_2 _10394_ (.A0(\w[18][5] ),
    .A1(\w[16][5] ),
    .A2(\w[22][5] ),
    .A3(\w[20][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06040_));
 sky130_fd_sc_hd__mux4_2 _10395_ (.A0(\w[26][5] ),
    .A1(\w[24][5] ),
    .A2(\w[30][5] ),
    .A3(\w[28][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06041_));
 sky130_fd_sc_hd__mux4_2 _10396_ (.A0(\w[2][5] ),
    .A1(\w[0][5] ),
    .A2(\w[6][5] ),
    .A3(\w[4][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06042_));
 sky130_fd_sc_hd__mux4_2 _10397_ (.A0(\w[10][5] ),
    .A1(\w[8][5] ),
    .A2(\w[14][5] ),
    .A3(\w[12][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06043_));
 sky130_fd_sc_hd__mux4_2 _10398_ (.A0(_06040_),
    .A1(_06041_),
    .A2(_06042_),
    .A3(_06043_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06044_));
 sky130_fd_sc_hd__mux4_2 _10399_ (.A0(\w[50][5] ),
    .A1(\w[48][5] ),
    .A2(\w[54][5] ),
    .A3(\w[52][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06045_));
 sky130_fd_sc_hd__mux4_2 _10401_ (.A0(\w[58][5] ),
    .A1(\w[56][5] ),
    .A2(\w[62][5] ),
    .A3(\w[60][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06047_));
 sky130_fd_sc_hd__mux4_2 _10402_ (.A0(\w[34][5] ),
    .A1(\w[32][5] ),
    .A2(\w[38][5] ),
    .A3(\w[36][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06048_));
 sky130_fd_sc_hd__mux4_2 _10403_ (.A0(\w[42][5] ),
    .A1(\w[40][5] ),
    .A2(\w[46][5] ),
    .A3(\w[44][5] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06049_));
 sky130_fd_sc_hd__mux4_2 _10404_ (.A0(_06045_),
    .A1(_06047_),
    .A2(_06048_),
    .A3(_06049_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06050_));
 sky130_fd_sc_hd__mux2i_1 _10405_ (.A0(_06044_),
    .A1(_06050_),
    .S(_05978_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand2_1 _10406_ (.A(reset_hash),
    .B(\w[0][5] ),
    .Y(_06052_));
 sky130_fd_sc_hd__o21ai_0 _10407_ (.A1(_05482_),
    .A2(_06051_),
    .B1(_06052_),
    .Y(_00027_));
 sky130_fd_sc_hd__mux4_2 _10408_ (.A0(\w[18][6] ),
    .A1(\w[16][6] ),
    .A2(\w[22][6] ),
    .A3(\w[20][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06053_));
 sky130_fd_sc_hd__mux4_2 _10410_ (.A0(\w[26][6] ),
    .A1(\w[24][6] ),
    .A2(\w[30][6] ),
    .A3(\w[28][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06055_));
 sky130_fd_sc_hd__mux4_2 _10411_ (.A0(\w[2][6] ),
    .A1(\w[0][6] ),
    .A2(\w[6][6] ),
    .A3(\w[4][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06056_));
 sky130_fd_sc_hd__mux4_2 _10412_ (.A0(\w[10][6] ),
    .A1(\w[8][6] ),
    .A2(\w[14][6] ),
    .A3(\w[12][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06057_));
 sky130_fd_sc_hd__mux4_2 _10414_ (.A0(_06053_),
    .A1(_06055_),
    .A2(_06056_),
    .A3(_06057_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06059_));
 sky130_fd_sc_hd__mux4_2 _10415_ (.A0(\w[50][6] ),
    .A1(\w[48][6] ),
    .A2(\w[54][6] ),
    .A3(\w[52][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06060_));
 sky130_fd_sc_hd__mux4_2 _10416_ (.A0(\w[58][6] ),
    .A1(\w[56][6] ),
    .A2(\w[62][6] ),
    .A3(\w[60][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06061_));
 sky130_fd_sc_hd__mux4_2 _10417_ (.A0(\w[34][6] ),
    .A1(\w[32][6] ),
    .A2(\w[38][6] ),
    .A3(\w[36][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06062_));
 sky130_fd_sc_hd__mux4_2 _10419_ (.A0(\w[42][6] ),
    .A1(\w[40][6] ),
    .A2(\w[46][6] ),
    .A3(\w[44][6] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06064_));
 sky130_fd_sc_hd__mux4_2 _10421_ (.A0(_06060_),
    .A1(_06061_),
    .A2(_06062_),
    .A3(_06064_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06066_));
 sky130_fd_sc_hd__mux2i_1 _10423_ (.A0(_06059_),
    .A1(_06066_),
    .S(_05978_),
    .Y(_06068_));
 sky130_fd_sc_hd__nand2_1 _10424_ (.A(reset_hash),
    .B(\w[0][6] ),
    .Y(_06069_));
 sky130_fd_sc_hd__o21ai_0 _10425_ (.A1(_05482_),
    .A2(_06068_),
    .B1(_06069_),
    .Y(_00028_));
 sky130_fd_sc_hd__mux4_2 _10426_ (.A0(\w[18][7] ),
    .A1(\w[16][7] ),
    .A2(\w[22][7] ),
    .A3(\w[20][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06070_));
 sky130_fd_sc_hd__mux4_2 _10428_ (.A0(\w[26][7] ),
    .A1(\w[24][7] ),
    .A2(\w[30][7] ),
    .A3(\w[28][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06072_));
 sky130_fd_sc_hd__mux4_2 _10429_ (.A0(\w[2][7] ),
    .A1(\w[0][7] ),
    .A2(\w[6][7] ),
    .A3(\w[4][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06073_));
 sky130_fd_sc_hd__mux4_2 _10430_ (.A0(\w[10][7] ),
    .A1(\w[8][7] ),
    .A2(\w[14][7] ),
    .A3(\w[12][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06074_));
 sky130_fd_sc_hd__mux4_2 _10431_ (.A0(_06070_),
    .A1(_06072_),
    .A2(_06073_),
    .A3(_06074_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06075_));
 sky130_fd_sc_hd__mux4_2 _10432_ (.A0(\w[50][7] ),
    .A1(\w[48][7] ),
    .A2(\w[54][7] ),
    .A3(\w[52][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06076_));
 sky130_fd_sc_hd__mux4_2 _10433_ (.A0(\w[58][7] ),
    .A1(\w[56][7] ),
    .A2(\w[62][7] ),
    .A3(\w[60][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06077_));
 sky130_fd_sc_hd__mux4_2 _10434_ (.A0(\w[34][7] ),
    .A1(\w[32][7] ),
    .A2(\w[38][7] ),
    .A3(\w[36][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06078_));
 sky130_fd_sc_hd__mux4_2 _10436_ (.A0(\w[42][7] ),
    .A1(\w[40][7] ),
    .A2(\w[46][7] ),
    .A3(\w[44][7] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06080_));
 sky130_fd_sc_hd__mux4_2 _10437_ (.A0(_06076_),
    .A1(_06077_),
    .A2(_06078_),
    .A3(_06080_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06081_));
 sky130_fd_sc_hd__mux2i_1 _10438_ (.A0(_06075_),
    .A1(_06081_),
    .S(_05978_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand2_1 _10439_ (.A(reset_hash),
    .B(\w[0][7] ),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_0 _10440_ (.A1(_05482_),
    .A2(_06082_),
    .B1(_06083_),
    .Y(_00029_));
 sky130_fd_sc_hd__mux4_2 _10441_ (.A0(\w[18][8] ),
    .A1(\w[16][8] ),
    .A2(\w[22][8] ),
    .A3(\w[20][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06084_));
 sky130_fd_sc_hd__mux4_2 _10442_ (.A0(\w[26][8] ),
    .A1(\w[24][8] ),
    .A2(\w[30][8] ),
    .A3(\w[28][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06085_));
 sky130_fd_sc_hd__mux4_2 _10443_ (.A0(\w[2][8] ),
    .A1(\w[0][8] ),
    .A2(\w[6][8] ),
    .A3(\w[4][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06086_));
 sky130_fd_sc_hd__mux4_2 _10445_ (.A0(\w[10][8] ),
    .A1(\w[8][8] ),
    .A2(\w[14][8] ),
    .A3(\w[12][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06088_));
 sky130_fd_sc_hd__mux4_2 _10447_ (.A0(_06084_),
    .A1(_06085_),
    .A2(_06086_),
    .A3(_06088_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06090_));
 sky130_fd_sc_hd__mux4_2 _10448_ (.A0(\w[50][8] ),
    .A1(\w[48][8] ),
    .A2(\w[54][8] ),
    .A3(\w[52][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06091_));
 sky130_fd_sc_hd__mux4_2 _10449_ (.A0(\w[58][8] ),
    .A1(\w[56][8] ),
    .A2(\w[62][8] ),
    .A3(\w[60][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06092_));
 sky130_fd_sc_hd__mux4_2 _10451_ (.A0(\w[34][8] ),
    .A1(\w[32][8] ),
    .A2(\w[38][8] ),
    .A3(\w[36][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06094_));
 sky130_fd_sc_hd__mux4_2 _10452_ (.A0(\w[42][8] ),
    .A1(\w[40][8] ),
    .A2(\w[46][8] ),
    .A3(\w[44][8] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06095_));
 sky130_fd_sc_hd__mux4_2 _10453_ (.A0(_06091_),
    .A1(_06092_),
    .A2(_06094_),
    .A3(_06095_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06096_));
 sky130_fd_sc_hd__mux2i_1 _10454_ (.A0(_06090_),
    .A1(_06096_),
    .S(_05978_),
    .Y(_06097_));
 sky130_fd_sc_hd__nand2_1 _10455_ (.A(reset_hash),
    .B(\w[0][8] ),
    .Y(_06098_));
 sky130_fd_sc_hd__o21ai_0 _10456_ (.A1(_05482_),
    .A2(_06097_),
    .B1(_06098_),
    .Y(_00030_));
 sky130_fd_sc_hd__mux4_2 _10457_ (.A0(\w[18][9] ),
    .A1(\w[16][9] ),
    .A2(\w[22][9] ),
    .A3(\w[20][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06099_));
 sky130_fd_sc_hd__mux4_2 _10458_ (.A0(\w[26][9] ),
    .A1(\w[24][9] ),
    .A2(\w[30][9] ),
    .A3(\w[28][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06100_));
 sky130_fd_sc_hd__mux4_2 _10459_ (.A0(\w[2][9] ),
    .A1(\w[0][9] ),
    .A2(\w[6][9] ),
    .A3(\w[4][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06101_));
 sky130_fd_sc_hd__mux4_2 _10461_ (.A0(\w[10][9] ),
    .A1(\w[8][9] ),
    .A2(\w[14][9] ),
    .A3(\w[12][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06103_));
 sky130_fd_sc_hd__mux4_2 _10462_ (.A0(_06099_),
    .A1(_06100_),
    .A2(_06101_),
    .A3(_06103_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06104_));
 sky130_fd_sc_hd__mux4_2 _10463_ (.A0(\w[50][9] ),
    .A1(\w[48][9] ),
    .A2(\w[54][9] ),
    .A3(\w[52][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06105_));
 sky130_fd_sc_hd__mux4_2 _10464_ (.A0(\w[58][9] ),
    .A1(\w[56][9] ),
    .A2(\w[62][9] ),
    .A3(\w[60][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06106_));
 sky130_fd_sc_hd__mux4_2 _10466_ (.A0(\w[34][9] ),
    .A1(\w[32][9] ),
    .A2(\w[38][9] ),
    .A3(\w[36][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06108_));
 sky130_fd_sc_hd__mux4_2 _10467_ (.A0(\w[42][9] ),
    .A1(\w[40][9] ),
    .A2(\w[46][9] ),
    .A3(\w[44][9] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06109_));
 sky130_fd_sc_hd__mux4_2 _10468_ (.A0(_06105_),
    .A1(_06106_),
    .A2(_06108_),
    .A3(_06109_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06110_));
 sky130_fd_sc_hd__mux2i_1 _10469_ (.A0(_06104_),
    .A1(_06110_),
    .S(_05978_),
    .Y(_06111_));
 sky130_fd_sc_hd__nand2_1 _10470_ (.A(reset_hash),
    .B(\w[0][9] ),
    .Y(_06112_));
 sky130_fd_sc_hd__o21ai_0 _10471_ (.A1(_05482_),
    .A2(_06111_),
    .B1(_06112_),
    .Y(_00031_));
 sky130_fd_sc_hd__mux4_2 _10473_ (.A0(\w[18][10] ),
    .A1(\w[16][10] ),
    .A2(\w[22][10] ),
    .A3(\w[20][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06114_));
 sky130_fd_sc_hd__mux4_2 _10474_ (.A0(\w[26][10] ),
    .A1(\w[24][10] ),
    .A2(\w[30][10] ),
    .A3(\w[28][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06115_));
 sky130_fd_sc_hd__mux4_2 _10475_ (.A0(\w[2][10] ),
    .A1(\w[0][10] ),
    .A2(\w[6][10] ),
    .A3(\w[4][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06116_));
 sky130_fd_sc_hd__mux4_2 _10476_ (.A0(\w[10][10] ),
    .A1(\w[8][10] ),
    .A2(\w[14][10] ),
    .A3(\w[12][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06117_));
 sky130_fd_sc_hd__mux4_2 _10477_ (.A0(_06114_),
    .A1(_06115_),
    .A2(_06116_),
    .A3(_06117_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06118_));
 sky130_fd_sc_hd__mux4_2 _10479_ (.A0(\w[50][10] ),
    .A1(\w[48][10] ),
    .A2(\w[54][10] ),
    .A3(\w[52][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06120_));
 sky130_fd_sc_hd__mux4_2 _10480_ (.A0(\w[58][10] ),
    .A1(\w[56][10] ),
    .A2(\w[62][10] ),
    .A3(\w[60][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06121_));
 sky130_fd_sc_hd__mux4_2 _10481_ (.A0(\w[34][10] ),
    .A1(\w[32][10] ),
    .A2(\w[38][10] ),
    .A3(\w[36][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06122_));
 sky130_fd_sc_hd__mux4_2 _10482_ (.A0(\w[42][10] ),
    .A1(\w[40][10] ),
    .A2(\w[46][10] ),
    .A3(\w[44][10] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06123_));
 sky130_fd_sc_hd__mux4_2 _10483_ (.A0(_06120_),
    .A1(_06121_),
    .A2(_06122_),
    .A3(_06123_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06124_));
 sky130_fd_sc_hd__mux2i_1 _10484_ (.A0(_06118_),
    .A1(_06124_),
    .S(_05978_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_1 _10485_ (.A(reset_hash),
    .B(\w[0][10] ),
    .Y(_06126_));
 sky130_fd_sc_hd__o21ai_0 _10486_ (.A1(_05482_),
    .A2(_06125_),
    .B1(_06126_),
    .Y(_00001_));
 sky130_fd_sc_hd__mux4_2 _10487_ (.A0(\w[18][11] ),
    .A1(\w[16][11] ),
    .A2(\w[22][11] ),
    .A3(\w[20][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06127_));
 sky130_fd_sc_hd__mux4_2 _10488_ (.A0(\w[26][11] ),
    .A1(\w[24][11] ),
    .A2(\w[30][11] ),
    .A3(\w[28][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06128_));
 sky130_fd_sc_hd__mux4_2 _10489_ (.A0(\w[2][11] ),
    .A1(\w[0][11] ),
    .A2(\w[6][11] ),
    .A3(\w[4][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06129_));
 sky130_fd_sc_hd__mux4_2 _10490_ (.A0(\w[10][11] ),
    .A1(\w[8][11] ),
    .A2(\w[14][11] ),
    .A3(\w[12][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06130_));
 sky130_fd_sc_hd__mux4_2 _10491_ (.A0(_06127_),
    .A1(_06128_),
    .A2(_06129_),
    .A3(_06130_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06131_));
 sky130_fd_sc_hd__mux4_2 _10493_ (.A0(\w[50][11] ),
    .A1(\w[48][11] ),
    .A2(\w[54][11] ),
    .A3(\w[52][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06133_));
 sky130_fd_sc_hd__mux4_2 _10494_ (.A0(\w[58][11] ),
    .A1(\w[56][11] ),
    .A2(\w[62][11] ),
    .A3(\w[60][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06134_));
 sky130_fd_sc_hd__mux4_2 _10495_ (.A0(\w[34][11] ),
    .A1(\w[32][11] ),
    .A2(\w[38][11] ),
    .A3(\w[36][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06135_));
 sky130_fd_sc_hd__mux4_2 _10496_ (.A0(\w[42][11] ),
    .A1(\w[40][11] ),
    .A2(\w[46][11] ),
    .A3(\w[44][11] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06136_));
 sky130_fd_sc_hd__mux4_2 _10497_ (.A0(_06133_),
    .A1(_06134_),
    .A2(_06135_),
    .A3(_06136_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06137_));
 sky130_fd_sc_hd__mux2i_1 _10498_ (.A0(_06131_),
    .A1(_06137_),
    .S(_05978_),
    .Y(_06138_));
 sky130_fd_sc_hd__nand2_1 _10499_ (.A(reset_hash),
    .B(\w[0][11] ),
    .Y(_06139_));
 sky130_fd_sc_hd__o21ai_0 _10500_ (.A1(_05482_),
    .A2(_06138_),
    .B1(_06139_),
    .Y(_00002_));
 sky130_fd_sc_hd__mux4_2 _10501_ (.A0(\w[18][12] ),
    .A1(\w[16][12] ),
    .A2(\w[22][12] ),
    .A3(\w[20][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06140_));
 sky130_fd_sc_hd__mux4_2 _10502_ (.A0(\w[26][12] ),
    .A1(\w[24][12] ),
    .A2(\w[30][12] ),
    .A3(\w[28][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06141_));
 sky130_fd_sc_hd__mux4_2 _10504_ (.A0(\w[2][12] ),
    .A1(\w[0][12] ),
    .A2(\w[6][12] ),
    .A3(\w[4][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06143_));
 sky130_fd_sc_hd__mux4_2 _10505_ (.A0(\w[10][12] ),
    .A1(\w[8][12] ),
    .A2(\w[14][12] ),
    .A3(\w[12][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06144_));
 sky130_fd_sc_hd__mux4_2 _10506_ (.A0(_06140_),
    .A1(_06141_),
    .A2(_06143_),
    .A3(_06144_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06145_));
 sky130_fd_sc_hd__mux4_2 _10507_ (.A0(\w[50][12] ),
    .A1(\w[48][12] ),
    .A2(\w[54][12] ),
    .A3(\w[52][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06146_));
 sky130_fd_sc_hd__mux4_2 _10508_ (.A0(\w[58][12] ),
    .A1(\w[56][12] ),
    .A2(\w[62][12] ),
    .A3(\w[60][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06147_));
 sky130_fd_sc_hd__mux4_2 _10509_ (.A0(\w[34][12] ),
    .A1(\w[32][12] ),
    .A2(\w[38][12] ),
    .A3(\w[36][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06148_));
 sky130_fd_sc_hd__mux4_2 _10510_ (.A0(\w[42][12] ),
    .A1(\w[40][12] ),
    .A2(\w[46][12] ),
    .A3(\w[44][12] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06149_));
 sky130_fd_sc_hd__mux4_2 _10511_ (.A0(_06146_),
    .A1(_06147_),
    .A2(_06148_),
    .A3(_06149_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06150_));
 sky130_fd_sc_hd__mux2i_1 _10512_ (.A0(_06145_),
    .A1(_06150_),
    .S(_05978_),
    .Y(_06151_));
 sky130_fd_sc_hd__nand2_1 _10514_ (.A(reset_hash),
    .B(\w[0][12] ),
    .Y(_06153_));
 sky130_fd_sc_hd__o21ai_0 _10515_ (.A1(_05482_),
    .A2(_06151_),
    .B1(_06153_),
    .Y(_00003_));
 sky130_fd_sc_hd__mux4_2 _10516_ (.A0(\w[18][13] ),
    .A1(\w[16][13] ),
    .A2(\w[22][13] ),
    .A3(\w[20][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06154_));
 sky130_fd_sc_hd__mux4_2 _10517_ (.A0(\w[26][13] ),
    .A1(\w[24][13] ),
    .A2(\w[30][13] ),
    .A3(\w[28][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06155_));
 sky130_fd_sc_hd__mux4_2 _10519_ (.A0(\w[2][13] ),
    .A1(\w[0][13] ),
    .A2(\w[6][13] ),
    .A3(\w[4][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06157_));
 sky130_fd_sc_hd__mux4_2 _10520_ (.A0(\w[10][13] ),
    .A1(\w[8][13] ),
    .A2(\w[14][13] ),
    .A3(\w[12][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06158_));
 sky130_fd_sc_hd__mux4_2 _10521_ (.A0(_06154_),
    .A1(_06155_),
    .A2(_06157_),
    .A3(_06158_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06159_));
 sky130_fd_sc_hd__mux4_2 _10522_ (.A0(\w[50][13] ),
    .A1(\w[48][13] ),
    .A2(\w[54][13] ),
    .A3(\w[52][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06160_));
 sky130_fd_sc_hd__mux4_2 _10523_ (.A0(\w[58][13] ),
    .A1(\w[56][13] ),
    .A2(\w[62][13] ),
    .A3(\w[60][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06161_));
 sky130_fd_sc_hd__mux4_2 _10524_ (.A0(\w[34][13] ),
    .A1(\w[32][13] ),
    .A2(\w[38][13] ),
    .A3(\w[36][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06162_));
 sky130_fd_sc_hd__mux4_2 _10525_ (.A0(\w[42][13] ),
    .A1(\w[40][13] ),
    .A2(\w[46][13] ),
    .A3(\w[44][13] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06163_));
 sky130_fd_sc_hd__mux4_2 _10526_ (.A0(_06160_),
    .A1(_06161_),
    .A2(_06162_),
    .A3(_06163_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06164_));
 sky130_fd_sc_hd__mux2i_1 _10527_ (.A0(_06159_),
    .A1(_06164_),
    .S(_05978_),
    .Y(_06165_));
 sky130_fd_sc_hd__nand2_1 _10528_ (.A(reset_hash),
    .B(\w[0][13] ),
    .Y(_06166_));
 sky130_fd_sc_hd__o21ai_0 _10529_ (.A1(_05482_),
    .A2(_06165_),
    .B1(_06166_),
    .Y(_00004_));
 sky130_fd_sc_hd__mux4_2 _10531_ (.A0(\w[18][14] ),
    .A1(\w[16][14] ),
    .A2(\w[22][14] ),
    .A3(\w[20][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06168_));
 sky130_fd_sc_hd__mux4_2 _10532_ (.A0(\w[26][14] ),
    .A1(\w[24][14] ),
    .A2(\w[30][14] ),
    .A3(\w[28][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06169_));
 sky130_fd_sc_hd__mux4_2 _10533_ (.A0(\w[2][14] ),
    .A1(\w[0][14] ),
    .A2(\w[6][14] ),
    .A3(\w[4][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06170_));
 sky130_fd_sc_hd__mux4_2 _10534_ (.A0(\w[10][14] ),
    .A1(\w[8][14] ),
    .A2(\w[14][14] ),
    .A3(\w[12][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06171_));
 sky130_fd_sc_hd__mux4_2 _10535_ (.A0(_06168_),
    .A1(_06169_),
    .A2(_06170_),
    .A3(_06171_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06172_));
 sky130_fd_sc_hd__mux4_2 _10536_ (.A0(\w[50][14] ),
    .A1(\w[48][14] ),
    .A2(\w[54][14] ),
    .A3(\w[52][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06173_));
 sky130_fd_sc_hd__mux4_2 _10538_ (.A0(\w[58][14] ),
    .A1(\w[56][14] ),
    .A2(\w[62][14] ),
    .A3(\w[60][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06175_));
 sky130_fd_sc_hd__mux4_2 _10539_ (.A0(\w[34][14] ),
    .A1(\w[32][14] ),
    .A2(\w[38][14] ),
    .A3(\w[36][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06176_));
 sky130_fd_sc_hd__mux4_2 _10540_ (.A0(\w[42][14] ),
    .A1(\w[40][14] ),
    .A2(\w[46][14] ),
    .A3(\w[44][14] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06177_));
 sky130_fd_sc_hd__mux4_2 _10542_ (.A0(_06173_),
    .A1(_06175_),
    .A2(_06176_),
    .A3(_06177_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06179_));
 sky130_fd_sc_hd__mux2i_1 _10543_ (.A0(_06172_),
    .A1(_06179_),
    .S(_05978_),
    .Y(_06180_));
 sky130_fd_sc_hd__nand2_1 _10544_ (.A(reset_hash),
    .B(\w[0][14] ),
    .Y(_06181_));
 sky130_fd_sc_hd__o21ai_0 _10545_ (.A1(_05482_),
    .A2(_06180_),
    .B1(_06181_),
    .Y(_00005_));
 sky130_fd_sc_hd__mux4_2 _10547_ (.A0(\w[18][15] ),
    .A1(\w[16][15] ),
    .A2(\w[22][15] ),
    .A3(\w[20][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06183_));
 sky130_fd_sc_hd__mux4_2 _10548_ (.A0(\w[26][15] ),
    .A1(\w[24][15] ),
    .A2(\w[30][15] ),
    .A3(\w[28][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06184_));
 sky130_fd_sc_hd__mux4_2 _10549_ (.A0(\w[2][15] ),
    .A1(\w[0][15] ),
    .A2(\w[6][15] ),
    .A3(\w[4][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06185_));
 sky130_fd_sc_hd__mux4_2 _10550_ (.A0(\w[10][15] ),
    .A1(\w[8][15] ),
    .A2(\w[14][15] ),
    .A3(\w[12][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06186_));
 sky130_fd_sc_hd__mux4_2 _10551_ (.A0(_06183_),
    .A1(_06184_),
    .A2(_06185_),
    .A3(_06186_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06187_));
 sky130_fd_sc_hd__mux4_2 _10552_ (.A0(\w[50][15] ),
    .A1(\w[48][15] ),
    .A2(\w[54][15] ),
    .A3(\w[52][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06188_));
 sky130_fd_sc_hd__mux4_2 _10554_ (.A0(\w[58][15] ),
    .A1(\w[56][15] ),
    .A2(\w[62][15] ),
    .A3(\w[60][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06190_));
 sky130_fd_sc_hd__mux4_2 _10555_ (.A0(\w[34][15] ),
    .A1(\w[32][15] ),
    .A2(\w[38][15] ),
    .A3(\w[36][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06191_));
 sky130_fd_sc_hd__mux4_2 _10556_ (.A0(\w[42][15] ),
    .A1(\w[40][15] ),
    .A2(\w[46][15] ),
    .A3(\w[44][15] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06192_));
 sky130_fd_sc_hd__mux4_2 _10557_ (.A0(_06188_),
    .A1(_06190_),
    .A2(_06191_),
    .A3(_06192_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06193_));
 sky130_fd_sc_hd__mux2i_1 _10558_ (.A0(_06187_),
    .A1(_06193_),
    .S(_05978_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_1 _10559_ (.A(reset_hash),
    .B(\w[0][15] ),
    .Y(_06195_));
 sky130_fd_sc_hd__o21ai_0 _10560_ (.A1(_05482_),
    .A2(_06194_),
    .B1(_06195_),
    .Y(_00006_));
 sky130_fd_sc_hd__mux4_2 _10561_ (.A0(\w[18][16] ),
    .A1(\w[16][16] ),
    .A2(\w[22][16] ),
    .A3(\w[20][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06196_));
 sky130_fd_sc_hd__mux4_2 _10563_ (.A0(\w[26][16] ),
    .A1(\w[24][16] ),
    .A2(\w[30][16] ),
    .A3(\w[28][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06198_));
 sky130_fd_sc_hd__mux4_2 _10564_ (.A0(\w[2][16] ),
    .A1(\w[0][16] ),
    .A2(\w[6][16] ),
    .A3(\w[4][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06199_));
 sky130_fd_sc_hd__mux4_2 _10565_ (.A0(\w[10][16] ),
    .A1(\w[8][16] ),
    .A2(\w[14][16] ),
    .A3(\w[12][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06200_));
 sky130_fd_sc_hd__mux4_2 _10567_ (.A0(_06196_),
    .A1(_06198_),
    .A2(_06199_),
    .A3(_06200_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06202_));
 sky130_fd_sc_hd__mux4_2 _10568_ (.A0(\w[50][16] ),
    .A1(\w[48][16] ),
    .A2(\w[54][16] ),
    .A3(\w[52][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06203_));
 sky130_fd_sc_hd__mux4_2 _10569_ (.A0(\w[58][16] ),
    .A1(\w[56][16] ),
    .A2(\w[62][16] ),
    .A3(\w[60][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06204_));
 sky130_fd_sc_hd__mux4_2 _10570_ (.A0(\w[34][16] ),
    .A1(\w[32][16] ),
    .A2(\w[38][16] ),
    .A3(\w[36][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06205_));
 sky130_fd_sc_hd__mux4_2 _10572_ (.A0(\w[42][16] ),
    .A1(\w[40][16] ),
    .A2(\w[46][16] ),
    .A3(\w[44][16] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06207_));
 sky130_fd_sc_hd__mux4_2 _10574_ (.A0(_06203_),
    .A1(_06204_),
    .A2(_06205_),
    .A3(_06207_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06209_));
 sky130_fd_sc_hd__mux2i_1 _10576_ (.A0(_06202_),
    .A1(_06209_),
    .S(_05978_),
    .Y(_06211_));
 sky130_fd_sc_hd__nand2_1 _10577_ (.A(reset_hash),
    .B(\w[0][16] ),
    .Y(_06212_));
 sky130_fd_sc_hd__o21ai_0 _10578_ (.A1(_05482_),
    .A2(_06211_),
    .B1(_06212_),
    .Y(_00007_));
 sky130_fd_sc_hd__mux4_2 _10579_ (.A0(\w[18][17] ),
    .A1(\w[16][17] ),
    .A2(\w[22][17] ),
    .A3(\w[20][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06213_));
 sky130_fd_sc_hd__mux4_2 _10581_ (.A0(\w[26][17] ),
    .A1(\w[24][17] ),
    .A2(\w[30][17] ),
    .A3(\w[28][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06215_));
 sky130_fd_sc_hd__mux4_2 _10582_ (.A0(\w[2][17] ),
    .A1(\w[0][17] ),
    .A2(\w[6][17] ),
    .A3(\w[4][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06216_));
 sky130_fd_sc_hd__mux4_2 _10583_ (.A0(\w[10][17] ),
    .A1(\w[8][17] ),
    .A2(\w[14][17] ),
    .A3(\w[12][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06217_));
 sky130_fd_sc_hd__mux4_2 _10584_ (.A0(_06213_),
    .A1(_06215_),
    .A2(_06216_),
    .A3(_06217_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06218_));
 sky130_fd_sc_hd__mux4_2 _10585_ (.A0(\w[50][17] ),
    .A1(\w[48][17] ),
    .A2(\w[54][17] ),
    .A3(\w[52][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06219_));
 sky130_fd_sc_hd__mux4_2 _10586_ (.A0(\w[58][17] ),
    .A1(\w[56][17] ),
    .A2(\w[62][17] ),
    .A3(\w[60][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06220_));
 sky130_fd_sc_hd__mux4_2 _10587_ (.A0(\w[34][17] ),
    .A1(\w[32][17] ),
    .A2(\w[38][17] ),
    .A3(\w[36][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06221_));
 sky130_fd_sc_hd__mux4_2 _10589_ (.A0(\w[42][17] ),
    .A1(\w[40][17] ),
    .A2(\w[46][17] ),
    .A3(\w[44][17] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06223_));
 sky130_fd_sc_hd__mux4_2 _10590_ (.A0(_06219_),
    .A1(_06220_),
    .A2(_06221_),
    .A3(_06223_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06224_));
 sky130_fd_sc_hd__mux2i_1 _10591_ (.A0(_06218_),
    .A1(_06224_),
    .S(_05978_),
    .Y(_06225_));
 sky130_fd_sc_hd__nand2_1 _10592_ (.A(reset_hash),
    .B(\w[0][17] ),
    .Y(_06226_));
 sky130_fd_sc_hd__o21ai_0 _10593_ (.A1(_05482_),
    .A2(_06225_),
    .B1(_06226_),
    .Y(_00008_));
 sky130_fd_sc_hd__mux4_2 _10594_ (.A0(\w[18][18] ),
    .A1(\w[16][18] ),
    .A2(\w[22][18] ),
    .A3(\w[20][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06227_));
 sky130_fd_sc_hd__mux4_2 _10595_ (.A0(\w[26][18] ),
    .A1(\w[24][18] ),
    .A2(\w[30][18] ),
    .A3(\w[28][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06228_));
 sky130_fd_sc_hd__mux4_2 _10596_ (.A0(\w[2][18] ),
    .A1(\w[0][18] ),
    .A2(\w[6][18] ),
    .A3(\w[4][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06229_));
 sky130_fd_sc_hd__mux4_2 _10598_ (.A0(\w[10][18] ),
    .A1(\w[8][18] ),
    .A2(\w[14][18] ),
    .A3(\w[12][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06231_));
 sky130_fd_sc_hd__mux4_2 _10600_ (.A0(_06227_),
    .A1(_06228_),
    .A2(_06229_),
    .A3(_06231_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06233_));
 sky130_fd_sc_hd__mux4_2 _10601_ (.A0(\w[50][18] ),
    .A1(\w[48][18] ),
    .A2(\w[54][18] ),
    .A3(\w[52][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06234_));
 sky130_fd_sc_hd__mux4_2 _10602_ (.A0(\w[58][18] ),
    .A1(\w[56][18] ),
    .A2(\w[62][18] ),
    .A3(\w[60][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06235_));
 sky130_fd_sc_hd__mux4_2 _10604_ (.A0(\w[34][18] ),
    .A1(\w[32][18] ),
    .A2(\w[38][18] ),
    .A3(\w[36][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06237_));
 sky130_fd_sc_hd__mux4_2 _10605_ (.A0(\w[42][18] ),
    .A1(\w[40][18] ),
    .A2(\w[46][18] ),
    .A3(\w[44][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06238_));
 sky130_fd_sc_hd__mux4_2 _10606_ (.A0(_06234_),
    .A1(_06235_),
    .A2(_06237_),
    .A3(_06238_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06239_));
 sky130_fd_sc_hd__mux2i_1 _10607_ (.A0(_06233_),
    .A1(_06239_),
    .S(_05978_),
    .Y(_06240_));
 sky130_fd_sc_hd__nand2_1 _10608_ (.A(reset_hash),
    .B(\w[0][18] ),
    .Y(_06241_));
 sky130_fd_sc_hd__o21ai_0 _10609_ (.A1(_05482_),
    .A2(_06240_),
    .B1(_06241_),
    .Y(_00009_));
 sky130_fd_sc_hd__mux4_2 _10610_ (.A0(\w[18][19] ),
    .A1(\w[16][19] ),
    .A2(\w[22][19] ),
    .A3(\w[20][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06242_));
 sky130_fd_sc_hd__mux4_2 _10611_ (.A0(\w[26][19] ),
    .A1(\w[24][19] ),
    .A2(\w[30][19] ),
    .A3(\w[28][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06243_));
 sky130_fd_sc_hd__mux4_2 _10612_ (.A0(\w[2][19] ),
    .A1(\w[0][19] ),
    .A2(\w[6][19] ),
    .A3(\w[4][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06244_));
 sky130_fd_sc_hd__mux4_2 _10614_ (.A0(\w[10][19] ),
    .A1(\w[8][19] ),
    .A2(\w[14][19] ),
    .A3(\w[12][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06246_));
 sky130_fd_sc_hd__mux4_2 _10615_ (.A0(_06242_),
    .A1(_06243_),
    .A2(_06244_),
    .A3(_06246_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06247_));
 sky130_fd_sc_hd__mux4_2 _10616_ (.A0(\w[50][19] ),
    .A1(\w[48][19] ),
    .A2(\w[54][19] ),
    .A3(\w[52][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06248_));
 sky130_fd_sc_hd__mux4_2 _10617_ (.A0(\w[58][19] ),
    .A1(\w[56][19] ),
    .A2(\w[62][19] ),
    .A3(\w[60][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06249_));
 sky130_fd_sc_hd__mux4_2 _10619_ (.A0(\w[34][19] ),
    .A1(\w[32][19] ),
    .A2(\w[38][19] ),
    .A3(\w[36][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06251_));
 sky130_fd_sc_hd__mux4_2 _10620_ (.A0(\w[42][19] ),
    .A1(\w[40][19] ),
    .A2(\w[46][19] ),
    .A3(\w[44][19] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06252_));
 sky130_fd_sc_hd__mux4_2 _10621_ (.A0(_06248_),
    .A1(_06249_),
    .A2(_06251_),
    .A3(_06252_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06253_));
 sky130_fd_sc_hd__mux2i_1 _10622_ (.A0(_06247_),
    .A1(_06253_),
    .S(_05978_),
    .Y(_06254_));
 sky130_fd_sc_hd__nand2_1 _10623_ (.A(reset_hash),
    .B(\w[0][19] ),
    .Y(_06255_));
 sky130_fd_sc_hd__o21ai_0 _10624_ (.A1(_05482_),
    .A2(_06254_),
    .B1(_06255_),
    .Y(_00010_));
 sky130_fd_sc_hd__mux4_2 _10626_ (.A0(\w[18][20] ),
    .A1(\w[16][20] ),
    .A2(\w[22][20] ),
    .A3(\w[20][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06257_));
 sky130_fd_sc_hd__mux4_2 _10627_ (.A0(\w[26][20] ),
    .A1(\w[24][20] ),
    .A2(\w[30][20] ),
    .A3(\w[28][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06258_));
 sky130_fd_sc_hd__mux4_2 _10628_ (.A0(\w[2][20] ),
    .A1(\w[0][20] ),
    .A2(\w[6][20] ),
    .A3(\w[4][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06259_));
 sky130_fd_sc_hd__mux4_2 _10629_ (.A0(\w[10][20] ),
    .A1(\w[8][20] ),
    .A2(\w[14][20] ),
    .A3(\w[12][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06260_));
 sky130_fd_sc_hd__mux4_2 _10630_ (.A0(_06257_),
    .A1(_06258_),
    .A2(_06259_),
    .A3(_06260_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06261_));
 sky130_fd_sc_hd__mux4_2 _10632_ (.A0(\w[50][20] ),
    .A1(\w[48][20] ),
    .A2(\w[54][20] ),
    .A3(\w[52][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06263_));
 sky130_fd_sc_hd__mux4_2 _10633_ (.A0(\w[58][20] ),
    .A1(\w[56][20] ),
    .A2(\w[62][20] ),
    .A3(\w[60][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06264_));
 sky130_fd_sc_hd__mux4_2 _10634_ (.A0(\w[34][20] ),
    .A1(\w[32][20] ),
    .A2(\w[38][20] ),
    .A3(\w[36][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06265_));
 sky130_fd_sc_hd__mux4_2 _10635_ (.A0(\w[42][20] ),
    .A1(\w[40][20] ),
    .A2(\w[46][20] ),
    .A3(\w[44][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06266_));
 sky130_fd_sc_hd__mux4_2 _10636_ (.A0(_06263_),
    .A1(_06264_),
    .A2(_06265_),
    .A3(_06266_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06267_));
 sky130_fd_sc_hd__mux2i_1 _10637_ (.A0(_06261_),
    .A1(_06267_),
    .S(_05978_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_1 _10638_ (.A(reset_hash),
    .B(\w[0][20] ),
    .Y(_06269_));
 sky130_fd_sc_hd__o21ai_0 _10639_ (.A1(_05482_),
    .A2(_06268_),
    .B1(_06269_),
    .Y(_00012_));
 sky130_fd_sc_hd__mux4_2 _10640_ (.A0(\w[18][21] ),
    .A1(\w[16][21] ),
    .A2(\w[22][21] ),
    .A3(\w[20][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06270_));
 sky130_fd_sc_hd__mux4_2 _10641_ (.A0(\w[26][21] ),
    .A1(\w[24][21] ),
    .A2(\w[30][21] ),
    .A3(\w[28][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06271_));
 sky130_fd_sc_hd__mux4_2 _10642_ (.A0(\w[2][21] ),
    .A1(\w[0][21] ),
    .A2(\w[6][21] ),
    .A3(\w[4][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06272_));
 sky130_fd_sc_hd__mux4_2 _10643_ (.A0(\w[10][21] ),
    .A1(\w[8][21] ),
    .A2(\w[14][21] ),
    .A3(\w[12][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06273_));
 sky130_fd_sc_hd__mux4_2 _10644_ (.A0(_06270_),
    .A1(_06271_),
    .A2(_06272_),
    .A3(_06273_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06274_));
 sky130_fd_sc_hd__mux4_2 _10646_ (.A0(\w[50][21] ),
    .A1(\w[48][21] ),
    .A2(\w[54][21] ),
    .A3(\w[52][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06276_));
 sky130_fd_sc_hd__mux4_2 _10647_ (.A0(\w[58][21] ),
    .A1(\w[56][21] ),
    .A2(\w[62][21] ),
    .A3(\w[60][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06277_));
 sky130_fd_sc_hd__mux4_2 _10648_ (.A0(\w[34][21] ),
    .A1(\w[32][21] ),
    .A2(\w[38][21] ),
    .A3(\w[36][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06278_));
 sky130_fd_sc_hd__mux4_2 _10649_ (.A0(\w[42][21] ),
    .A1(\w[40][21] ),
    .A2(\w[46][21] ),
    .A3(\w[44][21] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06279_));
 sky130_fd_sc_hd__mux4_2 _10650_ (.A0(_06276_),
    .A1(_06277_),
    .A2(_06278_),
    .A3(_06279_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06280_));
 sky130_fd_sc_hd__mux2i_1 _10651_ (.A0(_06274_),
    .A1(_06280_),
    .S(_05978_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_1 _10652_ (.A(reset_hash),
    .B(\w[0][21] ),
    .Y(_06282_));
 sky130_fd_sc_hd__o21ai_0 _10653_ (.A1(_05482_),
    .A2(_06281_),
    .B1(_06282_),
    .Y(_00013_));
 sky130_fd_sc_hd__mux4_2 _10654_ (.A0(\w[18][22] ),
    .A1(\w[16][22] ),
    .A2(\w[22][22] ),
    .A3(\w[20][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06283_));
 sky130_fd_sc_hd__mux4_2 _10655_ (.A0(\w[26][22] ),
    .A1(\w[24][22] ),
    .A2(\w[30][22] ),
    .A3(\w[28][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06284_));
 sky130_fd_sc_hd__mux4_2 _10657_ (.A0(\w[2][22] ),
    .A1(\w[0][22] ),
    .A2(\w[6][22] ),
    .A3(\w[4][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06286_));
 sky130_fd_sc_hd__mux4_2 _10658_ (.A0(\w[10][22] ),
    .A1(\w[8][22] ),
    .A2(\w[14][22] ),
    .A3(\w[12][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06287_));
 sky130_fd_sc_hd__mux4_2 _10659_ (.A0(_06283_),
    .A1(_06284_),
    .A2(_06286_),
    .A3(_06287_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06288_));
 sky130_fd_sc_hd__mux4_2 _10660_ (.A0(\w[50][22] ),
    .A1(\w[48][22] ),
    .A2(\w[54][22] ),
    .A3(\w[52][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06289_));
 sky130_fd_sc_hd__mux4_2 _10661_ (.A0(\w[58][22] ),
    .A1(\w[56][22] ),
    .A2(\w[62][22] ),
    .A3(\w[60][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06290_));
 sky130_fd_sc_hd__mux4_2 _10662_ (.A0(\w[34][22] ),
    .A1(\w[32][22] ),
    .A2(\w[38][22] ),
    .A3(\w[36][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06291_));
 sky130_fd_sc_hd__mux4_2 _10663_ (.A0(\w[42][22] ),
    .A1(\w[40][22] ),
    .A2(\w[46][22] ),
    .A3(\w[44][22] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06292_));
 sky130_fd_sc_hd__mux4_2 _10664_ (.A0(_06289_),
    .A1(_06290_),
    .A2(_06291_),
    .A3(_06292_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06293_));
 sky130_fd_sc_hd__mux2i_1 _10665_ (.A0(_06288_),
    .A1(_06293_),
    .S(_05978_),
    .Y(_06294_));
 sky130_fd_sc_hd__nand2_1 _10667_ (.A(reset_hash),
    .B(\w[0][22] ),
    .Y(_06296_));
 sky130_fd_sc_hd__o21ai_0 _10668_ (.A1(_05482_),
    .A2(_06294_),
    .B1(_06296_),
    .Y(_00014_));
 sky130_fd_sc_hd__mux4_2 _10669_ (.A0(\w[18][23] ),
    .A1(\w[16][23] ),
    .A2(\w[22][23] ),
    .A3(\w[20][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06297_));
 sky130_fd_sc_hd__mux4_2 _10670_ (.A0(\w[26][23] ),
    .A1(\w[24][23] ),
    .A2(\w[30][23] ),
    .A3(\w[28][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06298_));
 sky130_fd_sc_hd__mux4_2 _10671_ (.A0(\w[2][23] ),
    .A1(\w[0][23] ),
    .A2(\w[6][23] ),
    .A3(\w[4][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06299_));
 sky130_fd_sc_hd__mux4_2 _10672_ (.A0(\w[10][23] ),
    .A1(\w[8][23] ),
    .A2(\w[14][23] ),
    .A3(\w[12][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06300_));
 sky130_fd_sc_hd__mux4_2 _10673_ (.A0(_06297_),
    .A1(_06298_),
    .A2(_06299_),
    .A3(_06300_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06301_));
 sky130_fd_sc_hd__mux4_2 _10674_ (.A0(\w[50][23] ),
    .A1(\w[48][23] ),
    .A2(\w[54][23] ),
    .A3(\w[52][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06302_));
 sky130_fd_sc_hd__mux4_2 _10675_ (.A0(\w[58][23] ),
    .A1(\w[56][23] ),
    .A2(\w[62][23] ),
    .A3(\w[60][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06303_));
 sky130_fd_sc_hd__mux4_2 _10676_ (.A0(\w[34][23] ),
    .A1(\w[32][23] ),
    .A2(\w[38][23] ),
    .A3(\w[36][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06304_));
 sky130_fd_sc_hd__mux4_2 _10677_ (.A0(\w[42][23] ),
    .A1(\w[40][23] ),
    .A2(\w[46][23] ),
    .A3(\w[44][23] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06305_));
 sky130_fd_sc_hd__mux4_2 _10678_ (.A0(_06302_),
    .A1(_06303_),
    .A2(_06304_),
    .A3(_06305_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06306_));
 sky130_fd_sc_hd__mux2i_1 _10679_ (.A0(_06301_),
    .A1(_06306_),
    .S(_05978_),
    .Y(_06307_));
 sky130_fd_sc_hd__nand2_1 _10680_ (.A(reset_hash),
    .B(\w[0][23] ),
    .Y(_06308_));
 sky130_fd_sc_hd__o21ai_0 _10681_ (.A1(_05482_),
    .A2(_06307_),
    .B1(_06308_),
    .Y(_00015_));
 sky130_fd_sc_hd__mux4_2 _10682_ (.A0(\w[18][24] ),
    .A1(\w[16][24] ),
    .A2(\w[22][24] ),
    .A3(\w[20][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06309_));
 sky130_fd_sc_hd__mux4_2 _10683_ (.A0(\w[26][24] ),
    .A1(\w[24][24] ),
    .A2(\w[30][24] ),
    .A3(\w[28][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06310_));
 sky130_fd_sc_hd__mux4_2 _10684_ (.A0(\w[2][24] ),
    .A1(\w[0][24] ),
    .A2(\w[6][24] ),
    .A3(\w[4][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06311_));
 sky130_fd_sc_hd__mux4_2 _10685_ (.A0(\w[10][24] ),
    .A1(\w[8][24] ),
    .A2(\w[14][24] ),
    .A3(\w[12][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06312_));
 sky130_fd_sc_hd__mux4_2 _10686_ (.A0(_06309_),
    .A1(_06310_),
    .A2(_06311_),
    .A3(_06312_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06313_));
 sky130_fd_sc_hd__mux4_2 _10687_ (.A0(\w[50][24] ),
    .A1(\w[48][24] ),
    .A2(\w[54][24] ),
    .A3(\w[52][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06314_));
 sky130_fd_sc_hd__mux4_2 _10688_ (.A0(\w[58][24] ),
    .A1(\w[56][24] ),
    .A2(\w[62][24] ),
    .A3(\w[60][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06315_));
 sky130_fd_sc_hd__mux4_2 _10689_ (.A0(\w[34][24] ),
    .A1(\w[32][24] ),
    .A2(\w[38][24] ),
    .A3(\w[36][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06316_));
 sky130_fd_sc_hd__mux4_2 _10690_ (.A0(\w[42][24] ),
    .A1(\w[40][24] ),
    .A2(\w[46][24] ),
    .A3(\w[44][24] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06317_));
 sky130_fd_sc_hd__mux4_2 _10692_ (.A0(_06314_),
    .A1(_06315_),
    .A2(_06316_),
    .A3(_06317_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06319_));
 sky130_fd_sc_hd__mux2i_1 _10693_ (.A0(_06313_),
    .A1(_06319_),
    .S(_05978_),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_1 _10694_ (.A(reset_hash),
    .B(\w[0][24] ),
    .Y(_06321_));
 sky130_fd_sc_hd__o21ai_0 _10695_ (.A1(_05482_),
    .A2(_06320_),
    .B1(_06321_),
    .Y(_00016_));
 sky130_fd_sc_hd__mux4_2 _10696_ (.A0(\w[18][25] ),
    .A1(\w[16][25] ),
    .A2(\w[22][25] ),
    .A3(\w[20][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06322_));
 sky130_fd_sc_hd__mux4_2 _10697_ (.A0(\w[26][25] ),
    .A1(\w[24][25] ),
    .A2(\w[30][25] ),
    .A3(\w[28][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06323_));
 sky130_fd_sc_hd__mux4_2 _10698_ (.A0(\w[2][25] ),
    .A1(\w[0][25] ),
    .A2(\w[6][25] ),
    .A3(\w[4][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06324_));
 sky130_fd_sc_hd__mux4_2 _10699_ (.A0(\w[10][25] ),
    .A1(\w[8][25] ),
    .A2(\w[14][25] ),
    .A3(\w[12][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06325_));
 sky130_fd_sc_hd__mux4_2 _10700_ (.A0(_06322_),
    .A1(_06323_),
    .A2(_06324_),
    .A3(_06325_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06326_));
 sky130_fd_sc_hd__mux4_2 _10701_ (.A0(\w[50][25] ),
    .A1(\w[48][25] ),
    .A2(\w[54][25] ),
    .A3(\w[52][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06327_));
 sky130_fd_sc_hd__mux4_2 _10702_ (.A0(\w[58][25] ),
    .A1(\w[56][25] ),
    .A2(\w[62][25] ),
    .A3(\w[60][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06328_));
 sky130_fd_sc_hd__mux4_2 _10703_ (.A0(\w[34][25] ),
    .A1(\w[32][25] ),
    .A2(\w[38][25] ),
    .A3(\w[36][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06329_));
 sky130_fd_sc_hd__mux4_2 _10704_ (.A0(\w[42][25] ),
    .A1(\w[40][25] ),
    .A2(\w[46][25] ),
    .A3(\w[44][25] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06330_));
 sky130_fd_sc_hd__mux4_2 _10705_ (.A0(_06327_),
    .A1(_06328_),
    .A2(_06329_),
    .A3(_06330_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06331_));
 sky130_fd_sc_hd__mux2i_1 _10706_ (.A0(_06326_),
    .A1(_06331_),
    .S(_05978_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_1 _10707_ (.A(reset_hash),
    .B(\w[0][25] ),
    .Y(_06333_));
 sky130_fd_sc_hd__o21ai_0 _10708_ (.A1(_05482_),
    .A2(_06332_),
    .B1(_06333_),
    .Y(_00017_));
 sky130_fd_sc_hd__mux4_2 _10709_ (.A0(\w[18][26] ),
    .A1(\w[16][26] ),
    .A2(\w[22][26] ),
    .A3(\w[20][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06334_));
 sky130_fd_sc_hd__mux4_2 _10710_ (.A0(\w[26][26] ),
    .A1(\w[24][26] ),
    .A2(\w[30][26] ),
    .A3(\w[28][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06335_));
 sky130_fd_sc_hd__mux4_2 _10711_ (.A0(\w[2][26] ),
    .A1(\w[0][26] ),
    .A2(\w[6][26] ),
    .A3(\w[4][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06336_));
 sky130_fd_sc_hd__mux4_2 _10712_ (.A0(\w[10][26] ),
    .A1(\w[8][26] ),
    .A2(\w[14][26] ),
    .A3(\w[12][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06337_));
 sky130_fd_sc_hd__mux4_2 _10713_ (.A0(_06334_),
    .A1(_06335_),
    .A2(_06336_),
    .A3(_06337_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06338_));
 sky130_fd_sc_hd__mux4_2 _10714_ (.A0(\w[50][26] ),
    .A1(\w[48][26] ),
    .A2(\w[54][26] ),
    .A3(\w[52][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06339_));
 sky130_fd_sc_hd__mux4_2 _10715_ (.A0(\w[58][26] ),
    .A1(\w[56][26] ),
    .A2(\w[62][26] ),
    .A3(\w[60][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06340_));
 sky130_fd_sc_hd__mux4_2 _10716_ (.A0(\w[34][26] ),
    .A1(\w[32][26] ),
    .A2(\w[38][26] ),
    .A3(\w[36][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06341_));
 sky130_fd_sc_hd__mux4_2 _10717_ (.A0(\w[42][26] ),
    .A1(\w[40][26] ),
    .A2(\w[46][26] ),
    .A3(\w[44][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06342_));
 sky130_fd_sc_hd__mux4_2 _10719_ (.A0(_06339_),
    .A1(_06340_),
    .A2(_06341_),
    .A3(_06342_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06344_));
 sky130_fd_sc_hd__mux2i_1 _10721_ (.A0(_06338_),
    .A1(_06344_),
    .S(_05978_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand2_1 _10722_ (.A(reset_hash),
    .B(\w[0][26] ),
    .Y(_06347_));
 sky130_fd_sc_hd__o21ai_0 _10723_ (.A1(_05482_),
    .A2(_06346_),
    .B1(_06347_),
    .Y(_00018_));
 sky130_fd_sc_hd__mux4_2 _10724_ (.A0(\w[18][27] ),
    .A1(\w[16][27] ),
    .A2(\w[22][27] ),
    .A3(\w[20][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06348_));
 sky130_fd_sc_hd__mux4_2 _10725_ (.A0(\w[26][27] ),
    .A1(\w[24][27] ),
    .A2(\w[30][27] ),
    .A3(\w[28][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06349_));
 sky130_fd_sc_hd__mux4_2 _10726_ (.A0(\w[2][27] ),
    .A1(\w[0][27] ),
    .A2(\w[6][27] ),
    .A3(\w[4][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06350_));
 sky130_fd_sc_hd__mux4_2 _10727_ (.A0(\w[10][27] ),
    .A1(\w[8][27] ),
    .A2(\w[14][27] ),
    .A3(\w[12][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06351_));
 sky130_fd_sc_hd__mux4_2 _10728_ (.A0(_06348_),
    .A1(_06349_),
    .A2(_06350_),
    .A3(_06351_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06352_));
 sky130_fd_sc_hd__mux4_2 _10729_ (.A0(\w[50][27] ),
    .A1(\w[48][27] ),
    .A2(\w[54][27] ),
    .A3(\w[52][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06353_));
 sky130_fd_sc_hd__mux4_2 _10730_ (.A0(\w[58][27] ),
    .A1(\w[56][27] ),
    .A2(\w[62][27] ),
    .A3(\w[60][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06354_));
 sky130_fd_sc_hd__mux4_2 _10731_ (.A0(\w[34][27] ),
    .A1(\w[32][27] ),
    .A2(\w[38][27] ),
    .A3(\w[36][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06355_));
 sky130_fd_sc_hd__mux4_2 _10732_ (.A0(\w[42][27] ),
    .A1(\w[40][27] ),
    .A2(\w[46][27] ),
    .A3(\w[44][27] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06356_));
 sky130_fd_sc_hd__mux4_2 _10733_ (.A0(_06353_),
    .A1(_06354_),
    .A2(_06355_),
    .A3(_06356_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06357_));
 sky130_fd_sc_hd__mux2i_1 _10734_ (.A0(_06352_),
    .A1(_06357_),
    .S(_05978_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand2_1 _10735_ (.A(reset_hash),
    .B(\w[0][27] ),
    .Y(_06359_));
 sky130_fd_sc_hd__o21ai_0 _10736_ (.A1(_05482_),
    .A2(_06358_),
    .B1(_06359_),
    .Y(_00019_));
 sky130_fd_sc_hd__mux4_2 _10737_ (.A0(\w[18][28] ),
    .A1(\w[16][28] ),
    .A2(\w[22][28] ),
    .A3(\w[20][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06360_));
 sky130_fd_sc_hd__mux4_2 _10738_ (.A0(\w[26][28] ),
    .A1(\w[24][28] ),
    .A2(\w[30][28] ),
    .A3(\w[28][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06361_));
 sky130_fd_sc_hd__mux4_2 _10739_ (.A0(\w[2][28] ),
    .A1(\w[0][28] ),
    .A2(\w[6][28] ),
    .A3(\w[4][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06362_));
 sky130_fd_sc_hd__mux4_2 _10740_ (.A0(\w[10][28] ),
    .A1(\w[8][28] ),
    .A2(\w[14][28] ),
    .A3(\w[12][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06363_));
 sky130_fd_sc_hd__mux4_2 _10741_ (.A0(_06360_),
    .A1(_06361_),
    .A2(_06362_),
    .A3(_06363_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06364_));
 sky130_fd_sc_hd__mux4_2 _10742_ (.A0(\w[50][28] ),
    .A1(\w[48][28] ),
    .A2(\w[54][28] ),
    .A3(\w[52][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06365_));
 sky130_fd_sc_hd__mux4_2 _10743_ (.A0(\w[58][28] ),
    .A1(\w[56][28] ),
    .A2(\w[62][28] ),
    .A3(\w[60][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06366_));
 sky130_fd_sc_hd__mux4_2 _10744_ (.A0(\w[34][28] ),
    .A1(\w[32][28] ),
    .A2(\w[38][28] ),
    .A3(\w[36][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06367_));
 sky130_fd_sc_hd__mux4_2 _10745_ (.A0(\w[42][28] ),
    .A1(\w[40][28] ),
    .A2(\w[46][28] ),
    .A3(\w[44][28] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06368_));
 sky130_fd_sc_hd__mux4_2 _10746_ (.A0(_06365_),
    .A1(_06366_),
    .A2(_06367_),
    .A3(_06368_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06369_));
 sky130_fd_sc_hd__mux2i_1 _10747_ (.A0(_06364_),
    .A1(_06369_),
    .S(_05978_),
    .Y(_06370_));
 sky130_fd_sc_hd__nand2_1 _10748_ (.A(reset_hash),
    .B(\w[0][28] ),
    .Y(_06371_));
 sky130_fd_sc_hd__o21ai_0 _10749_ (.A1(_05482_),
    .A2(_06370_),
    .B1(_06371_),
    .Y(_00020_));
 sky130_fd_sc_hd__mux4_2 _10750_ (.A0(\w[18][29] ),
    .A1(\w[16][29] ),
    .A2(\w[22][29] ),
    .A3(\w[20][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06372_));
 sky130_fd_sc_hd__mux4_2 _10751_ (.A0(\w[26][29] ),
    .A1(\w[24][29] ),
    .A2(\w[30][29] ),
    .A3(\w[28][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06373_));
 sky130_fd_sc_hd__mux4_2 _10752_ (.A0(\w[2][29] ),
    .A1(\w[0][29] ),
    .A2(\w[6][29] ),
    .A3(\w[4][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06374_));
 sky130_fd_sc_hd__mux4_2 _10753_ (.A0(\w[10][29] ),
    .A1(\w[8][29] ),
    .A2(\w[14][29] ),
    .A3(\w[12][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06375_));
 sky130_fd_sc_hd__mux4_2 _10754_ (.A0(_06372_),
    .A1(_06373_),
    .A2(_06374_),
    .A3(_06375_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06376_));
 sky130_fd_sc_hd__mux4_2 _10755_ (.A0(\w[50][29] ),
    .A1(\w[48][29] ),
    .A2(\w[54][29] ),
    .A3(\w[52][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06377_));
 sky130_fd_sc_hd__mux4_2 _10756_ (.A0(\w[58][29] ),
    .A1(\w[56][29] ),
    .A2(\w[62][29] ),
    .A3(\w[60][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06378_));
 sky130_fd_sc_hd__mux4_2 _10757_ (.A0(\w[34][29] ),
    .A1(\w[32][29] ),
    .A2(\w[38][29] ),
    .A3(\w[36][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06379_));
 sky130_fd_sc_hd__mux4_2 _10758_ (.A0(\w[42][29] ),
    .A1(\w[40][29] ),
    .A2(\w[46][29] ),
    .A3(\w[44][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06380_));
 sky130_fd_sc_hd__mux4_2 _10759_ (.A0(_06377_),
    .A1(_06378_),
    .A2(_06379_),
    .A3(_06380_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06381_));
 sky130_fd_sc_hd__mux2i_1 _10760_ (.A0(_06376_),
    .A1(_06381_),
    .S(_05978_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_1 _10761_ (.A(reset_hash),
    .B(\w[0][29] ),
    .Y(_06383_));
 sky130_fd_sc_hd__o21ai_0 _10762_ (.A1(_05482_),
    .A2(_06382_),
    .B1(_06383_),
    .Y(_00021_));
 sky130_fd_sc_hd__mux4_2 _10763_ (.A0(\w[18][30] ),
    .A1(\w[16][30] ),
    .A2(\w[22][30] ),
    .A3(\w[20][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06384_));
 sky130_fd_sc_hd__mux4_2 _10764_ (.A0(\w[26][30] ),
    .A1(\w[24][30] ),
    .A2(\w[30][30] ),
    .A3(\w[28][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06385_));
 sky130_fd_sc_hd__mux4_2 _10765_ (.A0(\w[2][30] ),
    .A1(\w[0][30] ),
    .A2(\w[6][30] ),
    .A3(\w[4][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06386_));
 sky130_fd_sc_hd__mux4_2 _10766_ (.A0(\w[10][30] ),
    .A1(\w[8][30] ),
    .A2(\w[14][30] ),
    .A3(\w[12][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06387_));
 sky130_fd_sc_hd__mux4_2 _10767_ (.A0(_06384_),
    .A1(_06385_),
    .A2(_06386_),
    .A3(_06387_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06388_));
 sky130_fd_sc_hd__mux4_2 _10768_ (.A0(\w[50][30] ),
    .A1(\w[48][30] ),
    .A2(\w[54][30] ),
    .A3(\w[52][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06389_));
 sky130_fd_sc_hd__mux4_2 _10769_ (.A0(\w[58][30] ),
    .A1(\w[56][30] ),
    .A2(\w[62][30] ),
    .A3(\w[60][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06390_));
 sky130_fd_sc_hd__mux4_2 _10770_ (.A0(\w[34][30] ),
    .A1(\w[32][30] ),
    .A2(\w[38][30] ),
    .A3(\w[36][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06391_));
 sky130_fd_sc_hd__mux4_2 _10771_ (.A0(\w[42][30] ),
    .A1(\w[40][30] ),
    .A2(\w[46][30] ),
    .A3(\w[44][30] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06392_));
 sky130_fd_sc_hd__mux4_2 _10772_ (.A0(_06389_),
    .A1(_06390_),
    .A2(_06391_),
    .A3(_06392_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06393_));
 sky130_fd_sc_hd__mux2i_1 _10773_ (.A0(_06388_),
    .A1(_06393_),
    .S(_05978_),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2_1 _10774_ (.A(reset_hash),
    .B(\w[0][30] ),
    .Y(_06395_));
 sky130_fd_sc_hd__o21ai_0 _10775_ (.A1(_05482_),
    .A2(_06394_),
    .B1(_06395_),
    .Y(_00023_));
 sky130_fd_sc_hd__mux4_2 _10776_ (.A0(\w[18][31] ),
    .A1(\w[16][31] ),
    .A2(\w[22][31] ),
    .A3(\w[20][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06396_));
 sky130_fd_sc_hd__mux4_2 _10777_ (.A0(\w[26][31] ),
    .A1(\w[24][31] ),
    .A2(\w[30][31] ),
    .A3(\w[28][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06397_));
 sky130_fd_sc_hd__mux4_2 _10778_ (.A0(\w[2][31] ),
    .A1(\w[0][31] ),
    .A2(\w[6][31] ),
    .A3(\w[4][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06398_));
 sky130_fd_sc_hd__mux4_2 _10779_ (.A0(\w[10][31] ),
    .A1(\w[8][31] ),
    .A2(\w[14][31] ),
    .A3(\w[12][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06399_));
 sky130_fd_sc_hd__mux4_2 _10780_ (.A0(_06396_),
    .A1(_06397_),
    .A2(_06398_),
    .A3(_06399_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06400_));
 sky130_fd_sc_hd__mux4_2 _10781_ (.A0(\w[50][31] ),
    .A1(\w[48][31] ),
    .A2(\w[54][31] ),
    .A3(\w[52][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06401_));
 sky130_fd_sc_hd__mux4_2 _10782_ (.A0(\w[58][31] ),
    .A1(\w[56][31] ),
    .A2(\w[62][31] ),
    .A3(\w[60][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06402_));
 sky130_fd_sc_hd__mux4_2 _10783_ (.A0(\w[34][31] ),
    .A1(\w[32][31] ),
    .A2(\w[38][31] ),
    .A3(\w[36][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06403_));
 sky130_fd_sc_hd__mux4_2 _10784_ (.A0(\w[42][31] ),
    .A1(\w[40][31] ),
    .A2(\w[46][31] ),
    .A3(\w[44][31] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_06404_));
 sky130_fd_sc_hd__mux4_2 _10785_ (.A0(_06401_),
    .A1(_06402_),
    .A2(_06403_),
    .A3(_06404_),
    .S0(_05953_),
    .S1(_05958_),
    .X(_06405_));
 sky130_fd_sc_hd__mux2i_1 _10786_ (.A0(_06400_),
    .A1(_06405_),
    .S(_05978_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand2_1 _10787_ (.A(reset_hash),
    .B(\w[0][31] ),
    .Y(_06407_));
 sky130_fd_sc_hd__o21ai_0 _10788_ (.A1(_05482_),
    .A2(_06406_),
    .B1(_06407_),
    .Y(_00024_));
 sky130_fd_sc_hd__mux4_2 _10795_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06414_));
 sky130_fd_sc_hd__mux4_2 _10798_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06417_));
 sky130_fd_sc_hd__mux4_2 _10803_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06422_));
 sky130_fd_sc_hd__mux4_2 _10806_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06425_));
 sky130_fd_sc_hd__mux4_2 _10812_ (.A0(_06414_),
    .A1(_06417_),
    .A2(_06422_),
    .A3(_06425_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06431_));
 sky130_fd_sc_hd__mux4_2 _10815_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06434_));
 sky130_fd_sc_hd__mux4_2 _10818_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06437_));
 sky130_fd_sc_hd__mux4_2 _10821_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06440_));
 sky130_fd_sc_hd__mux4_2 _10825_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06444_));
 sky130_fd_sc_hd__mux4_2 _10828_ (.A0(_06434_),
    .A1(_06437_),
    .A2(_06440_),
    .A3(_06444_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06447_));
 sky130_fd_sc_hd__mux2_2 _10831_ (.A0(_06431_),
    .A1(_06447_),
    .S(\count16_1[5] ),
    .X(_08822_));
 sky130_fd_sc_hd__mux4_2 _10832_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06450_));
 sky130_fd_sc_hd__mux4_2 _10834_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06452_));
 sky130_fd_sc_hd__mux4_2 _10835_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06453_));
 sky130_fd_sc_hd__mux4_2 _10836_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06454_));
 sky130_fd_sc_hd__mux4_2 _10837_ (.A0(_06450_),
    .A1(_06452_),
    .A2(_06453_),
    .A3(_06454_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06455_));
 sky130_fd_sc_hd__mux4_2 _10838_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06456_));
 sky130_fd_sc_hd__mux4_2 _10839_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06457_));
 sky130_fd_sc_hd__mux4_2 _10840_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06458_));
 sky130_fd_sc_hd__mux4_2 _10841_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06459_));
 sky130_fd_sc_hd__mux4_2 _10842_ (.A0(_06456_),
    .A1(_06457_),
    .A2(_06458_),
    .A3(_06459_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06460_));
 sky130_fd_sc_hd__mux2_2 _10843_ (.A0(_06455_),
    .A1(_06460_),
    .S(\count16_1[5] ),
    .X(_08825_));
 sky130_fd_sc_hd__mux4_2 _10851_ (.A0(\w[1][1] ),
    .A1(\w[3][1] ),
    .A2(\w[5][1] ),
    .A3(\w[7][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06468_));
 sky130_fd_sc_hd__mux4_2 _10856_ (.A0(\w[9][1] ),
    .A1(\w[11][1] ),
    .A2(\w[13][1] ),
    .A3(\w[15][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06473_));
 sky130_fd_sc_hd__mux4_2 _10859_ (.A0(\w[17][1] ),
    .A1(\w[19][1] ),
    .A2(\w[21][1] ),
    .A3(\w[23][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06476_));
 sky130_fd_sc_hd__mux4_2 _10863_ (.A0(\w[25][1] ),
    .A1(\w[27][1] ),
    .A2(\w[29][1] ),
    .A3(\w[31][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06480_));
 sky130_fd_sc_hd__mux4_2 _10870_ (.A0(_06468_),
    .A1(_06473_),
    .A2(_06476_),
    .A3(_06480_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06487_));
 sky130_fd_sc_hd__mux4_2 _10873_ (.A0(\w[33][1] ),
    .A1(\w[35][1] ),
    .A2(\w[37][1] ),
    .A3(\w[39][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06490_));
 sky130_fd_sc_hd__mux4_2 _10876_ (.A0(\w[41][1] ),
    .A1(\w[43][1] ),
    .A2(\w[45][1] ),
    .A3(\w[47][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06493_));
 sky130_fd_sc_hd__mux4_2 _10879_ (.A0(\w[49][1] ),
    .A1(\w[51][1] ),
    .A2(\w[53][1] ),
    .A3(\w[55][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06496_));
 sky130_fd_sc_hd__mux4_2 _10882_ (.A0(\w[57][1] ),
    .A1(\w[59][1] ),
    .A2(\w[61][1] ),
    .A3(\w[63][1] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06499_));
 sky130_fd_sc_hd__mux4_2 _10885_ (.A0(_06490_),
    .A1(_06493_),
    .A2(_06496_),
    .A3(_06499_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06502_));
 sky130_fd_sc_hd__mux2i_1 _10888_ (.A0(_06487_),
    .A1(_06502_),
    .S(\count7_1[5] ),
    .Y(_08828_));
 sky130_fd_sc_hd__mux4_2 _10889_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06505_));
 sky130_fd_sc_hd__mux4_2 _10891_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06507_));
 sky130_fd_sc_hd__mux4_2 _10892_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06508_));
 sky130_fd_sc_hd__mux4_2 _10893_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06509_));
 sky130_fd_sc_hd__mux4_2 _10894_ (.A0(_06505_),
    .A1(_06507_),
    .A2(_06508_),
    .A3(_06509_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06510_));
 sky130_fd_sc_hd__mux4_2 _10895_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06511_));
 sky130_fd_sc_hd__mux4_2 _10897_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06513_));
 sky130_fd_sc_hd__mux4_2 _10898_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06514_));
 sky130_fd_sc_hd__mux4_2 _10899_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06515_));
 sky130_fd_sc_hd__mux4_2 _10900_ (.A0(_06511_),
    .A1(_06513_),
    .A2(_06514_),
    .A3(_06515_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06516_));
 sky130_fd_sc_hd__mux2_2 _10901_ (.A0(_06510_),
    .A1(_06516_),
    .S(\count16_1[5] ),
    .X(_08833_));
 sky130_fd_sc_hd__mux4_2 _10902_ (.A0(\w[1][2] ),
    .A1(\w[3][2] ),
    .A2(\w[5][2] ),
    .A3(\w[7][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06517_));
 sky130_fd_sc_hd__mux4_2 _10903_ (.A0(\w[9][2] ),
    .A1(\w[11][2] ),
    .A2(\w[13][2] ),
    .A3(\w[15][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06518_));
 sky130_fd_sc_hd__mux4_2 _10904_ (.A0(\w[17][2] ),
    .A1(\w[19][2] ),
    .A2(\w[21][2] ),
    .A3(\w[23][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06519_));
 sky130_fd_sc_hd__mux4_2 _10905_ (.A0(\w[25][2] ),
    .A1(\w[27][2] ),
    .A2(\w[29][2] ),
    .A3(\w[31][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06520_));
 sky130_fd_sc_hd__mux4_2 _10906_ (.A0(_06517_),
    .A1(_06518_),
    .A2(_06519_),
    .A3(_06520_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06521_));
 sky130_fd_sc_hd__mux4_2 _10907_ (.A0(\w[33][2] ),
    .A1(\w[35][2] ),
    .A2(\w[37][2] ),
    .A3(\w[39][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06522_));
 sky130_fd_sc_hd__mux4_2 _10908_ (.A0(\w[41][2] ),
    .A1(\w[43][2] ),
    .A2(\w[45][2] ),
    .A3(\w[47][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06523_));
 sky130_fd_sc_hd__mux4_2 _10909_ (.A0(\w[49][2] ),
    .A1(\w[51][2] ),
    .A2(\w[53][2] ),
    .A3(\w[55][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06524_));
 sky130_fd_sc_hd__mux4_2 _10910_ (.A0(\w[57][2] ),
    .A1(\w[59][2] ),
    .A2(\w[61][2] ),
    .A3(\w[63][2] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06525_));
 sky130_fd_sc_hd__mux4_2 _10911_ (.A0(_06522_),
    .A1(_06523_),
    .A2(_06524_),
    .A3(_06525_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06526_));
 sky130_fd_sc_hd__mux2i_1 _10912_ (.A0(_06521_),
    .A1(_06526_),
    .S(\count7_1[5] ),
    .Y(_08836_));
 sky130_fd_sc_hd__mux4_2 _10913_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06527_));
 sky130_fd_sc_hd__mux4_2 _10914_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06528_));
 sky130_fd_sc_hd__mux4_2 _10916_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06530_));
 sky130_fd_sc_hd__mux4_2 _10917_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06531_));
 sky130_fd_sc_hd__mux4_2 _10918_ (.A0(_06527_),
    .A1(_06528_),
    .A2(_06530_),
    .A3(_06531_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06532_));
 sky130_fd_sc_hd__mux4_2 _10919_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06533_));
 sky130_fd_sc_hd__mux4_2 _10921_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06535_));
 sky130_fd_sc_hd__mux4_2 _10922_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06536_));
 sky130_fd_sc_hd__mux4_2 _10923_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06537_));
 sky130_fd_sc_hd__mux4_2 _10924_ (.A0(_06533_),
    .A1(_06535_),
    .A2(_06536_),
    .A3(_06537_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06538_));
 sky130_fd_sc_hd__mux2_2 _10925_ (.A0(_06532_),
    .A1(_06538_),
    .S(\count16_1[5] ),
    .X(_08846_));
 sky130_fd_sc_hd__mux4_2 _10926_ (.A0(\w[1][3] ),
    .A1(\w[3][3] ),
    .A2(\w[5][3] ),
    .A3(\w[7][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06539_));
 sky130_fd_sc_hd__mux4_2 _10927_ (.A0(\w[9][3] ),
    .A1(\w[11][3] ),
    .A2(\w[13][3] ),
    .A3(\w[15][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06540_));
 sky130_fd_sc_hd__mux4_2 _10928_ (.A0(\w[17][3] ),
    .A1(\w[19][3] ),
    .A2(\w[21][3] ),
    .A3(\w[23][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06541_));
 sky130_fd_sc_hd__mux4_2 _10929_ (.A0(\w[25][3] ),
    .A1(\w[27][3] ),
    .A2(\w[29][3] ),
    .A3(\w[31][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06542_));
 sky130_fd_sc_hd__mux4_2 _10930_ (.A0(_06539_),
    .A1(_06540_),
    .A2(_06541_),
    .A3(_06542_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06543_));
 sky130_fd_sc_hd__mux4_2 _10931_ (.A0(\w[33][3] ),
    .A1(\w[35][3] ),
    .A2(\w[37][3] ),
    .A3(\w[39][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06544_));
 sky130_fd_sc_hd__mux4_2 _10932_ (.A0(\w[41][3] ),
    .A1(\w[43][3] ),
    .A2(\w[45][3] ),
    .A3(\w[47][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06545_));
 sky130_fd_sc_hd__mux4_2 _10933_ (.A0(\w[49][3] ),
    .A1(\w[51][3] ),
    .A2(\w[53][3] ),
    .A3(\w[55][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06546_));
 sky130_fd_sc_hd__mux4_2 _10934_ (.A0(\w[57][3] ),
    .A1(\w[59][3] ),
    .A2(\w[61][3] ),
    .A3(\w[63][3] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06547_));
 sky130_fd_sc_hd__mux4_2 _10935_ (.A0(_06544_),
    .A1(_06545_),
    .A2(_06546_),
    .A3(_06547_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06548_));
 sky130_fd_sc_hd__mux2i_1 _10936_ (.A0(_06543_),
    .A1(_06548_),
    .S(\count7_1[5] ),
    .Y(_08849_));
 sky130_fd_sc_hd__mux4_2 _10937_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06549_));
 sky130_fd_sc_hd__mux4_2 _10938_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06550_));
 sky130_fd_sc_hd__mux4_2 _10940_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06552_));
 sky130_fd_sc_hd__mux4_2 _10941_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06553_));
 sky130_fd_sc_hd__mux4_2 _10942_ (.A0(_06549_),
    .A1(_06550_),
    .A2(_06552_),
    .A3(_06553_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06554_));
 sky130_fd_sc_hd__mux4_2 _10943_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06555_));
 sky130_fd_sc_hd__mux4_2 _10944_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06556_));
 sky130_fd_sc_hd__mux4_2 _10946_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06558_));
 sky130_fd_sc_hd__mux4_2 _10947_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06559_));
 sky130_fd_sc_hd__mux4_2 _10948_ (.A0(_06555_),
    .A1(_06556_),
    .A2(_06558_),
    .A3(_06559_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06560_));
 sky130_fd_sc_hd__mux2_2 _10949_ (.A0(_06554_),
    .A1(_06560_),
    .S(\count16_1[5] ),
    .X(_08854_));
 sky130_fd_sc_hd__mux4_2 _10950_ (.A0(\w[1][4] ),
    .A1(\w[3][4] ),
    .A2(\w[5][4] ),
    .A3(\w[7][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06561_));
 sky130_fd_sc_hd__mux4_2 _10951_ (.A0(\w[9][4] ),
    .A1(\w[11][4] ),
    .A2(\w[13][4] ),
    .A3(\w[15][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06562_));
 sky130_fd_sc_hd__mux4_2 _10952_ (.A0(\w[17][4] ),
    .A1(\w[19][4] ),
    .A2(\w[21][4] ),
    .A3(\w[23][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06563_));
 sky130_fd_sc_hd__mux4_2 _10953_ (.A0(\w[25][4] ),
    .A1(\w[27][4] ),
    .A2(\w[29][4] ),
    .A3(\w[31][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06564_));
 sky130_fd_sc_hd__mux4_2 _10954_ (.A0(_06561_),
    .A1(_06562_),
    .A2(_06563_),
    .A3(_06564_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06565_));
 sky130_fd_sc_hd__mux4_2 _10955_ (.A0(\w[33][4] ),
    .A1(\w[35][4] ),
    .A2(\w[37][4] ),
    .A3(\w[39][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06566_));
 sky130_fd_sc_hd__mux4_2 _10956_ (.A0(\w[41][4] ),
    .A1(\w[43][4] ),
    .A2(\w[45][4] ),
    .A3(\w[47][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06567_));
 sky130_fd_sc_hd__mux4_2 _10957_ (.A0(\w[49][4] ),
    .A1(\w[51][4] ),
    .A2(\w[53][4] ),
    .A3(\w[55][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06568_));
 sky130_fd_sc_hd__mux4_2 _10958_ (.A0(\w[57][4] ),
    .A1(\w[59][4] ),
    .A2(\w[61][4] ),
    .A3(\w[63][4] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06569_));
 sky130_fd_sc_hd__mux4_2 _10959_ (.A0(_06566_),
    .A1(_06567_),
    .A2(_06568_),
    .A3(_06569_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06570_));
 sky130_fd_sc_hd__mux2i_1 _10960_ (.A0(_06565_),
    .A1(_06570_),
    .S(\count7_1[5] ),
    .Y(_08857_));
 sky130_fd_sc_hd__mux4_2 _10962_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06572_));
 sky130_fd_sc_hd__mux4_2 _10963_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06573_));
 sky130_fd_sc_hd__mux4_2 _10964_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06574_));
 sky130_fd_sc_hd__mux4_2 _10965_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06575_));
 sky130_fd_sc_hd__mux4_2 _10966_ (.A0(_06572_),
    .A1(_06573_),
    .A2(_06574_),
    .A3(_06575_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06576_));
 sky130_fd_sc_hd__mux4_2 _10967_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06577_));
 sky130_fd_sc_hd__mux4_2 _10968_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06578_));
 sky130_fd_sc_hd__mux4_2 _10970_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06580_));
 sky130_fd_sc_hd__mux4_2 _10971_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06581_));
 sky130_fd_sc_hd__mux4_2 _10972_ (.A0(_06577_),
    .A1(_06578_),
    .A2(_06580_),
    .A3(_06581_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06582_));
 sky130_fd_sc_hd__mux2_2 _10973_ (.A0(_06576_),
    .A1(_06582_),
    .S(\count16_1[5] ),
    .X(_08862_));
 sky130_fd_sc_hd__mux4_2 _10974_ (.A0(\w[1][5] ),
    .A1(\w[3][5] ),
    .A2(\w[5][5] ),
    .A3(\w[7][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06583_));
 sky130_fd_sc_hd__mux4_2 _10975_ (.A0(\w[9][5] ),
    .A1(\w[11][5] ),
    .A2(\w[13][5] ),
    .A3(\w[15][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06584_));
 sky130_fd_sc_hd__mux4_2 _10976_ (.A0(\w[17][5] ),
    .A1(\w[19][5] ),
    .A2(\w[21][5] ),
    .A3(\w[23][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06585_));
 sky130_fd_sc_hd__mux4_2 _10977_ (.A0(\w[25][5] ),
    .A1(\w[27][5] ),
    .A2(\w[29][5] ),
    .A3(\w[31][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06586_));
 sky130_fd_sc_hd__mux4_2 _10978_ (.A0(_06583_),
    .A1(_06584_),
    .A2(_06585_),
    .A3(_06586_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06587_));
 sky130_fd_sc_hd__mux4_2 _10979_ (.A0(\w[33][5] ),
    .A1(\w[35][5] ),
    .A2(\w[37][5] ),
    .A3(\w[39][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06588_));
 sky130_fd_sc_hd__mux4_2 _10980_ (.A0(\w[41][5] ),
    .A1(\w[43][5] ),
    .A2(\w[45][5] ),
    .A3(\w[47][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06589_));
 sky130_fd_sc_hd__mux4_2 _10981_ (.A0(\w[49][5] ),
    .A1(\w[51][5] ),
    .A2(\w[53][5] ),
    .A3(\w[55][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06590_));
 sky130_fd_sc_hd__mux4_2 _10982_ (.A0(\w[57][5] ),
    .A1(\w[59][5] ),
    .A2(\w[61][5] ),
    .A3(\w[63][5] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06591_));
 sky130_fd_sc_hd__mux4_2 _10983_ (.A0(_06588_),
    .A1(_06589_),
    .A2(_06590_),
    .A3(_06591_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06592_));
 sky130_fd_sc_hd__mux2i_1 _10984_ (.A0(_06587_),
    .A1(_06592_),
    .S(\count7_1[5] ),
    .Y(_08865_));
 sky130_fd_sc_hd__mux4_2 _10986_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06594_));
 sky130_fd_sc_hd__mux4_2 _10987_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06595_));
 sky130_fd_sc_hd__mux4_2 _10988_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06596_));
 sky130_fd_sc_hd__mux4_2 _10989_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06597_));
 sky130_fd_sc_hd__mux4_2 _10991_ (.A0(_06594_),
    .A1(_06595_),
    .A2(_06596_),
    .A3(_06597_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06599_));
 sky130_fd_sc_hd__mux4_2 _10993_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06601_));
 sky130_fd_sc_hd__mux4_2 _10994_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06602_));
 sky130_fd_sc_hd__mux4_2 _10995_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06603_));
 sky130_fd_sc_hd__mux4_2 _10996_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06604_));
 sky130_fd_sc_hd__mux4_2 _10997_ (.A0(_06601_),
    .A1(_06602_),
    .A2(_06603_),
    .A3(_06604_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06605_));
 sky130_fd_sc_hd__mux2_2 _10998_ (.A0(_06599_),
    .A1(_06605_),
    .S(\count16_1[5] ),
    .X(_08870_));
 sky130_fd_sc_hd__mux4_2 _10999_ (.A0(\w[1][6] ),
    .A1(\w[3][6] ),
    .A2(\w[5][6] ),
    .A3(\w[7][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06606_));
 sky130_fd_sc_hd__mux4_2 _11000_ (.A0(\w[9][6] ),
    .A1(\w[11][6] ),
    .A2(\w[13][6] ),
    .A3(\w[15][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06607_));
 sky130_fd_sc_hd__mux4_2 _11001_ (.A0(\w[17][6] ),
    .A1(\w[19][6] ),
    .A2(\w[21][6] ),
    .A3(\w[23][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06608_));
 sky130_fd_sc_hd__mux4_2 _11002_ (.A0(\w[25][6] ),
    .A1(\w[27][6] ),
    .A2(\w[29][6] ),
    .A3(\w[31][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06609_));
 sky130_fd_sc_hd__mux4_2 _11003_ (.A0(_06606_),
    .A1(_06607_),
    .A2(_06608_),
    .A3(_06609_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06610_));
 sky130_fd_sc_hd__mux4_2 _11004_ (.A0(\w[33][6] ),
    .A1(\w[35][6] ),
    .A2(\w[37][6] ),
    .A3(\w[39][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06611_));
 sky130_fd_sc_hd__mux4_2 _11005_ (.A0(\w[41][6] ),
    .A1(\w[43][6] ),
    .A2(\w[45][6] ),
    .A3(\w[47][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06612_));
 sky130_fd_sc_hd__mux4_2 _11006_ (.A0(\w[49][6] ),
    .A1(\w[51][6] ),
    .A2(\w[53][6] ),
    .A3(\w[55][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06613_));
 sky130_fd_sc_hd__mux4_2 _11007_ (.A0(\w[57][6] ),
    .A1(\w[59][6] ),
    .A2(\w[61][6] ),
    .A3(\w[63][6] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06614_));
 sky130_fd_sc_hd__mux4_2 _11008_ (.A0(_06611_),
    .A1(_06612_),
    .A2(_06613_),
    .A3(_06614_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06615_));
 sky130_fd_sc_hd__mux2i_1 _11009_ (.A0(_06610_),
    .A1(_06615_),
    .S(\count7_1[5] ),
    .Y(_08873_));
 sky130_fd_sc_hd__mux4_2 _11010_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06616_));
 sky130_fd_sc_hd__mux4_2 _11011_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06617_));
 sky130_fd_sc_hd__mux4_2 _11012_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06618_));
 sky130_fd_sc_hd__mux4_2 _11014_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06620_));
 sky130_fd_sc_hd__mux4_2 _11016_ (.A0(_06616_),
    .A1(_06617_),
    .A2(_06618_),
    .A3(_06620_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06622_));
 sky130_fd_sc_hd__mux4_2 _11018_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06624_));
 sky130_fd_sc_hd__mux4_2 _11019_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06625_));
 sky130_fd_sc_hd__mux4_2 _11020_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06626_));
 sky130_fd_sc_hd__mux4_2 _11021_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06627_));
 sky130_fd_sc_hd__mux4_2 _11023_ (.A0(_06624_),
    .A1(_06625_),
    .A2(_06626_),
    .A3(_06627_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06629_));
 sky130_fd_sc_hd__mux2_2 _11024_ (.A0(_06622_),
    .A1(_06629_),
    .S(\count16_1[5] ),
    .X(_08878_));
 sky130_fd_sc_hd__mux4_2 _11025_ (.A0(\w[1][7] ),
    .A1(\w[3][7] ),
    .A2(\w[5][7] ),
    .A3(\w[7][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06630_));
 sky130_fd_sc_hd__mux4_2 _11026_ (.A0(\w[9][7] ),
    .A1(\w[11][7] ),
    .A2(\w[13][7] ),
    .A3(\w[15][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06631_));
 sky130_fd_sc_hd__mux4_2 _11027_ (.A0(\w[17][7] ),
    .A1(\w[19][7] ),
    .A2(\w[21][7] ),
    .A3(\w[23][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06632_));
 sky130_fd_sc_hd__mux4_2 _11028_ (.A0(\w[25][7] ),
    .A1(\w[27][7] ),
    .A2(\w[29][7] ),
    .A3(\w[31][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06633_));
 sky130_fd_sc_hd__mux4_2 _11029_ (.A0(_06630_),
    .A1(_06631_),
    .A2(_06632_),
    .A3(_06633_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06634_));
 sky130_fd_sc_hd__mux4_2 _11030_ (.A0(\w[33][7] ),
    .A1(\w[35][7] ),
    .A2(\w[37][7] ),
    .A3(\w[39][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06635_));
 sky130_fd_sc_hd__mux4_2 _11031_ (.A0(\w[41][7] ),
    .A1(\w[43][7] ),
    .A2(\w[45][7] ),
    .A3(\w[47][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06636_));
 sky130_fd_sc_hd__mux4_2 _11032_ (.A0(\w[49][7] ),
    .A1(\w[51][7] ),
    .A2(\w[53][7] ),
    .A3(\w[55][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06637_));
 sky130_fd_sc_hd__mux4_2 _11033_ (.A0(\w[57][7] ),
    .A1(\w[59][7] ),
    .A2(\w[61][7] ),
    .A3(\w[63][7] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06638_));
 sky130_fd_sc_hd__mux4_2 _11034_ (.A0(_06635_),
    .A1(_06636_),
    .A2(_06637_),
    .A3(_06638_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06639_));
 sky130_fd_sc_hd__mux2i_1 _11035_ (.A0(_06634_),
    .A1(_06639_),
    .S(\count7_1[5] ),
    .Y(_08881_));
 sky130_fd_sc_hd__mux4_2 _11036_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06640_));
 sky130_fd_sc_hd__mux4_2 _11037_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06641_));
 sky130_fd_sc_hd__mux4_2 _11038_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06642_));
 sky130_fd_sc_hd__mux4_2 _11040_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06644_));
 sky130_fd_sc_hd__mux4_2 _11041_ (.A0(_06640_),
    .A1(_06641_),
    .A2(_06642_),
    .A3(_06644_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06645_));
 sky130_fd_sc_hd__mux4_2 _11042_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06646_));
 sky130_fd_sc_hd__mux4_2 _11043_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06647_));
 sky130_fd_sc_hd__mux4_2 _11044_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06648_));
 sky130_fd_sc_hd__mux4_2 _11046_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06650_));
 sky130_fd_sc_hd__mux4_2 _11048_ (.A0(_06646_),
    .A1(_06647_),
    .A2(_06648_),
    .A3(_06650_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06652_));
 sky130_fd_sc_hd__mux2_2 _11049_ (.A0(_06645_),
    .A1(_06652_),
    .S(\count16_1[5] ),
    .X(_08886_));
 sky130_fd_sc_hd__mux4_2 _11050_ (.A0(\w[1][8] ),
    .A1(\w[3][8] ),
    .A2(\w[5][8] ),
    .A3(\w[7][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06653_));
 sky130_fd_sc_hd__mux4_2 _11051_ (.A0(\w[9][8] ),
    .A1(\w[11][8] ),
    .A2(\w[13][8] ),
    .A3(\w[15][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06654_));
 sky130_fd_sc_hd__mux4_2 _11052_ (.A0(\w[17][8] ),
    .A1(\w[19][8] ),
    .A2(\w[21][8] ),
    .A3(\w[23][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06655_));
 sky130_fd_sc_hd__mux4_2 _11053_ (.A0(\w[25][8] ),
    .A1(\w[27][8] ),
    .A2(\w[29][8] ),
    .A3(\w[31][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06656_));
 sky130_fd_sc_hd__mux4_2 _11055_ (.A0(_06653_),
    .A1(_06654_),
    .A2(_06655_),
    .A3(_06656_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06658_));
 sky130_fd_sc_hd__mux4_2 _11056_ (.A0(\w[33][8] ),
    .A1(\w[35][8] ),
    .A2(\w[37][8] ),
    .A3(\w[39][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06659_));
 sky130_fd_sc_hd__mux4_2 _11057_ (.A0(\w[41][8] ),
    .A1(\w[43][8] ),
    .A2(\w[45][8] ),
    .A3(\w[47][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06660_));
 sky130_fd_sc_hd__mux4_2 _11058_ (.A0(\w[49][8] ),
    .A1(\w[51][8] ),
    .A2(\w[53][8] ),
    .A3(\w[55][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06661_));
 sky130_fd_sc_hd__mux4_2 _11059_ (.A0(\w[57][8] ),
    .A1(\w[59][8] ),
    .A2(\w[61][8] ),
    .A3(\w[63][8] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06662_));
 sky130_fd_sc_hd__mux4_2 _11061_ (.A0(_06659_),
    .A1(_06660_),
    .A2(_06661_),
    .A3(_06662_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06664_));
 sky130_fd_sc_hd__mux2i_1 _11062_ (.A0(_06658_),
    .A1(_06664_),
    .S(\count7_1[5] ),
    .Y(_08889_));
 sky130_fd_sc_hd__mux4_2 _11063_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06665_));
 sky130_fd_sc_hd__mux4_2 _11064_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06666_));
 sky130_fd_sc_hd__mux4_2 _11065_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06667_));
 sky130_fd_sc_hd__mux4_2 _11066_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06668_));
 sky130_fd_sc_hd__mux4_2 _11067_ (.A0(_06665_),
    .A1(_06666_),
    .A2(_06667_),
    .A3(_06668_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06669_));
 sky130_fd_sc_hd__mux4_2 _11068_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06670_));
 sky130_fd_sc_hd__mux4_2 _11069_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06671_));
 sky130_fd_sc_hd__mux4_2 _11070_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06672_));
 sky130_fd_sc_hd__mux4_2 _11072_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06674_));
 sky130_fd_sc_hd__mux4_2 _11073_ (.A0(_06670_),
    .A1(_06671_),
    .A2(_06672_),
    .A3(_06674_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06675_));
 sky130_fd_sc_hd__mux2_2 _11075_ (.A0(_06669_),
    .A1(_06675_),
    .S(\count16_1[5] ),
    .X(_08894_));
 sky130_fd_sc_hd__mux4_2 _11077_ (.A0(\w[1][9] ),
    .A1(\w[3][9] ),
    .A2(\w[5][9] ),
    .A3(\w[7][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06678_));
 sky130_fd_sc_hd__mux4_2 _11079_ (.A0(\w[9][9] ),
    .A1(\w[11][9] ),
    .A2(\w[13][9] ),
    .A3(\w[15][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06680_));
 sky130_fd_sc_hd__mux4_2 _11081_ (.A0(\w[17][9] ),
    .A1(\w[19][9] ),
    .A2(\w[21][9] ),
    .A3(\w[23][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06682_));
 sky130_fd_sc_hd__mux4_2 _11083_ (.A0(\w[25][9] ),
    .A1(\w[27][9] ),
    .A2(\w[29][9] ),
    .A3(\w[31][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06684_));
 sky130_fd_sc_hd__mux4_2 _11085_ (.A0(_06678_),
    .A1(_06680_),
    .A2(_06682_),
    .A3(_06684_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06686_));
 sky130_fd_sc_hd__mux4_2 _11087_ (.A0(\w[33][9] ),
    .A1(\w[35][9] ),
    .A2(\w[37][9] ),
    .A3(\w[39][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06688_));
 sky130_fd_sc_hd__mux4_2 _11089_ (.A0(\w[41][9] ),
    .A1(\w[43][9] ),
    .A2(\w[45][9] ),
    .A3(\w[47][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06690_));
 sky130_fd_sc_hd__mux4_2 _11091_ (.A0(\w[49][9] ),
    .A1(\w[51][9] ),
    .A2(\w[53][9] ),
    .A3(\w[55][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06692_));
 sky130_fd_sc_hd__mux4_2 _11093_ (.A0(\w[57][9] ),
    .A1(\w[59][9] ),
    .A2(\w[61][9] ),
    .A3(\w[63][9] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06694_));
 sky130_fd_sc_hd__mux4_2 _11095_ (.A0(_06688_),
    .A1(_06690_),
    .A2(_06692_),
    .A3(_06694_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06696_));
 sky130_fd_sc_hd__mux2i_1 _11096_ (.A0(_06686_),
    .A1(_06696_),
    .S(\count7_1[5] ),
    .Y(_08897_));
 sky130_fd_sc_hd__mux4_2 _11097_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06697_));
 sky130_fd_sc_hd__mux4_2 _11098_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06698_));
 sky130_fd_sc_hd__mux4_2 _11099_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06699_));
 sky130_fd_sc_hd__mux4_2 _11100_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06700_));
 sky130_fd_sc_hd__mux4_2 _11101_ (.A0(_06697_),
    .A1(_06698_),
    .A2(_06699_),
    .A3(_06700_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06701_));
 sky130_fd_sc_hd__mux4_2 _11102_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06702_));
 sky130_fd_sc_hd__mux4_2 _11103_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06703_));
 sky130_fd_sc_hd__mux4_2 _11104_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06704_));
 sky130_fd_sc_hd__mux4_2 _11105_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06705_));
 sky130_fd_sc_hd__mux4_2 _11106_ (.A0(_06702_),
    .A1(_06703_),
    .A2(_06704_),
    .A3(_06705_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06706_));
 sky130_fd_sc_hd__mux2_2 _11107_ (.A0(_06701_),
    .A1(_06706_),
    .S(\count16_1[5] ),
    .X(_08902_));
 sky130_fd_sc_hd__mux4_2 _11109_ (.A0(\w[1][10] ),
    .A1(\w[3][10] ),
    .A2(\w[5][10] ),
    .A3(\w[7][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06708_));
 sky130_fd_sc_hd__mux4_2 _11111_ (.A0(\w[9][10] ),
    .A1(\w[11][10] ),
    .A2(\w[13][10] ),
    .A3(\w[15][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06710_));
 sky130_fd_sc_hd__mux4_2 _11113_ (.A0(\w[17][10] ),
    .A1(\w[19][10] ),
    .A2(\w[21][10] ),
    .A3(\w[23][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06712_));
 sky130_fd_sc_hd__mux4_2 _11115_ (.A0(\w[25][10] ),
    .A1(\w[27][10] ),
    .A2(\w[29][10] ),
    .A3(\w[31][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06714_));
 sky130_fd_sc_hd__mux4_2 _11116_ (.A0(_06708_),
    .A1(_06710_),
    .A2(_06712_),
    .A3(_06714_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06715_));
 sky130_fd_sc_hd__mux4_2 _11118_ (.A0(\w[33][10] ),
    .A1(\w[35][10] ),
    .A2(\w[37][10] ),
    .A3(\w[39][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06717_));
 sky130_fd_sc_hd__mux4_2 _11120_ (.A0(\w[41][10] ),
    .A1(\w[43][10] ),
    .A2(\w[45][10] ),
    .A3(\w[47][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06719_));
 sky130_fd_sc_hd__mux4_2 _11122_ (.A0(\w[49][10] ),
    .A1(\w[51][10] ),
    .A2(\w[53][10] ),
    .A3(\w[55][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06721_));
 sky130_fd_sc_hd__mux4_2 _11124_ (.A0(\w[57][10] ),
    .A1(\w[59][10] ),
    .A2(\w[61][10] ),
    .A3(\w[63][10] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06723_));
 sky130_fd_sc_hd__mux4_2 _11125_ (.A0(_06717_),
    .A1(_06719_),
    .A2(_06721_),
    .A3(_06723_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06724_));
 sky130_fd_sc_hd__mux2i_1 _11126_ (.A0(_06715_),
    .A1(_06724_),
    .S(\count7_1[5] ),
    .Y(_08905_));
 sky130_fd_sc_hd__mux4_2 _11127_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06725_));
 sky130_fd_sc_hd__mux4_2 _11129_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06727_));
 sky130_fd_sc_hd__mux4_2 _11130_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06728_));
 sky130_fd_sc_hd__mux4_2 _11131_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06729_));
 sky130_fd_sc_hd__mux4_2 _11132_ (.A0(_06725_),
    .A1(_06727_),
    .A2(_06728_),
    .A3(_06729_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06730_));
 sky130_fd_sc_hd__mux4_2 _11133_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06731_));
 sky130_fd_sc_hd__mux4_2 _11134_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06732_));
 sky130_fd_sc_hd__mux4_2 _11135_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06733_));
 sky130_fd_sc_hd__mux4_2 _11136_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06734_));
 sky130_fd_sc_hd__mux4_2 _11137_ (.A0(_06731_),
    .A1(_06732_),
    .A2(_06733_),
    .A3(_06734_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06735_));
 sky130_fd_sc_hd__mux2_2 _11138_ (.A0(_06730_),
    .A1(_06735_),
    .S(\count16_1[5] ),
    .X(_08910_));
 sky130_fd_sc_hd__mux4_2 _11139_ (.A0(\w[1][11] ),
    .A1(\w[3][11] ),
    .A2(\w[5][11] ),
    .A3(\w[7][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06736_));
 sky130_fd_sc_hd__mux4_2 _11140_ (.A0(\w[9][11] ),
    .A1(\w[11][11] ),
    .A2(\w[13][11] ),
    .A3(\w[15][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06737_));
 sky130_fd_sc_hd__mux4_2 _11141_ (.A0(\w[17][11] ),
    .A1(\w[19][11] ),
    .A2(\w[21][11] ),
    .A3(\w[23][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06738_));
 sky130_fd_sc_hd__mux4_2 _11142_ (.A0(\w[25][11] ),
    .A1(\w[27][11] ),
    .A2(\w[29][11] ),
    .A3(\w[31][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06739_));
 sky130_fd_sc_hd__mux4_2 _11143_ (.A0(_06736_),
    .A1(_06737_),
    .A2(_06738_),
    .A3(_06739_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06740_));
 sky130_fd_sc_hd__mux4_2 _11144_ (.A0(\w[33][11] ),
    .A1(\w[35][11] ),
    .A2(\w[37][11] ),
    .A3(\w[39][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06741_));
 sky130_fd_sc_hd__mux4_2 _11145_ (.A0(\w[41][11] ),
    .A1(\w[43][11] ),
    .A2(\w[45][11] ),
    .A3(\w[47][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06742_));
 sky130_fd_sc_hd__mux4_2 _11146_ (.A0(\w[49][11] ),
    .A1(\w[51][11] ),
    .A2(\w[53][11] ),
    .A3(\w[55][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06743_));
 sky130_fd_sc_hd__mux4_2 _11147_ (.A0(\w[57][11] ),
    .A1(\w[59][11] ),
    .A2(\w[61][11] ),
    .A3(\w[63][11] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06744_));
 sky130_fd_sc_hd__mux4_2 _11148_ (.A0(_06741_),
    .A1(_06742_),
    .A2(_06743_),
    .A3(_06744_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06745_));
 sky130_fd_sc_hd__mux2i_1 _11150_ (.A0(_06740_),
    .A1(_06745_),
    .S(\count7_1[5] ),
    .Y(_08913_));
 sky130_fd_sc_hd__mux4_2 _11151_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06747_));
 sky130_fd_sc_hd__mux4_2 _11153_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06749_));
 sky130_fd_sc_hd__mux4_2 _11154_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06750_));
 sky130_fd_sc_hd__mux4_2 _11155_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06751_));
 sky130_fd_sc_hd__mux4_2 _11156_ (.A0(_06747_),
    .A1(_06749_),
    .A2(_06750_),
    .A3(_06751_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06752_));
 sky130_fd_sc_hd__mux4_2 _11157_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06753_));
 sky130_fd_sc_hd__mux4_2 _11159_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06755_));
 sky130_fd_sc_hd__mux4_2 _11160_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06756_));
 sky130_fd_sc_hd__mux4_2 _11161_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06757_));
 sky130_fd_sc_hd__mux4_2 _11162_ (.A0(_06753_),
    .A1(_06755_),
    .A2(_06756_),
    .A3(_06757_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06758_));
 sky130_fd_sc_hd__mux2_2 _11163_ (.A0(_06752_),
    .A1(_06758_),
    .S(\count16_1[5] ),
    .X(_08918_));
 sky130_fd_sc_hd__mux4_2 _11164_ (.A0(\w[1][12] ),
    .A1(\w[3][12] ),
    .A2(\w[5][12] ),
    .A3(\w[7][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06759_));
 sky130_fd_sc_hd__mux4_2 _11165_ (.A0(\w[9][12] ),
    .A1(\w[11][12] ),
    .A2(\w[13][12] ),
    .A3(\w[15][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06760_));
 sky130_fd_sc_hd__mux4_2 _11166_ (.A0(\w[17][12] ),
    .A1(\w[19][12] ),
    .A2(\w[21][12] ),
    .A3(\w[23][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06761_));
 sky130_fd_sc_hd__mux4_2 _11167_ (.A0(\w[25][12] ),
    .A1(\w[27][12] ),
    .A2(\w[29][12] ),
    .A3(\w[31][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06762_));
 sky130_fd_sc_hd__mux4_2 _11168_ (.A0(_06759_),
    .A1(_06760_),
    .A2(_06761_),
    .A3(_06762_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06763_));
 sky130_fd_sc_hd__mux4_2 _11169_ (.A0(\w[33][12] ),
    .A1(\w[35][12] ),
    .A2(\w[37][12] ),
    .A3(\w[39][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06764_));
 sky130_fd_sc_hd__mux4_2 _11170_ (.A0(\w[41][12] ),
    .A1(\w[43][12] ),
    .A2(\w[45][12] ),
    .A3(\w[47][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06765_));
 sky130_fd_sc_hd__mux4_2 _11171_ (.A0(\w[49][12] ),
    .A1(\w[51][12] ),
    .A2(\w[53][12] ),
    .A3(\w[55][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06766_));
 sky130_fd_sc_hd__mux4_2 _11172_ (.A0(\w[57][12] ),
    .A1(\w[59][12] ),
    .A2(\w[61][12] ),
    .A3(\w[63][12] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06767_));
 sky130_fd_sc_hd__mux4_2 _11173_ (.A0(_06764_),
    .A1(_06765_),
    .A2(_06766_),
    .A3(_06767_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06768_));
 sky130_fd_sc_hd__mux2i_1 _11174_ (.A0(_06763_),
    .A1(_06768_),
    .S(\count7_1[5] ),
    .Y(_08921_));
 sky130_fd_sc_hd__mux4_2 _11175_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06769_));
 sky130_fd_sc_hd__mux4_2 _11176_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06770_));
 sky130_fd_sc_hd__mux4_2 _11178_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06772_));
 sky130_fd_sc_hd__mux4_2 _11179_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06773_));
 sky130_fd_sc_hd__mux4_2 _11180_ (.A0(_06769_),
    .A1(_06770_),
    .A2(_06772_),
    .A3(_06773_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06774_));
 sky130_fd_sc_hd__mux4_2 _11181_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06775_));
 sky130_fd_sc_hd__mux4_2 _11183_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06777_));
 sky130_fd_sc_hd__mux4_2 _11184_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06778_));
 sky130_fd_sc_hd__mux4_2 _11185_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06779_));
 sky130_fd_sc_hd__mux4_2 _11186_ (.A0(_06775_),
    .A1(_06777_),
    .A2(_06778_),
    .A3(_06779_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06780_));
 sky130_fd_sc_hd__mux2_2 _11187_ (.A0(_06774_),
    .A1(_06780_),
    .S(\count16_1[5] ),
    .X(_08926_));
 sky130_fd_sc_hd__mux4_2 _11188_ (.A0(\w[1][13] ),
    .A1(\w[3][13] ),
    .A2(\w[5][13] ),
    .A3(\w[7][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06781_));
 sky130_fd_sc_hd__mux4_2 _11189_ (.A0(\w[9][13] ),
    .A1(\w[11][13] ),
    .A2(\w[13][13] ),
    .A3(\w[15][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06782_));
 sky130_fd_sc_hd__mux4_2 _11190_ (.A0(\w[17][13] ),
    .A1(\w[19][13] ),
    .A2(\w[21][13] ),
    .A3(\w[23][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06783_));
 sky130_fd_sc_hd__mux4_2 _11191_ (.A0(\w[25][13] ),
    .A1(\w[27][13] ),
    .A2(\w[29][13] ),
    .A3(\w[31][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06784_));
 sky130_fd_sc_hd__mux4_2 _11192_ (.A0(_06781_),
    .A1(_06782_),
    .A2(_06783_),
    .A3(_06784_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06785_));
 sky130_fd_sc_hd__mux4_2 _11193_ (.A0(\w[33][13] ),
    .A1(\w[35][13] ),
    .A2(\w[37][13] ),
    .A3(\w[39][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06786_));
 sky130_fd_sc_hd__mux4_2 _11194_ (.A0(\w[41][13] ),
    .A1(\w[43][13] ),
    .A2(\w[45][13] ),
    .A3(\w[47][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06787_));
 sky130_fd_sc_hd__mux4_2 _11195_ (.A0(\w[49][13] ),
    .A1(\w[51][13] ),
    .A2(\w[53][13] ),
    .A3(\w[55][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06788_));
 sky130_fd_sc_hd__mux4_2 _11196_ (.A0(\w[57][13] ),
    .A1(\w[59][13] ),
    .A2(\w[61][13] ),
    .A3(\w[63][13] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06789_));
 sky130_fd_sc_hd__mux4_2 _11197_ (.A0(_06786_),
    .A1(_06787_),
    .A2(_06788_),
    .A3(_06789_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06790_));
 sky130_fd_sc_hd__mux2i_1 _11198_ (.A0(_06785_),
    .A1(_06790_),
    .S(\count7_1[5] ),
    .Y(_08929_));
 sky130_fd_sc_hd__mux4_2 _11199_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06791_));
 sky130_fd_sc_hd__mux4_2 _11200_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06792_));
 sky130_fd_sc_hd__mux4_2 _11202_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06794_));
 sky130_fd_sc_hd__mux4_2 _11203_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06795_));
 sky130_fd_sc_hd__mux4_2 _11204_ (.A0(_06791_),
    .A1(_06792_),
    .A2(_06794_),
    .A3(_06795_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06796_));
 sky130_fd_sc_hd__mux4_2 _11205_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06797_));
 sky130_fd_sc_hd__mux4_2 _11206_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06798_));
 sky130_fd_sc_hd__mux4_2 _11208_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06800_));
 sky130_fd_sc_hd__mux4_2 _11209_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06801_));
 sky130_fd_sc_hd__mux4_2 _11210_ (.A0(_06797_),
    .A1(_06798_),
    .A2(_06800_),
    .A3(_06801_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06802_));
 sky130_fd_sc_hd__mux2_2 _11211_ (.A0(_06796_),
    .A1(_06802_),
    .S(\count16_1[5] ),
    .X(_08934_));
 sky130_fd_sc_hd__mux4_2 _11212_ (.A0(\w[1][14] ),
    .A1(\w[3][14] ),
    .A2(\w[5][14] ),
    .A3(\w[7][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06803_));
 sky130_fd_sc_hd__mux4_2 _11213_ (.A0(\w[9][14] ),
    .A1(\w[11][14] ),
    .A2(\w[13][14] ),
    .A3(\w[15][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06804_));
 sky130_fd_sc_hd__mux4_2 _11214_ (.A0(\w[17][14] ),
    .A1(\w[19][14] ),
    .A2(\w[21][14] ),
    .A3(\w[23][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06805_));
 sky130_fd_sc_hd__mux4_2 _11215_ (.A0(\w[25][14] ),
    .A1(\w[27][14] ),
    .A2(\w[29][14] ),
    .A3(\w[31][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06806_));
 sky130_fd_sc_hd__mux4_2 _11216_ (.A0(_06803_),
    .A1(_06804_),
    .A2(_06805_),
    .A3(_06806_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06807_));
 sky130_fd_sc_hd__mux4_2 _11217_ (.A0(\w[33][14] ),
    .A1(\w[35][14] ),
    .A2(\w[37][14] ),
    .A3(\w[39][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06808_));
 sky130_fd_sc_hd__mux4_2 _11218_ (.A0(\w[41][14] ),
    .A1(\w[43][14] ),
    .A2(\w[45][14] ),
    .A3(\w[47][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06809_));
 sky130_fd_sc_hd__mux4_2 _11219_ (.A0(\w[49][14] ),
    .A1(\w[51][14] ),
    .A2(\w[53][14] ),
    .A3(\w[55][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06810_));
 sky130_fd_sc_hd__mux4_2 _11220_ (.A0(\w[57][14] ),
    .A1(\w[59][14] ),
    .A2(\w[61][14] ),
    .A3(\w[63][14] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06811_));
 sky130_fd_sc_hd__mux4_2 _11221_ (.A0(_06808_),
    .A1(_06809_),
    .A2(_06810_),
    .A3(_06811_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06812_));
 sky130_fd_sc_hd__mux2i_1 _11222_ (.A0(_06807_),
    .A1(_06812_),
    .S(\count7_1[5] ),
    .Y(_08937_));
 sky130_fd_sc_hd__mux4_2 _11224_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06814_));
 sky130_fd_sc_hd__mux4_2 _11225_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06815_));
 sky130_fd_sc_hd__mux4_2 _11226_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06816_));
 sky130_fd_sc_hd__mux4_2 _11227_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06817_));
 sky130_fd_sc_hd__mux4_2 _11228_ (.A0(_06814_),
    .A1(_06815_),
    .A2(_06816_),
    .A3(_06817_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06818_));
 sky130_fd_sc_hd__mux4_2 _11229_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06819_));
 sky130_fd_sc_hd__mux4_2 _11230_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06820_));
 sky130_fd_sc_hd__mux4_2 _11232_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06822_));
 sky130_fd_sc_hd__mux4_2 _11233_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06823_));
 sky130_fd_sc_hd__mux4_2 _11234_ (.A0(_06819_),
    .A1(_06820_),
    .A2(_06822_),
    .A3(_06823_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06824_));
 sky130_fd_sc_hd__mux2_2 _11235_ (.A0(_06818_),
    .A1(_06824_),
    .S(\count16_1[5] ),
    .X(_08942_));
 sky130_fd_sc_hd__mux4_2 _11236_ (.A0(\w[1][15] ),
    .A1(\w[3][15] ),
    .A2(\w[5][15] ),
    .A3(\w[7][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06825_));
 sky130_fd_sc_hd__mux4_2 _11237_ (.A0(\w[9][15] ),
    .A1(\w[11][15] ),
    .A2(\w[13][15] ),
    .A3(\w[15][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06826_));
 sky130_fd_sc_hd__mux4_2 _11238_ (.A0(\w[17][15] ),
    .A1(\w[19][15] ),
    .A2(\w[21][15] ),
    .A3(\w[23][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06827_));
 sky130_fd_sc_hd__mux4_2 _11239_ (.A0(\w[25][15] ),
    .A1(\w[27][15] ),
    .A2(\w[29][15] ),
    .A3(\w[31][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06828_));
 sky130_fd_sc_hd__mux4_2 _11240_ (.A0(_06825_),
    .A1(_06826_),
    .A2(_06827_),
    .A3(_06828_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06829_));
 sky130_fd_sc_hd__mux4_2 _11241_ (.A0(\w[33][15] ),
    .A1(\w[35][15] ),
    .A2(\w[37][15] ),
    .A3(\w[39][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06830_));
 sky130_fd_sc_hd__mux4_2 _11242_ (.A0(\w[41][15] ),
    .A1(\w[43][15] ),
    .A2(\w[45][15] ),
    .A3(\w[47][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06831_));
 sky130_fd_sc_hd__mux4_2 _11243_ (.A0(\w[49][15] ),
    .A1(\w[51][15] ),
    .A2(\w[53][15] ),
    .A3(\w[55][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06832_));
 sky130_fd_sc_hd__mux4_2 _11244_ (.A0(\w[57][15] ),
    .A1(\w[59][15] ),
    .A2(\w[61][15] ),
    .A3(\w[63][15] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06833_));
 sky130_fd_sc_hd__mux4_2 _11245_ (.A0(_06830_),
    .A1(_06831_),
    .A2(_06832_),
    .A3(_06833_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06834_));
 sky130_fd_sc_hd__mux2i_1 _11246_ (.A0(_06829_),
    .A1(_06834_),
    .S(\count7_1[5] ),
    .Y(_08945_));
 sky130_fd_sc_hd__mux4_2 _11248_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06836_));
 sky130_fd_sc_hd__mux4_2 _11249_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06837_));
 sky130_fd_sc_hd__mux4_2 _11250_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06838_));
 sky130_fd_sc_hd__mux4_2 _11251_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06839_));
 sky130_fd_sc_hd__mux4_2 _11253_ (.A0(_06836_),
    .A1(_06837_),
    .A2(_06838_),
    .A3(_06839_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06841_));
 sky130_fd_sc_hd__mux4_2 _11255_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06843_));
 sky130_fd_sc_hd__mux4_2 _11256_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06844_));
 sky130_fd_sc_hd__mux4_2 _11257_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06845_));
 sky130_fd_sc_hd__mux4_2 _11258_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06846_));
 sky130_fd_sc_hd__mux4_2 _11259_ (.A0(_06843_),
    .A1(_06844_),
    .A2(_06845_),
    .A3(_06846_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06847_));
 sky130_fd_sc_hd__mux2_2 _11260_ (.A0(_06841_),
    .A1(_06847_),
    .S(\count16_1[5] ),
    .X(_08950_));
 sky130_fd_sc_hd__mux4_2 _11261_ (.A0(\w[1][16] ),
    .A1(\w[3][16] ),
    .A2(\w[5][16] ),
    .A3(\w[7][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06848_));
 sky130_fd_sc_hd__mux4_2 _11262_ (.A0(\w[9][16] ),
    .A1(\w[11][16] ),
    .A2(\w[13][16] ),
    .A3(\w[15][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06849_));
 sky130_fd_sc_hd__mux4_2 _11263_ (.A0(\w[17][16] ),
    .A1(\w[19][16] ),
    .A2(\w[21][16] ),
    .A3(\w[23][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06850_));
 sky130_fd_sc_hd__mux4_2 _11264_ (.A0(\w[25][16] ),
    .A1(\w[27][16] ),
    .A2(\w[29][16] ),
    .A3(\w[31][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06851_));
 sky130_fd_sc_hd__mux4_2 _11265_ (.A0(_06848_),
    .A1(_06849_),
    .A2(_06850_),
    .A3(_06851_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06852_));
 sky130_fd_sc_hd__mux4_2 _11266_ (.A0(\w[33][16] ),
    .A1(\w[35][16] ),
    .A2(\w[37][16] ),
    .A3(\w[39][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06853_));
 sky130_fd_sc_hd__mux4_2 _11267_ (.A0(\w[41][16] ),
    .A1(\w[43][16] ),
    .A2(\w[45][16] ),
    .A3(\w[47][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06854_));
 sky130_fd_sc_hd__mux4_2 _11268_ (.A0(\w[49][16] ),
    .A1(\w[51][16] ),
    .A2(\w[53][16] ),
    .A3(\w[55][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06855_));
 sky130_fd_sc_hd__mux4_2 _11269_ (.A0(\w[57][16] ),
    .A1(\w[59][16] ),
    .A2(\w[61][16] ),
    .A3(\w[63][16] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06856_));
 sky130_fd_sc_hd__mux4_2 _11270_ (.A0(_06853_),
    .A1(_06854_),
    .A2(_06855_),
    .A3(_06856_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06857_));
 sky130_fd_sc_hd__mux2i_1 _11271_ (.A0(_06852_),
    .A1(_06857_),
    .S(\count7_1[5] ),
    .Y(_08953_));
 sky130_fd_sc_hd__mux4_2 _11272_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06858_));
 sky130_fd_sc_hd__mux4_2 _11273_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06859_));
 sky130_fd_sc_hd__mux4_2 _11274_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06860_));
 sky130_fd_sc_hd__mux4_2 _11276_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06862_));
 sky130_fd_sc_hd__mux4_2 _11278_ (.A0(_06858_),
    .A1(_06859_),
    .A2(_06860_),
    .A3(_06862_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06864_));
 sky130_fd_sc_hd__mux4_2 _11280_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06866_));
 sky130_fd_sc_hd__mux4_2 _11281_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06867_));
 sky130_fd_sc_hd__mux4_2 _11282_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06868_));
 sky130_fd_sc_hd__mux4_2 _11283_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06869_));
 sky130_fd_sc_hd__mux4_2 _11285_ (.A0(_06866_),
    .A1(_06867_),
    .A2(_06868_),
    .A3(_06869_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06871_));
 sky130_fd_sc_hd__mux2_2 _11286_ (.A0(_06864_),
    .A1(_06871_),
    .S(\count16_1[5] ),
    .X(_08958_));
 sky130_fd_sc_hd__mux4_2 _11287_ (.A0(\w[1][17] ),
    .A1(\w[3][17] ),
    .A2(\w[5][17] ),
    .A3(\w[7][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06872_));
 sky130_fd_sc_hd__mux4_2 _11288_ (.A0(\w[9][17] ),
    .A1(\w[11][17] ),
    .A2(\w[13][17] ),
    .A3(\w[15][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06873_));
 sky130_fd_sc_hd__mux4_2 _11289_ (.A0(\w[17][17] ),
    .A1(\w[19][17] ),
    .A2(\w[21][17] ),
    .A3(\w[23][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06874_));
 sky130_fd_sc_hd__mux4_2 _11290_ (.A0(\w[25][17] ),
    .A1(\w[27][17] ),
    .A2(\w[29][17] ),
    .A3(\w[31][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06875_));
 sky130_fd_sc_hd__mux4_2 _11291_ (.A0(_06872_),
    .A1(_06873_),
    .A2(_06874_),
    .A3(_06875_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06876_));
 sky130_fd_sc_hd__mux4_2 _11292_ (.A0(\w[33][17] ),
    .A1(\w[35][17] ),
    .A2(\w[37][17] ),
    .A3(\w[39][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06877_));
 sky130_fd_sc_hd__mux4_2 _11293_ (.A0(\w[41][17] ),
    .A1(\w[43][17] ),
    .A2(\w[45][17] ),
    .A3(\w[47][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06878_));
 sky130_fd_sc_hd__mux4_2 _11294_ (.A0(\w[49][17] ),
    .A1(\w[51][17] ),
    .A2(\w[53][17] ),
    .A3(\w[55][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06879_));
 sky130_fd_sc_hd__mux4_2 _11295_ (.A0(\w[57][17] ),
    .A1(\w[59][17] ),
    .A2(\w[61][17] ),
    .A3(\w[63][17] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06880_));
 sky130_fd_sc_hd__mux4_2 _11296_ (.A0(_06877_),
    .A1(_06878_),
    .A2(_06879_),
    .A3(_06880_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06881_));
 sky130_fd_sc_hd__mux2i_1 _11297_ (.A0(_06876_),
    .A1(_06881_),
    .S(\count7_1[5] ),
    .Y(_08961_));
 sky130_fd_sc_hd__mux4_2 _11298_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06882_));
 sky130_fd_sc_hd__mux4_2 _11299_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06883_));
 sky130_fd_sc_hd__mux4_2 _11300_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06884_));
 sky130_fd_sc_hd__mux4_2 _11302_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06886_));
 sky130_fd_sc_hd__mux4_2 _11303_ (.A0(_06882_),
    .A1(_06883_),
    .A2(_06884_),
    .A3(_06886_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06887_));
 sky130_fd_sc_hd__mux4_2 _11304_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06888_));
 sky130_fd_sc_hd__mux4_2 _11305_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06889_));
 sky130_fd_sc_hd__mux4_2 _11306_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06890_));
 sky130_fd_sc_hd__mux4_2 _11308_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06892_));
 sky130_fd_sc_hd__mux4_2 _11310_ (.A0(_06888_),
    .A1(_06889_),
    .A2(_06890_),
    .A3(_06892_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06894_));
 sky130_fd_sc_hd__mux2_2 _11311_ (.A0(_06887_),
    .A1(_06894_),
    .S(\count16_1[5] ),
    .X(_08966_));
 sky130_fd_sc_hd__mux4_2 _11312_ (.A0(\w[1][18] ),
    .A1(\w[3][18] ),
    .A2(\w[5][18] ),
    .A3(\w[7][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06895_));
 sky130_fd_sc_hd__mux4_2 _11313_ (.A0(\w[9][18] ),
    .A1(\w[11][18] ),
    .A2(\w[13][18] ),
    .A3(\w[15][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06896_));
 sky130_fd_sc_hd__mux4_2 _11314_ (.A0(\w[17][18] ),
    .A1(\w[19][18] ),
    .A2(\w[21][18] ),
    .A3(\w[23][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06897_));
 sky130_fd_sc_hd__mux4_2 _11315_ (.A0(\w[25][18] ),
    .A1(\w[27][18] ),
    .A2(\w[29][18] ),
    .A3(\w[31][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06898_));
 sky130_fd_sc_hd__mux4_2 _11317_ (.A0(_06895_),
    .A1(_06896_),
    .A2(_06897_),
    .A3(_06898_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06900_));
 sky130_fd_sc_hd__mux4_2 _11318_ (.A0(\w[33][18] ),
    .A1(\w[35][18] ),
    .A2(\w[37][18] ),
    .A3(\w[39][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06901_));
 sky130_fd_sc_hd__mux4_2 _11319_ (.A0(\w[41][18] ),
    .A1(\w[43][18] ),
    .A2(\w[45][18] ),
    .A3(\w[47][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06902_));
 sky130_fd_sc_hd__mux4_2 _11320_ (.A0(\w[49][18] ),
    .A1(\w[51][18] ),
    .A2(\w[53][18] ),
    .A3(\w[55][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06903_));
 sky130_fd_sc_hd__mux4_2 _11321_ (.A0(\w[57][18] ),
    .A1(\w[59][18] ),
    .A2(\w[61][18] ),
    .A3(\w[63][18] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06904_));
 sky130_fd_sc_hd__mux4_2 _11323_ (.A0(_06901_),
    .A1(_06902_),
    .A2(_06903_),
    .A3(_06904_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06906_));
 sky130_fd_sc_hd__mux2i_1 _11324_ (.A0(_06900_),
    .A1(_06906_),
    .S(\count7_1[5] ),
    .Y(_08969_));
 sky130_fd_sc_hd__mux4_2 _11325_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06907_));
 sky130_fd_sc_hd__mux4_2 _11326_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06908_));
 sky130_fd_sc_hd__mux4_2 _11327_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06909_));
 sky130_fd_sc_hd__mux4_2 _11328_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06910_));
 sky130_fd_sc_hd__mux4_2 _11329_ (.A0(_06907_),
    .A1(_06908_),
    .A2(_06909_),
    .A3(_06910_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06911_));
 sky130_fd_sc_hd__mux4_2 _11330_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06912_));
 sky130_fd_sc_hd__mux4_2 _11331_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06913_));
 sky130_fd_sc_hd__mux4_2 _11332_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06914_));
 sky130_fd_sc_hd__mux4_2 _11334_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06916_));
 sky130_fd_sc_hd__mux4_2 _11335_ (.A0(_06912_),
    .A1(_06913_),
    .A2(_06914_),
    .A3(_06916_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06917_));
 sky130_fd_sc_hd__mux2_2 _11337_ (.A0(_06911_),
    .A1(_06917_),
    .S(\count16_1[5] ),
    .X(_08974_));
 sky130_fd_sc_hd__mux4_2 _11339_ (.A0(\w[1][19] ),
    .A1(\w[3][19] ),
    .A2(\w[5][19] ),
    .A3(\w[7][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06920_));
 sky130_fd_sc_hd__mux4_2 _11341_ (.A0(\w[9][19] ),
    .A1(\w[11][19] ),
    .A2(\w[13][19] ),
    .A3(\w[15][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06922_));
 sky130_fd_sc_hd__mux4_2 _11343_ (.A0(\w[17][19] ),
    .A1(\w[19][19] ),
    .A2(\w[21][19] ),
    .A3(\w[23][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06924_));
 sky130_fd_sc_hd__mux4_2 _11345_ (.A0(\w[25][19] ),
    .A1(\w[27][19] ),
    .A2(\w[29][19] ),
    .A3(\w[31][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06926_));
 sky130_fd_sc_hd__mux4_2 _11347_ (.A0(_06920_),
    .A1(_06922_),
    .A2(_06924_),
    .A3(_06926_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06928_));
 sky130_fd_sc_hd__mux4_2 _11349_ (.A0(\w[33][19] ),
    .A1(\w[35][19] ),
    .A2(\w[37][19] ),
    .A3(\w[39][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06930_));
 sky130_fd_sc_hd__mux4_2 _11351_ (.A0(\w[41][19] ),
    .A1(\w[43][19] ),
    .A2(\w[45][19] ),
    .A3(\w[47][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06932_));
 sky130_fd_sc_hd__mux4_2 _11353_ (.A0(\w[49][19] ),
    .A1(\w[51][19] ),
    .A2(\w[53][19] ),
    .A3(\w[55][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06934_));
 sky130_fd_sc_hd__mux4_2 _11355_ (.A0(\w[57][19] ),
    .A1(\w[59][19] ),
    .A2(\w[61][19] ),
    .A3(\w[63][19] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06936_));
 sky130_fd_sc_hd__mux4_2 _11357_ (.A0(_06930_),
    .A1(_06932_),
    .A2(_06934_),
    .A3(_06936_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06938_));
 sky130_fd_sc_hd__mux2i_1 _11358_ (.A0(_06928_),
    .A1(_06938_),
    .S(\count7_1[5] ),
    .Y(_08977_));
 sky130_fd_sc_hd__mux4_2 _11359_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06939_));
 sky130_fd_sc_hd__mux4_2 _11360_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06940_));
 sky130_fd_sc_hd__mux4_2 _11361_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06941_));
 sky130_fd_sc_hd__mux4_2 _11362_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06942_));
 sky130_fd_sc_hd__mux4_2 _11363_ (.A0(_06939_),
    .A1(_06940_),
    .A2(_06941_),
    .A3(_06942_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06943_));
 sky130_fd_sc_hd__mux4_2 _11364_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06944_));
 sky130_fd_sc_hd__mux4_2 _11365_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06945_));
 sky130_fd_sc_hd__mux4_2 _11366_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06946_));
 sky130_fd_sc_hd__mux4_2 _11367_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06947_));
 sky130_fd_sc_hd__mux4_2 _11368_ (.A0(_06944_),
    .A1(_06945_),
    .A2(_06946_),
    .A3(_06947_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06948_));
 sky130_fd_sc_hd__mux2_2 _11369_ (.A0(_06943_),
    .A1(_06948_),
    .S(\count16_1[5] ),
    .X(_08982_));
 sky130_fd_sc_hd__mux4_2 _11371_ (.A0(\w[1][20] ),
    .A1(\w[3][20] ),
    .A2(\w[5][20] ),
    .A3(\w[7][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06950_));
 sky130_fd_sc_hd__mux4_2 _11373_ (.A0(\w[9][20] ),
    .A1(\w[11][20] ),
    .A2(\w[13][20] ),
    .A3(\w[15][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06952_));
 sky130_fd_sc_hd__mux4_2 _11375_ (.A0(\w[17][20] ),
    .A1(\w[19][20] ),
    .A2(\w[21][20] ),
    .A3(\w[23][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06954_));
 sky130_fd_sc_hd__mux4_2 _11377_ (.A0(\w[25][20] ),
    .A1(\w[27][20] ),
    .A2(\w[29][20] ),
    .A3(\w[31][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06956_));
 sky130_fd_sc_hd__mux4_2 _11378_ (.A0(_06950_),
    .A1(_06952_),
    .A2(_06954_),
    .A3(_06956_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06957_));
 sky130_fd_sc_hd__mux4_2 _11380_ (.A0(\w[33][20] ),
    .A1(\w[35][20] ),
    .A2(\w[37][20] ),
    .A3(\w[39][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06959_));
 sky130_fd_sc_hd__mux4_2 _11382_ (.A0(\w[41][20] ),
    .A1(\w[43][20] ),
    .A2(\w[45][20] ),
    .A3(\w[47][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06961_));
 sky130_fd_sc_hd__mux4_2 _11384_ (.A0(\w[49][20] ),
    .A1(\w[51][20] ),
    .A2(\w[53][20] ),
    .A3(\w[55][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06963_));
 sky130_fd_sc_hd__mux4_2 _11386_ (.A0(\w[57][20] ),
    .A1(\w[59][20] ),
    .A2(\w[61][20] ),
    .A3(\w[63][20] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06965_));
 sky130_fd_sc_hd__mux4_2 _11387_ (.A0(_06959_),
    .A1(_06961_),
    .A2(_06963_),
    .A3(_06965_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06966_));
 sky130_fd_sc_hd__mux2i_1 _11388_ (.A0(_06957_),
    .A1(_06966_),
    .S(\count7_1[5] ),
    .Y(_08985_));
 sky130_fd_sc_hd__mux4_2 _11389_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06967_));
 sky130_fd_sc_hd__mux4_2 _11391_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06969_));
 sky130_fd_sc_hd__mux4_2 _11392_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06970_));
 sky130_fd_sc_hd__mux4_2 _11393_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06971_));
 sky130_fd_sc_hd__mux4_2 _11394_ (.A0(_06967_),
    .A1(_06969_),
    .A2(_06970_),
    .A3(_06971_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06972_));
 sky130_fd_sc_hd__mux4_2 _11395_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06973_));
 sky130_fd_sc_hd__mux4_2 _11396_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06974_));
 sky130_fd_sc_hd__mux4_2 _11397_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06975_));
 sky130_fd_sc_hd__mux4_2 _11398_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06976_));
 sky130_fd_sc_hd__mux4_2 _11399_ (.A0(_06973_),
    .A1(_06974_),
    .A2(_06975_),
    .A3(_06976_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06977_));
 sky130_fd_sc_hd__mux2_2 _11400_ (.A0(_06972_),
    .A1(_06977_),
    .S(\count16_1[5] ),
    .X(_08990_));
 sky130_fd_sc_hd__mux4_2 _11401_ (.A0(\w[1][21] ),
    .A1(\w[3][21] ),
    .A2(\w[5][21] ),
    .A3(\w[7][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06978_));
 sky130_fd_sc_hd__mux4_2 _11402_ (.A0(\w[9][21] ),
    .A1(\w[11][21] ),
    .A2(\w[13][21] ),
    .A3(\w[15][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06979_));
 sky130_fd_sc_hd__mux4_2 _11403_ (.A0(\w[17][21] ),
    .A1(\w[19][21] ),
    .A2(\w[21][21] ),
    .A3(\w[23][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06980_));
 sky130_fd_sc_hd__mux4_2 _11404_ (.A0(\w[25][21] ),
    .A1(\w[27][21] ),
    .A2(\w[29][21] ),
    .A3(\w[31][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06981_));
 sky130_fd_sc_hd__mux4_2 _11405_ (.A0(_06978_),
    .A1(_06979_),
    .A2(_06980_),
    .A3(_06981_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06982_));
 sky130_fd_sc_hd__mux4_2 _11406_ (.A0(\w[33][21] ),
    .A1(\w[35][21] ),
    .A2(\w[37][21] ),
    .A3(\w[39][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06983_));
 sky130_fd_sc_hd__mux4_2 _11407_ (.A0(\w[41][21] ),
    .A1(\w[43][21] ),
    .A2(\w[45][21] ),
    .A3(\w[47][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06984_));
 sky130_fd_sc_hd__mux4_2 _11408_ (.A0(\w[49][21] ),
    .A1(\w[51][21] ),
    .A2(\w[53][21] ),
    .A3(\w[55][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06985_));
 sky130_fd_sc_hd__mux4_2 _11409_ (.A0(\w[57][21] ),
    .A1(\w[59][21] ),
    .A2(\w[61][21] ),
    .A3(\w[63][21] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06986_));
 sky130_fd_sc_hd__mux4_2 _11410_ (.A0(_06983_),
    .A1(_06984_),
    .A2(_06985_),
    .A3(_06986_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_06987_));
 sky130_fd_sc_hd__mux2i_1 _11412_ (.A0(_06982_),
    .A1(_06987_),
    .S(\count7_1[5] ),
    .Y(_08993_));
 sky130_fd_sc_hd__mux4_2 _11413_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06989_));
 sky130_fd_sc_hd__mux4_2 _11414_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06990_));
 sky130_fd_sc_hd__mux4_2 _11415_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06991_));
 sky130_fd_sc_hd__mux4_2 _11416_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06992_));
 sky130_fd_sc_hd__mux4_2 _11417_ (.A0(_06989_),
    .A1(_06990_),
    .A2(_06991_),
    .A3(_06992_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06993_));
 sky130_fd_sc_hd__mux4_2 _11418_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06994_));
 sky130_fd_sc_hd__mux4_2 _11419_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06995_));
 sky130_fd_sc_hd__mux4_2 _11420_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06996_));
 sky130_fd_sc_hd__mux4_2 _11421_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_06997_));
 sky130_fd_sc_hd__mux4_2 _11422_ (.A0(_06994_),
    .A1(_06995_),
    .A2(_06996_),
    .A3(_06997_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_06998_));
 sky130_fd_sc_hd__mux2_2 _11423_ (.A0(_06993_),
    .A1(_06998_),
    .S(\count16_1[5] ),
    .X(_08998_));
 sky130_fd_sc_hd__mux4_2 _11424_ (.A0(\w[1][22] ),
    .A1(\w[3][22] ),
    .A2(\w[5][22] ),
    .A3(\w[7][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_06999_));
 sky130_fd_sc_hd__mux4_2 _11425_ (.A0(\w[9][22] ),
    .A1(\w[11][22] ),
    .A2(\w[13][22] ),
    .A3(\w[15][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07000_));
 sky130_fd_sc_hd__mux4_2 _11426_ (.A0(\w[17][22] ),
    .A1(\w[19][22] ),
    .A2(\w[21][22] ),
    .A3(\w[23][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07001_));
 sky130_fd_sc_hd__mux4_2 _11427_ (.A0(\w[25][22] ),
    .A1(\w[27][22] ),
    .A2(\w[29][22] ),
    .A3(\w[31][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07002_));
 sky130_fd_sc_hd__mux4_2 _11428_ (.A0(_06999_),
    .A1(_07000_),
    .A2(_07001_),
    .A3(_07002_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07003_));
 sky130_fd_sc_hd__mux4_2 _11429_ (.A0(\w[33][22] ),
    .A1(\w[35][22] ),
    .A2(\w[37][22] ),
    .A3(\w[39][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07004_));
 sky130_fd_sc_hd__mux4_2 _11430_ (.A0(\w[41][22] ),
    .A1(\w[43][22] ),
    .A2(\w[45][22] ),
    .A3(\w[47][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07005_));
 sky130_fd_sc_hd__mux4_2 _11431_ (.A0(\w[49][22] ),
    .A1(\w[51][22] ),
    .A2(\w[53][22] ),
    .A3(\w[55][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07006_));
 sky130_fd_sc_hd__mux4_2 _11432_ (.A0(\w[57][22] ),
    .A1(\w[59][22] ),
    .A2(\w[61][22] ),
    .A3(\w[63][22] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07007_));
 sky130_fd_sc_hd__mux4_2 _11433_ (.A0(_07004_),
    .A1(_07005_),
    .A2(_07006_),
    .A3(_07007_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07008_));
 sky130_fd_sc_hd__mux2i_1 _11434_ (.A0(_07003_),
    .A1(_07008_),
    .S(\count7_1[5] ),
    .Y(_09001_));
 sky130_fd_sc_hd__mux4_2 _11435_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07009_));
 sky130_fd_sc_hd__mux4_2 _11436_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07010_));
 sky130_fd_sc_hd__mux4_2 _11437_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07011_));
 sky130_fd_sc_hd__mux4_2 _11438_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07012_));
 sky130_fd_sc_hd__mux4_2 _11439_ (.A0(_07009_),
    .A1(_07010_),
    .A2(_07011_),
    .A3(_07012_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07013_));
 sky130_fd_sc_hd__mux4_2 _11440_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07014_));
 sky130_fd_sc_hd__mux4_2 _11441_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07015_));
 sky130_fd_sc_hd__mux4_2 _11442_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07016_));
 sky130_fd_sc_hd__mux4_2 _11443_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07017_));
 sky130_fd_sc_hd__mux4_2 _11444_ (.A0(_07014_),
    .A1(_07015_),
    .A2(_07016_),
    .A3(_07017_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07018_));
 sky130_fd_sc_hd__mux2_2 _11445_ (.A0(_07013_),
    .A1(_07018_),
    .S(\count16_1[5] ),
    .X(_09006_));
 sky130_fd_sc_hd__mux4_2 _11446_ (.A0(\w[1][23] ),
    .A1(\w[3][23] ),
    .A2(\w[5][23] ),
    .A3(\w[7][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07019_));
 sky130_fd_sc_hd__mux4_2 _11447_ (.A0(\w[9][23] ),
    .A1(\w[11][23] ),
    .A2(\w[13][23] ),
    .A3(\w[15][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07020_));
 sky130_fd_sc_hd__mux4_2 _11448_ (.A0(\w[17][23] ),
    .A1(\w[19][23] ),
    .A2(\w[21][23] ),
    .A3(\w[23][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07021_));
 sky130_fd_sc_hd__mux4_2 _11449_ (.A0(\w[25][23] ),
    .A1(\w[27][23] ),
    .A2(\w[29][23] ),
    .A3(\w[31][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07022_));
 sky130_fd_sc_hd__mux4_2 _11450_ (.A0(_07019_),
    .A1(_07020_),
    .A2(_07021_),
    .A3(_07022_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07023_));
 sky130_fd_sc_hd__mux4_2 _11451_ (.A0(\w[33][23] ),
    .A1(\w[35][23] ),
    .A2(\w[37][23] ),
    .A3(\w[39][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07024_));
 sky130_fd_sc_hd__mux4_2 _11452_ (.A0(\w[41][23] ),
    .A1(\w[43][23] ),
    .A2(\w[45][23] ),
    .A3(\w[47][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07025_));
 sky130_fd_sc_hd__mux4_2 _11453_ (.A0(\w[49][23] ),
    .A1(\w[51][23] ),
    .A2(\w[53][23] ),
    .A3(\w[55][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07026_));
 sky130_fd_sc_hd__mux4_2 _11454_ (.A0(\w[57][23] ),
    .A1(\w[59][23] ),
    .A2(\w[61][23] ),
    .A3(\w[63][23] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07027_));
 sky130_fd_sc_hd__mux4_2 _11455_ (.A0(_07024_),
    .A1(_07025_),
    .A2(_07026_),
    .A3(_07027_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07028_));
 sky130_fd_sc_hd__mux2i_1 _11456_ (.A0(_07023_),
    .A1(_07028_),
    .S(\count7_1[5] ),
    .Y(_09009_));
 sky130_fd_sc_hd__mux4_2 _11457_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07029_));
 sky130_fd_sc_hd__mux4_2 _11458_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07030_));
 sky130_fd_sc_hd__mux4_2 _11459_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07031_));
 sky130_fd_sc_hd__mux4_2 _11460_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07032_));
 sky130_fd_sc_hd__mux4_2 _11461_ (.A0(_07029_),
    .A1(_07030_),
    .A2(_07031_),
    .A3(_07032_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07033_));
 sky130_fd_sc_hd__mux4_2 _11462_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07034_));
 sky130_fd_sc_hd__mux4_2 _11463_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07035_));
 sky130_fd_sc_hd__mux4_2 _11464_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07036_));
 sky130_fd_sc_hd__mux4_2 _11465_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07037_));
 sky130_fd_sc_hd__mux4_2 _11466_ (.A0(_07034_),
    .A1(_07035_),
    .A2(_07036_),
    .A3(_07037_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07038_));
 sky130_fd_sc_hd__mux2_2 _11467_ (.A0(_07033_),
    .A1(_07038_),
    .S(\count16_1[5] ),
    .X(_09014_));
 sky130_fd_sc_hd__mux4_2 _11468_ (.A0(\w[1][24] ),
    .A1(\w[3][24] ),
    .A2(\w[5][24] ),
    .A3(\w[7][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07039_));
 sky130_fd_sc_hd__mux4_2 _11469_ (.A0(\w[9][24] ),
    .A1(\w[11][24] ),
    .A2(\w[13][24] ),
    .A3(\w[15][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07040_));
 sky130_fd_sc_hd__mux4_2 _11470_ (.A0(\w[17][24] ),
    .A1(\w[19][24] ),
    .A2(\w[21][24] ),
    .A3(\w[23][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07041_));
 sky130_fd_sc_hd__mux4_2 _11471_ (.A0(\w[25][24] ),
    .A1(\w[27][24] ),
    .A2(\w[29][24] ),
    .A3(\w[31][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07042_));
 sky130_fd_sc_hd__mux4_2 _11472_ (.A0(_07039_),
    .A1(_07040_),
    .A2(_07041_),
    .A3(_07042_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07043_));
 sky130_fd_sc_hd__mux4_2 _11473_ (.A0(\w[33][24] ),
    .A1(\w[35][24] ),
    .A2(\w[37][24] ),
    .A3(\w[39][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07044_));
 sky130_fd_sc_hd__mux4_2 _11474_ (.A0(\w[41][24] ),
    .A1(\w[43][24] ),
    .A2(\w[45][24] ),
    .A3(\w[47][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07045_));
 sky130_fd_sc_hd__mux4_2 _11475_ (.A0(\w[49][24] ),
    .A1(\w[51][24] ),
    .A2(\w[53][24] ),
    .A3(\w[55][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07046_));
 sky130_fd_sc_hd__mux4_2 _11476_ (.A0(\w[57][24] ),
    .A1(\w[59][24] ),
    .A2(\w[61][24] ),
    .A3(\w[63][24] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07047_));
 sky130_fd_sc_hd__mux4_2 _11477_ (.A0(_07044_),
    .A1(_07045_),
    .A2(_07046_),
    .A3(_07047_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07048_));
 sky130_fd_sc_hd__mux2i_1 _11478_ (.A0(_07043_),
    .A1(_07048_),
    .S(\count7_1[5] ),
    .Y(_09017_));
 sky130_fd_sc_hd__mux4_2 _11479_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07049_));
 sky130_fd_sc_hd__mux4_2 _11480_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07050_));
 sky130_fd_sc_hd__mux4_2 _11481_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07051_));
 sky130_fd_sc_hd__mux4_2 _11482_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07052_));
 sky130_fd_sc_hd__mux4_2 _11483_ (.A0(_07049_),
    .A1(_07050_),
    .A2(_07051_),
    .A3(_07052_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07053_));
 sky130_fd_sc_hd__mux4_2 _11484_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07054_));
 sky130_fd_sc_hd__mux4_2 _11485_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07055_));
 sky130_fd_sc_hd__mux4_2 _11486_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07056_));
 sky130_fd_sc_hd__mux4_2 _11487_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07057_));
 sky130_fd_sc_hd__mux4_2 _11488_ (.A0(_07054_),
    .A1(_07055_),
    .A2(_07056_),
    .A3(_07057_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07058_));
 sky130_fd_sc_hd__mux2_2 _11489_ (.A0(_07053_),
    .A1(_07058_),
    .S(\count16_1[5] ),
    .X(_09022_));
 sky130_fd_sc_hd__mux4_2 _11490_ (.A0(\w[1][25] ),
    .A1(\w[3][25] ),
    .A2(\w[5][25] ),
    .A3(\w[7][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07059_));
 sky130_fd_sc_hd__mux4_2 _11491_ (.A0(\w[9][25] ),
    .A1(\w[11][25] ),
    .A2(\w[13][25] ),
    .A3(\w[15][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07060_));
 sky130_fd_sc_hd__mux4_2 _11492_ (.A0(\w[17][25] ),
    .A1(\w[19][25] ),
    .A2(\w[21][25] ),
    .A3(\w[23][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07061_));
 sky130_fd_sc_hd__mux4_2 _11493_ (.A0(\w[25][25] ),
    .A1(\w[27][25] ),
    .A2(\w[29][25] ),
    .A3(\w[31][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07062_));
 sky130_fd_sc_hd__mux4_2 _11494_ (.A0(_07059_),
    .A1(_07060_),
    .A2(_07061_),
    .A3(_07062_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07063_));
 sky130_fd_sc_hd__mux4_2 _11495_ (.A0(\w[33][25] ),
    .A1(\w[35][25] ),
    .A2(\w[37][25] ),
    .A3(\w[39][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07064_));
 sky130_fd_sc_hd__mux4_2 _11496_ (.A0(\w[41][25] ),
    .A1(\w[43][25] ),
    .A2(\w[45][25] ),
    .A3(\w[47][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07065_));
 sky130_fd_sc_hd__mux4_2 _11497_ (.A0(\w[49][25] ),
    .A1(\w[51][25] ),
    .A2(\w[53][25] ),
    .A3(\w[55][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07066_));
 sky130_fd_sc_hd__mux4_2 _11498_ (.A0(\w[57][25] ),
    .A1(\w[59][25] ),
    .A2(\w[61][25] ),
    .A3(\w[63][25] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07067_));
 sky130_fd_sc_hd__mux4_2 _11499_ (.A0(_07064_),
    .A1(_07065_),
    .A2(_07066_),
    .A3(_07067_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07068_));
 sky130_fd_sc_hd__mux2i_1 _11500_ (.A0(_07063_),
    .A1(_07068_),
    .S(\count7_1[5] ),
    .Y(_09025_));
 sky130_fd_sc_hd__mux4_2 _11501_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07069_));
 sky130_fd_sc_hd__mux4_2 _11502_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07070_));
 sky130_fd_sc_hd__mux4_2 _11503_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07071_));
 sky130_fd_sc_hd__mux4_2 _11504_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07072_));
 sky130_fd_sc_hd__mux4_2 _11505_ (.A0(_07069_),
    .A1(_07070_),
    .A2(_07071_),
    .A3(_07072_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07073_));
 sky130_fd_sc_hd__mux4_2 _11506_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07074_));
 sky130_fd_sc_hd__mux4_2 _11507_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07075_));
 sky130_fd_sc_hd__mux4_2 _11508_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07076_));
 sky130_fd_sc_hd__mux4_2 _11509_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07077_));
 sky130_fd_sc_hd__mux4_2 _11510_ (.A0(_07074_),
    .A1(_07075_),
    .A2(_07076_),
    .A3(_07077_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07078_));
 sky130_fd_sc_hd__mux2_2 _11511_ (.A0(_07073_),
    .A1(_07078_),
    .S(\count16_1[5] ),
    .X(_09030_));
 sky130_fd_sc_hd__mux4_2 _11512_ (.A0(\w[1][26] ),
    .A1(\w[3][26] ),
    .A2(\w[5][26] ),
    .A3(\w[7][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07079_));
 sky130_fd_sc_hd__mux4_2 _11513_ (.A0(\w[9][26] ),
    .A1(\w[11][26] ),
    .A2(\w[13][26] ),
    .A3(\w[15][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07080_));
 sky130_fd_sc_hd__mux4_2 _11514_ (.A0(\w[17][26] ),
    .A1(\w[19][26] ),
    .A2(\w[21][26] ),
    .A3(\w[23][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07081_));
 sky130_fd_sc_hd__mux4_2 _11515_ (.A0(\w[25][26] ),
    .A1(\w[27][26] ),
    .A2(\w[29][26] ),
    .A3(\w[31][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07082_));
 sky130_fd_sc_hd__mux4_2 _11516_ (.A0(_07079_),
    .A1(_07080_),
    .A2(_07081_),
    .A3(_07082_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07083_));
 sky130_fd_sc_hd__mux4_2 _11517_ (.A0(\w[33][26] ),
    .A1(\w[35][26] ),
    .A2(\w[37][26] ),
    .A3(\w[39][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07084_));
 sky130_fd_sc_hd__mux4_2 _11518_ (.A0(\w[41][26] ),
    .A1(\w[43][26] ),
    .A2(\w[45][26] ),
    .A3(\w[47][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07085_));
 sky130_fd_sc_hd__mux4_2 _11519_ (.A0(\w[49][26] ),
    .A1(\w[51][26] ),
    .A2(\w[53][26] ),
    .A3(\w[55][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07086_));
 sky130_fd_sc_hd__mux4_2 _11520_ (.A0(\w[57][26] ),
    .A1(\w[59][26] ),
    .A2(\w[61][26] ),
    .A3(\w[63][26] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07087_));
 sky130_fd_sc_hd__mux4_2 _11521_ (.A0(_07084_),
    .A1(_07085_),
    .A2(_07086_),
    .A3(_07087_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07088_));
 sky130_fd_sc_hd__mux2i_1 _11522_ (.A0(_07083_),
    .A1(_07088_),
    .S(\count7_1[5] ),
    .Y(_09033_));
 sky130_fd_sc_hd__mux4_2 _11523_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07089_));
 sky130_fd_sc_hd__mux4_2 _11524_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07090_));
 sky130_fd_sc_hd__mux4_2 _11525_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07091_));
 sky130_fd_sc_hd__mux4_2 _11526_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07092_));
 sky130_fd_sc_hd__mux4_2 _11527_ (.A0(_07089_),
    .A1(_07090_),
    .A2(_07091_),
    .A3(_07092_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07093_));
 sky130_fd_sc_hd__mux4_2 _11528_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07094_));
 sky130_fd_sc_hd__mux4_2 _11529_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07095_));
 sky130_fd_sc_hd__mux4_2 _11530_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07096_));
 sky130_fd_sc_hd__mux4_2 _11531_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07097_));
 sky130_fd_sc_hd__mux4_2 _11532_ (.A0(_07094_),
    .A1(_07095_),
    .A2(_07096_),
    .A3(_07097_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07098_));
 sky130_fd_sc_hd__mux2_2 _11533_ (.A0(_07093_),
    .A1(_07098_),
    .S(\count16_1[5] ),
    .X(_09038_));
 sky130_fd_sc_hd__mux4_2 _11534_ (.A0(\w[1][27] ),
    .A1(\w[3][27] ),
    .A2(\w[5][27] ),
    .A3(\w[7][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07099_));
 sky130_fd_sc_hd__mux4_2 _11535_ (.A0(\w[9][27] ),
    .A1(\w[11][27] ),
    .A2(\w[13][27] ),
    .A3(\w[15][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07100_));
 sky130_fd_sc_hd__mux4_2 _11536_ (.A0(\w[17][27] ),
    .A1(\w[19][27] ),
    .A2(\w[21][27] ),
    .A3(\w[23][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07101_));
 sky130_fd_sc_hd__mux4_2 _11537_ (.A0(\w[25][27] ),
    .A1(\w[27][27] ),
    .A2(\w[29][27] ),
    .A3(\w[31][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07102_));
 sky130_fd_sc_hd__mux4_2 _11538_ (.A0(_07099_),
    .A1(_07100_),
    .A2(_07101_),
    .A3(_07102_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07103_));
 sky130_fd_sc_hd__mux4_2 _11539_ (.A0(\w[33][27] ),
    .A1(\w[35][27] ),
    .A2(\w[37][27] ),
    .A3(\w[39][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07104_));
 sky130_fd_sc_hd__mux4_2 _11540_ (.A0(\w[41][27] ),
    .A1(\w[43][27] ),
    .A2(\w[45][27] ),
    .A3(\w[47][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07105_));
 sky130_fd_sc_hd__mux4_2 _11541_ (.A0(\w[49][27] ),
    .A1(\w[51][27] ),
    .A2(\w[53][27] ),
    .A3(\w[55][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07106_));
 sky130_fd_sc_hd__mux4_2 _11542_ (.A0(\w[57][27] ),
    .A1(\w[59][27] ),
    .A2(\w[61][27] ),
    .A3(\w[63][27] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07107_));
 sky130_fd_sc_hd__mux4_2 _11543_ (.A0(_07104_),
    .A1(_07105_),
    .A2(_07106_),
    .A3(_07107_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07108_));
 sky130_fd_sc_hd__mux2i_1 _11544_ (.A0(_07103_),
    .A1(_07108_),
    .S(\count7_1[5] ),
    .Y(_09041_));
 sky130_fd_sc_hd__mux4_2 _11545_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07109_));
 sky130_fd_sc_hd__mux4_2 _11546_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07110_));
 sky130_fd_sc_hd__mux4_2 _11547_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07111_));
 sky130_fd_sc_hd__mux4_2 _11548_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07112_));
 sky130_fd_sc_hd__mux4_2 _11549_ (.A0(_07109_),
    .A1(_07110_),
    .A2(_07111_),
    .A3(_07112_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07113_));
 sky130_fd_sc_hd__mux4_2 _11550_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07114_));
 sky130_fd_sc_hd__mux4_2 _11551_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07115_));
 sky130_fd_sc_hd__mux4_2 _11552_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07116_));
 sky130_fd_sc_hd__mux4_2 _11553_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07117_));
 sky130_fd_sc_hd__mux4_2 _11554_ (.A0(_07114_),
    .A1(_07115_),
    .A2(_07116_),
    .A3(_07117_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07118_));
 sky130_fd_sc_hd__mux2_2 _11555_ (.A0(_07113_),
    .A1(_07118_),
    .S(\count16_1[5] ),
    .X(_09046_));
 sky130_fd_sc_hd__mux4_2 _11556_ (.A0(\w[1][28] ),
    .A1(\w[3][28] ),
    .A2(\w[5][28] ),
    .A3(\w[7][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07119_));
 sky130_fd_sc_hd__mux4_2 _11557_ (.A0(\w[9][28] ),
    .A1(\w[11][28] ),
    .A2(\w[13][28] ),
    .A3(\w[15][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07120_));
 sky130_fd_sc_hd__mux4_2 _11558_ (.A0(\w[17][28] ),
    .A1(\w[19][28] ),
    .A2(\w[21][28] ),
    .A3(\w[23][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07121_));
 sky130_fd_sc_hd__mux4_2 _11559_ (.A0(\w[25][28] ),
    .A1(\w[27][28] ),
    .A2(\w[29][28] ),
    .A3(\w[31][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07122_));
 sky130_fd_sc_hd__mux4_2 _11560_ (.A0(_07119_),
    .A1(_07120_),
    .A2(_07121_),
    .A3(_07122_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07123_));
 sky130_fd_sc_hd__mux4_2 _11561_ (.A0(\w[33][28] ),
    .A1(\w[35][28] ),
    .A2(\w[37][28] ),
    .A3(\w[39][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07124_));
 sky130_fd_sc_hd__mux4_2 _11562_ (.A0(\w[41][28] ),
    .A1(\w[43][28] ),
    .A2(\w[45][28] ),
    .A3(\w[47][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07125_));
 sky130_fd_sc_hd__mux4_2 _11563_ (.A0(\w[49][28] ),
    .A1(\w[51][28] ),
    .A2(\w[53][28] ),
    .A3(\w[55][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07126_));
 sky130_fd_sc_hd__mux4_2 _11564_ (.A0(\w[57][28] ),
    .A1(\w[59][28] ),
    .A2(\w[61][28] ),
    .A3(\w[63][28] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07127_));
 sky130_fd_sc_hd__mux4_2 _11565_ (.A0(_07124_),
    .A1(_07125_),
    .A2(_07126_),
    .A3(_07127_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07128_));
 sky130_fd_sc_hd__mux2i_1 _11566_ (.A0(_07123_),
    .A1(_07128_),
    .S(\count7_1[5] ),
    .Y(_09049_));
 sky130_fd_sc_hd__mux4_2 _11567_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07129_));
 sky130_fd_sc_hd__mux4_2 _11568_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07130_));
 sky130_fd_sc_hd__mux4_2 _11569_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07131_));
 sky130_fd_sc_hd__mux4_2 _11570_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07132_));
 sky130_fd_sc_hd__mux4_2 _11571_ (.A0(_07129_),
    .A1(_07130_),
    .A2(_07131_),
    .A3(_07132_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07133_));
 sky130_fd_sc_hd__mux4_2 _11572_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07134_));
 sky130_fd_sc_hd__mux4_2 _11573_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07135_));
 sky130_fd_sc_hd__mux4_2 _11574_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07136_));
 sky130_fd_sc_hd__mux4_2 _11575_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07137_));
 sky130_fd_sc_hd__mux4_2 _11576_ (.A0(_07134_),
    .A1(_07135_),
    .A2(_07136_),
    .A3(_07137_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07138_));
 sky130_fd_sc_hd__mux2_2 _11577_ (.A0(_07133_),
    .A1(_07138_),
    .S(\count16_1[5] ),
    .X(_09054_));
 sky130_fd_sc_hd__mux4_2 _11578_ (.A0(\w[1][29] ),
    .A1(\w[3][29] ),
    .A2(\w[5][29] ),
    .A3(\w[7][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07139_));
 sky130_fd_sc_hd__mux4_2 _11579_ (.A0(\w[9][29] ),
    .A1(\w[11][29] ),
    .A2(\w[13][29] ),
    .A3(\w[15][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07140_));
 sky130_fd_sc_hd__mux4_2 _11580_ (.A0(\w[17][29] ),
    .A1(\w[19][29] ),
    .A2(\w[21][29] ),
    .A3(\w[23][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07141_));
 sky130_fd_sc_hd__mux4_2 _11581_ (.A0(\w[25][29] ),
    .A1(\w[27][29] ),
    .A2(\w[29][29] ),
    .A3(\w[31][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07142_));
 sky130_fd_sc_hd__mux4_2 _11582_ (.A0(_07139_),
    .A1(_07140_),
    .A2(_07141_),
    .A3(_07142_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07143_));
 sky130_fd_sc_hd__mux4_2 _11583_ (.A0(\w[33][29] ),
    .A1(\w[35][29] ),
    .A2(\w[37][29] ),
    .A3(\w[39][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07144_));
 sky130_fd_sc_hd__mux4_2 _11585_ (.A0(\w[41][29] ),
    .A1(\w[43][29] ),
    .A2(\w[45][29] ),
    .A3(\w[47][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07146_));
 sky130_fd_sc_hd__mux4_2 _11586_ (.A0(\w[49][29] ),
    .A1(\w[51][29] ),
    .A2(\w[53][29] ),
    .A3(\w[55][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07147_));
 sky130_fd_sc_hd__mux4_2 _11587_ (.A0(\w[57][29] ),
    .A1(\w[59][29] ),
    .A2(\w[61][29] ),
    .A3(\w[63][29] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07148_));
 sky130_fd_sc_hd__mux4_2 _11588_ (.A0(_07144_),
    .A1(_07146_),
    .A2(_07147_),
    .A3(_07148_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07149_));
 sky130_fd_sc_hd__mux2i_1 _11589_ (.A0(_07143_),
    .A1(_07149_),
    .S(\count7_1[5] ),
    .Y(_09057_));
 sky130_fd_sc_hd__mux4_2 _11590_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07150_));
 sky130_fd_sc_hd__mux4_2 _11591_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07151_));
 sky130_fd_sc_hd__mux4_2 _11592_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07152_));
 sky130_fd_sc_hd__mux4_2 _11593_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07153_));
 sky130_fd_sc_hd__mux4_2 _11594_ (.A0(_07150_),
    .A1(_07151_),
    .A2(_07152_),
    .A3(_07153_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07154_));
 sky130_fd_sc_hd__mux4_2 _11595_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07155_));
 sky130_fd_sc_hd__mux4_2 _11596_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07156_));
 sky130_fd_sc_hd__mux4_2 _11597_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07157_));
 sky130_fd_sc_hd__mux4_2 _11598_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07158_));
 sky130_fd_sc_hd__mux4_2 _11599_ (.A0(_07155_),
    .A1(_07156_),
    .A2(_07157_),
    .A3(_07158_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07159_));
 sky130_fd_sc_hd__mux2_2 _11600_ (.A0(_07154_),
    .A1(_07159_),
    .S(\count16_1[5] ),
    .X(_09062_));
 sky130_fd_sc_hd__mux4_2 _11601_ (.A0(\w[1][30] ),
    .A1(\w[3][30] ),
    .A2(\w[5][30] ),
    .A3(\w[7][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07160_));
 sky130_fd_sc_hd__mux4_2 _11602_ (.A0(\w[9][30] ),
    .A1(\w[11][30] ),
    .A2(\w[13][30] ),
    .A3(\w[15][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07161_));
 sky130_fd_sc_hd__mux4_2 _11603_ (.A0(\w[17][30] ),
    .A1(\w[19][30] ),
    .A2(\w[21][30] ),
    .A3(\w[23][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07162_));
 sky130_fd_sc_hd__mux4_2 _11604_ (.A0(\w[25][30] ),
    .A1(\w[27][30] ),
    .A2(\w[29][30] ),
    .A3(\w[31][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07163_));
 sky130_fd_sc_hd__mux4_2 _11605_ (.A0(_07160_),
    .A1(_07161_),
    .A2(_07162_),
    .A3(_07163_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07164_));
 sky130_fd_sc_hd__mux4_2 _11606_ (.A0(\w[33][30] ),
    .A1(\w[35][30] ),
    .A2(\w[37][30] ),
    .A3(\w[39][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07165_));
 sky130_fd_sc_hd__mux4_2 _11607_ (.A0(\w[41][30] ),
    .A1(\w[43][30] ),
    .A2(\w[45][30] ),
    .A3(\w[47][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07166_));
 sky130_fd_sc_hd__mux4_2 _11608_ (.A0(\w[49][30] ),
    .A1(\w[51][30] ),
    .A2(\w[53][30] ),
    .A3(\w[55][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07167_));
 sky130_fd_sc_hd__mux4_2 _11609_ (.A0(\w[57][30] ),
    .A1(\w[59][30] ),
    .A2(\w[61][30] ),
    .A3(\w[63][30] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07168_));
 sky130_fd_sc_hd__mux4_2 _11610_ (.A0(_07165_),
    .A1(_07166_),
    .A2(_07167_),
    .A3(_07168_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07169_));
 sky130_fd_sc_hd__mux2i_1 _11611_ (.A0(_07164_),
    .A1(_07169_),
    .S(\count7_1[5] ),
    .Y(_09065_));
 sky130_fd_sc_hd__mux4_2 _11619_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07177_));
 sky130_fd_sc_hd__mux4_2 _11624_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07182_));
 sky130_fd_sc_hd__mux4_2 _11627_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07185_));
 sky130_fd_sc_hd__mux4_2 _11631_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07189_));
 sky130_fd_sc_hd__mux4_2 _11637_ (.A0(_07177_),
    .A1(_07182_),
    .A2(_07185_),
    .A3(_07189_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07195_));
 sky130_fd_sc_hd__mux4_2 _11640_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07198_));
 sky130_fd_sc_hd__mux4_2 _11643_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07201_));
 sky130_fd_sc_hd__mux4_2 _11646_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07204_));
 sky130_fd_sc_hd__mux4_2 _11649_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07207_));
 sky130_fd_sc_hd__mux4_2 _11652_ (.A0(_07198_),
    .A1(_07201_),
    .A2(_07204_),
    .A3(_07207_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07210_));
 sky130_fd_sc_hd__mux2i_1 _11655_ (.A0(_07195_),
    .A1(_07210_),
    .S(\count7_2[5] ),
    .Y(_09071_));
 sky130_fd_sc_hd__mux4_2 _11656_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07213_));
 sky130_fd_sc_hd__mux4_2 _11657_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07214_));
 sky130_fd_sc_hd__mux4_2 _11659_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07216_));
 sky130_fd_sc_hd__mux4_2 _11660_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07217_));
 sky130_fd_sc_hd__mux4_2 _11661_ (.A0(_07213_),
    .A1(_07214_),
    .A2(_07216_),
    .A3(_07217_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07218_));
 sky130_fd_sc_hd__mux4_2 _11662_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07219_));
 sky130_fd_sc_hd__mux4_2 _11663_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07220_));
 sky130_fd_sc_hd__mux4_2 _11664_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07221_));
 sky130_fd_sc_hd__mux4_2 _11666_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07223_));
 sky130_fd_sc_hd__mux4_2 _11667_ (.A0(_07219_),
    .A1(_07220_),
    .A2(_07221_),
    .A3(_07223_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07224_));
 sky130_fd_sc_hd__mux2i_1 _11668_ (.A0(_07218_),
    .A1(_07224_),
    .S(\count7_2[5] ),
    .Y(_09076_));
 sky130_fd_sc_hd__mux4_2 _11669_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07225_));
 sky130_fd_sc_hd__mux4_2 _11670_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07226_));
 sky130_fd_sc_hd__mux4_2 _11672_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07228_));
 sky130_fd_sc_hd__mux4_2 _11673_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07229_));
 sky130_fd_sc_hd__mux4_2 _11674_ (.A0(_07225_),
    .A1(_07226_),
    .A2(_07228_),
    .A3(_07229_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07230_));
 sky130_fd_sc_hd__mux4_2 _11676_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07232_));
 sky130_fd_sc_hd__mux4_2 _11677_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07233_));
 sky130_fd_sc_hd__mux4_2 _11678_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07234_));
 sky130_fd_sc_hd__mux4_2 _11679_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07235_));
 sky130_fd_sc_hd__mux4_2 _11680_ (.A0(_07232_),
    .A1(_07233_),
    .A2(_07234_),
    .A3(_07235_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07236_));
 sky130_fd_sc_hd__mux2i_1 _11681_ (.A0(_07230_),
    .A1(_07236_),
    .S(\count7_2[5] ),
    .Y(_09085_));
 sky130_fd_sc_hd__mux4_2 _11682_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07237_));
 sky130_fd_sc_hd__mux4_2 _11683_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07238_));
 sky130_fd_sc_hd__mux4_2 _11684_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07239_));
 sky130_fd_sc_hd__mux4_2 _11685_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07240_));
 sky130_fd_sc_hd__mux4_2 _11686_ (.A0(_07237_),
    .A1(_07238_),
    .A2(_07239_),
    .A3(_07240_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07241_));
 sky130_fd_sc_hd__mux4_2 _11688_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07243_));
 sky130_fd_sc_hd__mux4_2 _11689_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07244_));
 sky130_fd_sc_hd__mux4_2 _11691_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07246_));
 sky130_fd_sc_hd__mux4_2 _11692_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07247_));
 sky130_fd_sc_hd__mux4_2 _11693_ (.A0(_07243_),
    .A1(_07244_),
    .A2(_07246_),
    .A3(_07247_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07248_));
 sky130_fd_sc_hd__mux2i_1 _11694_ (.A0(_07241_),
    .A1(_07248_),
    .S(\count7_2[5] ),
    .Y(_09097_));
 sky130_fd_sc_hd__mux4_2 _11695_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07249_));
 sky130_fd_sc_hd__mux4_2 _11697_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07251_));
 sky130_fd_sc_hd__mux4_2 _11698_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07252_));
 sky130_fd_sc_hd__mux4_2 _11699_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07253_));
 sky130_fd_sc_hd__mux4_2 _11700_ (.A0(_07249_),
    .A1(_07251_),
    .A2(_07252_),
    .A3(_07253_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07254_));
 sky130_fd_sc_hd__mux4_2 _11701_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07255_));
 sky130_fd_sc_hd__mux4_2 _11702_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07256_));
 sky130_fd_sc_hd__mux4_2 _11704_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07258_));
 sky130_fd_sc_hd__mux4_2 _11705_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07259_));
 sky130_fd_sc_hd__mux4_2 _11706_ (.A0(_07255_),
    .A1(_07256_),
    .A2(_07258_),
    .A3(_07259_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07260_));
 sky130_fd_sc_hd__mux2i_1 _11707_ (.A0(_07254_),
    .A1(_07260_),
    .S(\count7_2[5] ),
    .Y(_09106_));
 sky130_fd_sc_hd__mux4_2 _11708_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07261_));
 sky130_fd_sc_hd__mux4_2 _11710_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07263_));
 sky130_fd_sc_hd__mux4_2 _11711_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07264_));
 sky130_fd_sc_hd__mux4_2 _11712_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07265_));
 sky130_fd_sc_hd__mux4_2 _11713_ (.A0(_07261_),
    .A1(_07263_),
    .A2(_07264_),
    .A3(_07265_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07266_));
 sky130_fd_sc_hd__mux4_2 _11714_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07267_));
 sky130_fd_sc_hd__mux4_2 _11716_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07269_));
 sky130_fd_sc_hd__mux4_2 _11717_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07270_));
 sky130_fd_sc_hd__mux4_2 _11718_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07271_));
 sky130_fd_sc_hd__mux4_2 _11719_ (.A0(_07267_),
    .A1(_07269_),
    .A2(_07270_),
    .A3(_07271_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07272_));
 sky130_fd_sc_hd__mux2i_1 _11720_ (.A0(_07266_),
    .A1(_07272_),
    .S(\count7_2[5] ),
    .Y(_09115_));
 sky130_fd_sc_hd__mux4_2 _11721_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07273_));
 sky130_fd_sc_hd__mux4_2 _11722_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07274_));
 sky130_fd_sc_hd__mux4_2 _11723_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07275_));
 sky130_fd_sc_hd__mux4_2 _11724_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07276_));
 sky130_fd_sc_hd__mux4_2 _11725_ (.A0(_07273_),
    .A1(_07274_),
    .A2(_07275_),
    .A3(_07276_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07277_));
 sky130_fd_sc_hd__mux4_2 _11726_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07278_));
 sky130_fd_sc_hd__mux4_2 _11728_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07280_));
 sky130_fd_sc_hd__mux4_2 _11729_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07281_));
 sky130_fd_sc_hd__mux4_2 _11730_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07282_));
 sky130_fd_sc_hd__mux4_2 _11731_ (.A0(_07278_),
    .A1(_07280_),
    .A2(_07281_),
    .A3(_07282_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07283_));
 sky130_fd_sc_hd__mux2i_1 _11732_ (.A0(_07277_),
    .A1(_07283_),
    .S(\count7_2[5] ),
    .Y(_09124_));
 sky130_fd_sc_hd__mux4_2 _11733_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07284_));
 sky130_fd_sc_hd__mux4_2 _11734_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07285_));
 sky130_fd_sc_hd__mux4_2 _11735_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07286_));
 sky130_fd_sc_hd__mux4_2 _11736_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07287_));
 sky130_fd_sc_hd__mux4_2 _11738_ (.A0(_07284_),
    .A1(_07285_),
    .A2(_07286_),
    .A3(_07287_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07289_));
 sky130_fd_sc_hd__mux4_2 _11739_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07290_));
 sky130_fd_sc_hd__mux4_2 _11740_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07291_));
 sky130_fd_sc_hd__mux4_2 _11741_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07292_));
 sky130_fd_sc_hd__mux4_2 _11742_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07293_));
 sky130_fd_sc_hd__mux4_2 _11743_ (.A0(_07290_),
    .A1(_07291_),
    .A2(_07292_),
    .A3(_07293_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07294_));
 sky130_fd_sc_hd__mux2i_1 _11744_ (.A0(_07289_),
    .A1(_07294_),
    .S(\count7_2[5] ),
    .Y(_09133_));
 sky130_fd_sc_hd__mux4_2 _11745_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07295_));
 sky130_fd_sc_hd__mux4_2 _11746_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07296_));
 sky130_fd_sc_hd__mux4_2 _11747_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07297_));
 sky130_fd_sc_hd__mux4_2 _11749_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07299_));
 sky130_fd_sc_hd__mux4_2 _11751_ (.A0(_07295_),
    .A1(_07296_),
    .A2(_07297_),
    .A3(_07299_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07301_));
 sky130_fd_sc_hd__mux4_2 _11752_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07302_));
 sky130_fd_sc_hd__mux4_2 _11753_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07303_));
 sky130_fd_sc_hd__mux4_2 _11754_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07304_));
 sky130_fd_sc_hd__mux4_2 _11755_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07305_));
 sky130_fd_sc_hd__mux4_2 _11757_ (.A0(_07302_),
    .A1(_07303_),
    .A2(_07304_),
    .A3(_07305_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07307_));
 sky130_fd_sc_hd__mux2i_1 _11758_ (.A0(_07301_),
    .A1(_07307_),
    .S(\count7_2[5] ),
    .Y(_09142_));
 sky130_fd_sc_hd__mux4_2 _11760_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07309_));
 sky130_fd_sc_hd__mux4_2 _11761_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07310_));
 sky130_fd_sc_hd__mux4_2 _11762_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07311_));
 sky130_fd_sc_hd__mux4_2 _11764_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07313_));
 sky130_fd_sc_hd__mux4_2 _11765_ (.A0(_07309_),
    .A1(_07310_),
    .A2(_07311_),
    .A3(_07313_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07314_));
 sky130_fd_sc_hd__mux4_2 _11766_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07315_));
 sky130_fd_sc_hd__mux4_2 _11767_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07316_));
 sky130_fd_sc_hd__mux4_2 _11768_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07317_));
 sky130_fd_sc_hd__mux4_2 _11769_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07318_));
 sky130_fd_sc_hd__mux4_2 _11771_ (.A0(_07315_),
    .A1(_07316_),
    .A2(_07317_),
    .A3(_07318_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07320_));
 sky130_fd_sc_hd__mux2i_1 _11772_ (.A0(_07314_),
    .A1(_07320_),
    .S(\count7_2[5] ),
    .Y(_09151_));
 sky130_fd_sc_hd__mux4_2 _11774_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07322_));
 sky130_fd_sc_hd__mux4_2 _11775_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07323_));
 sky130_fd_sc_hd__mux4_2 _11776_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07324_));
 sky130_fd_sc_hd__mux4_2 _11777_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07325_));
 sky130_fd_sc_hd__mux4_2 _11778_ (.A0(_07322_),
    .A1(_07323_),
    .A2(_07324_),
    .A3(_07325_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07326_));
 sky130_fd_sc_hd__mux4_2 _11779_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07327_));
 sky130_fd_sc_hd__mux4_2 _11780_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07328_));
 sky130_fd_sc_hd__mux4_2 _11781_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07329_));
 sky130_fd_sc_hd__mux4_2 _11783_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07331_));
 sky130_fd_sc_hd__mux4_2 _11784_ (.A0(_07327_),
    .A1(_07328_),
    .A2(_07329_),
    .A3(_07331_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07332_));
 sky130_fd_sc_hd__mux2i_1 _11786_ (.A0(_07326_),
    .A1(_07332_),
    .S(\count7_2[5] ),
    .Y(_09160_));
 sky130_fd_sc_hd__mux4_2 _11787_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07334_));
 sky130_fd_sc_hd__mux4_2 _11788_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07335_));
 sky130_fd_sc_hd__mux4_2 _11790_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07337_));
 sky130_fd_sc_hd__mux4_2 _11791_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07338_));
 sky130_fd_sc_hd__mux4_2 _11792_ (.A0(_07334_),
    .A1(_07335_),
    .A2(_07337_),
    .A3(_07338_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07339_));
 sky130_fd_sc_hd__mux4_2 _11793_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07340_));
 sky130_fd_sc_hd__mux4_2 _11794_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07341_));
 sky130_fd_sc_hd__mux4_2 _11795_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07342_));
 sky130_fd_sc_hd__mux4_2 _11797_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07344_));
 sky130_fd_sc_hd__mux4_2 _11798_ (.A0(_07340_),
    .A1(_07341_),
    .A2(_07342_),
    .A3(_07344_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07345_));
 sky130_fd_sc_hd__mux2i_1 _11799_ (.A0(_07339_),
    .A1(_07345_),
    .S(\count7_2[5] ),
    .Y(_09169_));
 sky130_fd_sc_hd__mux4_2 _11800_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07346_));
 sky130_fd_sc_hd__mux4_2 _11801_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07347_));
 sky130_fd_sc_hd__mux4_2 _11803_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07349_));
 sky130_fd_sc_hd__mux4_2 _11804_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07350_));
 sky130_fd_sc_hd__mux4_2 _11805_ (.A0(_07346_),
    .A1(_07347_),
    .A2(_07349_),
    .A3(_07350_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07351_));
 sky130_fd_sc_hd__mux4_2 _11807_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07353_));
 sky130_fd_sc_hd__mux4_2 _11808_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07354_));
 sky130_fd_sc_hd__mux4_2 _11809_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07355_));
 sky130_fd_sc_hd__mux4_2 _11810_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07356_));
 sky130_fd_sc_hd__mux4_2 _11811_ (.A0(_07353_),
    .A1(_07354_),
    .A2(_07355_),
    .A3(_07356_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07357_));
 sky130_fd_sc_hd__mux2i_1 _11812_ (.A0(_07351_),
    .A1(_07357_),
    .S(\count7_2[5] ),
    .Y(_09178_));
 sky130_fd_sc_hd__mux4_2 _11813_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07358_));
 sky130_fd_sc_hd__mux4_2 _11814_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07359_));
 sky130_fd_sc_hd__mux4_2 _11815_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07360_));
 sky130_fd_sc_hd__mux4_2 _11816_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07361_));
 sky130_fd_sc_hd__mux4_2 _11817_ (.A0(_07358_),
    .A1(_07359_),
    .A2(_07360_),
    .A3(_07361_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07362_));
 sky130_fd_sc_hd__mux4_2 _11819_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07364_));
 sky130_fd_sc_hd__mux4_2 _11820_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07365_));
 sky130_fd_sc_hd__mux4_2 _11822_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07367_));
 sky130_fd_sc_hd__mux4_2 _11823_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07368_));
 sky130_fd_sc_hd__mux4_2 _11824_ (.A0(_07364_),
    .A1(_07365_),
    .A2(_07367_),
    .A3(_07368_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07369_));
 sky130_fd_sc_hd__mux2i_1 _11825_ (.A0(_07362_),
    .A1(_07369_),
    .S(\count7_2[5] ),
    .Y(_09187_));
 sky130_fd_sc_hd__mux4_2 _11826_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07370_));
 sky130_fd_sc_hd__mux4_2 _11828_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07372_));
 sky130_fd_sc_hd__mux4_2 _11829_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07373_));
 sky130_fd_sc_hd__mux4_2 _11830_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07374_));
 sky130_fd_sc_hd__mux4_2 _11831_ (.A0(_07370_),
    .A1(_07372_),
    .A2(_07373_),
    .A3(_07374_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07375_));
 sky130_fd_sc_hd__mux4_2 _11832_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07376_));
 sky130_fd_sc_hd__mux4_2 _11833_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07377_));
 sky130_fd_sc_hd__mux4_2 _11835_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07379_));
 sky130_fd_sc_hd__mux4_2 _11836_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07380_));
 sky130_fd_sc_hd__mux4_2 _11837_ (.A0(_07376_),
    .A1(_07377_),
    .A2(_07379_),
    .A3(_07380_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07381_));
 sky130_fd_sc_hd__mux2i_1 _11838_ (.A0(_07375_),
    .A1(_07381_),
    .S(\count7_2[5] ),
    .Y(_09196_));
 sky130_fd_sc_hd__mux4_2 _11839_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07382_));
 sky130_fd_sc_hd__mux4_2 _11841_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07384_));
 sky130_fd_sc_hd__mux4_2 _11842_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07385_));
 sky130_fd_sc_hd__mux4_2 _11843_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07386_));
 sky130_fd_sc_hd__mux4_2 _11844_ (.A0(_07382_),
    .A1(_07384_),
    .A2(_07385_),
    .A3(_07386_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07387_));
 sky130_fd_sc_hd__mux4_2 _11845_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07388_));
 sky130_fd_sc_hd__mux4_2 _11847_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07390_));
 sky130_fd_sc_hd__mux4_2 _11848_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07391_));
 sky130_fd_sc_hd__mux4_2 _11849_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07392_));
 sky130_fd_sc_hd__mux4_2 _11850_ (.A0(_07388_),
    .A1(_07390_),
    .A2(_07391_),
    .A3(_07392_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07393_));
 sky130_fd_sc_hd__mux2i_1 _11851_ (.A0(_07387_),
    .A1(_07393_),
    .S(\count7_2[5] ),
    .Y(_09205_));
 sky130_fd_sc_hd__mux4_2 _11852_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07394_));
 sky130_fd_sc_hd__mux4_2 _11853_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07395_));
 sky130_fd_sc_hd__mux4_2 _11854_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07396_));
 sky130_fd_sc_hd__mux4_2 _11855_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07397_));
 sky130_fd_sc_hd__mux4_2 _11856_ (.A0(_07394_),
    .A1(_07395_),
    .A2(_07396_),
    .A3(_07397_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07398_));
 sky130_fd_sc_hd__mux4_2 _11857_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07399_));
 sky130_fd_sc_hd__mux4_2 _11859_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07401_));
 sky130_fd_sc_hd__mux4_2 _11860_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07402_));
 sky130_fd_sc_hd__mux4_2 _11861_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07403_));
 sky130_fd_sc_hd__mux4_2 _11862_ (.A0(_07399_),
    .A1(_07401_),
    .A2(_07402_),
    .A3(_07403_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07404_));
 sky130_fd_sc_hd__mux2i_1 _11863_ (.A0(_07398_),
    .A1(_07404_),
    .S(\count7_2[5] ),
    .Y(_09214_));
 sky130_fd_sc_hd__mux4_2 _11864_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07405_));
 sky130_fd_sc_hd__mux4_2 _11865_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07406_));
 sky130_fd_sc_hd__mux4_2 _11866_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07407_));
 sky130_fd_sc_hd__mux4_2 _11867_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07408_));
 sky130_fd_sc_hd__mux4_2 _11869_ (.A0(_07405_),
    .A1(_07406_),
    .A2(_07407_),
    .A3(_07408_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07410_));
 sky130_fd_sc_hd__mux4_2 _11870_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07411_));
 sky130_fd_sc_hd__mux4_2 _11871_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07412_));
 sky130_fd_sc_hd__mux4_2 _11872_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07413_));
 sky130_fd_sc_hd__mux4_2 _11873_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07414_));
 sky130_fd_sc_hd__mux4_2 _11874_ (.A0(_07411_),
    .A1(_07412_),
    .A2(_07413_),
    .A3(_07414_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07415_));
 sky130_fd_sc_hd__mux2i_1 _11875_ (.A0(_07410_),
    .A1(_07415_),
    .S(\count7_2[5] ),
    .Y(_09223_));
 sky130_fd_sc_hd__mux4_2 _11876_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07416_));
 sky130_fd_sc_hd__mux4_2 _11877_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07417_));
 sky130_fd_sc_hd__mux4_2 _11878_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07418_));
 sky130_fd_sc_hd__mux4_2 _11880_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07420_));
 sky130_fd_sc_hd__mux4_2 _11882_ (.A0(_07416_),
    .A1(_07417_),
    .A2(_07418_),
    .A3(_07420_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07422_));
 sky130_fd_sc_hd__mux4_2 _11883_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07423_));
 sky130_fd_sc_hd__mux4_2 _11884_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07424_));
 sky130_fd_sc_hd__mux4_2 _11885_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07425_));
 sky130_fd_sc_hd__mux4_2 _11886_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07426_));
 sky130_fd_sc_hd__mux4_2 _11888_ (.A0(_07423_),
    .A1(_07424_),
    .A2(_07425_),
    .A3(_07426_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07428_));
 sky130_fd_sc_hd__mux2i_1 _11889_ (.A0(_07422_),
    .A1(_07428_),
    .S(\count7_2[5] ),
    .Y(_09232_));
 sky130_fd_sc_hd__mux4_2 _11891_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07430_));
 sky130_fd_sc_hd__mux4_2 _11892_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07431_));
 sky130_fd_sc_hd__mux4_2 _11893_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07432_));
 sky130_fd_sc_hd__mux4_2 _11895_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07434_));
 sky130_fd_sc_hd__mux4_2 _11896_ (.A0(_07430_),
    .A1(_07431_),
    .A2(_07432_),
    .A3(_07434_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07435_));
 sky130_fd_sc_hd__mux4_2 _11897_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07436_));
 sky130_fd_sc_hd__mux4_2 _11898_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07437_));
 sky130_fd_sc_hd__mux4_2 _11899_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07438_));
 sky130_fd_sc_hd__mux4_2 _11900_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07439_));
 sky130_fd_sc_hd__mux4_2 _11902_ (.A0(_07436_),
    .A1(_07437_),
    .A2(_07438_),
    .A3(_07439_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07441_));
 sky130_fd_sc_hd__mux2i_1 _11903_ (.A0(_07435_),
    .A1(_07441_),
    .S(\count7_2[5] ),
    .Y(_09241_));
 sky130_fd_sc_hd__mux4_2 _11904_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07442_));
 sky130_fd_sc_hd__mux4_2 _11905_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07443_));
 sky130_fd_sc_hd__mux4_2 _11906_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07444_));
 sky130_fd_sc_hd__mux4_2 _11907_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07445_));
 sky130_fd_sc_hd__mux4_2 _11908_ (.A0(_07442_),
    .A1(_07443_),
    .A2(_07444_),
    .A3(_07445_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07446_));
 sky130_fd_sc_hd__mux4_2 _11909_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07447_));
 sky130_fd_sc_hd__mux4_2 _11910_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07448_));
 sky130_fd_sc_hd__mux4_2 _11911_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07449_));
 sky130_fd_sc_hd__mux4_2 _11912_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07450_));
 sky130_fd_sc_hd__mux4_2 _11913_ (.A0(_07447_),
    .A1(_07448_),
    .A2(_07449_),
    .A3(_07450_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07451_));
 sky130_fd_sc_hd__mux2i_1 _11915_ (.A0(_07446_),
    .A1(_07451_),
    .S(\count7_2[5] ),
    .Y(_09250_));
 sky130_fd_sc_hd__mux4_2 _11916_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07453_));
 sky130_fd_sc_hd__mux4_2 _11917_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07454_));
 sky130_fd_sc_hd__mux4_2 _11918_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07455_));
 sky130_fd_sc_hd__mux4_2 _11919_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07456_));
 sky130_fd_sc_hd__mux4_2 _11920_ (.A0(_07453_),
    .A1(_07454_),
    .A2(_07455_),
    .A3(_07456_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07457_));
 sky130_fd_sc_hd__mux4_2 _11921_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07458_));
 sky130_fd_sc_hd__mux4_2 _11922_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07459_));
 sky130_fd_sc_hd__mux4_2 _11923_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07460_));
 sky130_fd_sc_hd__mux4_2 _11924_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07461_));
 sky130_fd_sc_hd__mux4_2 _11925_ (.A0(_07458_),
    .A1(_07459_),
    .A2(_07460_),
    .A3(_07461_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07462_));
 sky130_fd_sc_hd__mux2i_1 _11926_ (.A0(_07457_),
    .A1(_07462_),
    .S(\count7_2[5] ),
    .Y(_09259_));
 sky130_fd_sc_hd__mux4_2 _11927_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07463_));
 sky130_fd_sc_hd__mux4_2 _11928_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07464_));
 sky130_fd_sc_hd__mux4_2 _11929_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07465_));
 sky130_fd_sc_hd__mux4_2 _11930_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07466_));
 sky130_fd_sc_hd__mux4_2 _11931_ (.A0(_07463_),
    .A1(_07464_),
    .A2(_07465_),
    .A3(_07466_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07467_));
 sky130_fd_sc_hd__mux4_2 _11932_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07468_));
 sky130_fd_sc_hd__mux4_2 _11933_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07469_));
 sky130_fd_sc_hd__mux4_2 _11934_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07470_));
 sky130_fd_sc_hd__mux4_2 _11935_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07471_));
 sky130_fd_sc_hd__mux4_2 _11936_ (.A0(_07468_),
    .A1(_07469_),
    .A2(_07470_),
    .A3(_07471_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07472_));
 sky130_fd_sc_hd__mux2i_1 _11937_ (.A0(_07467_),
    .A1(_07472_),
    .S(\count7_2[5] ),
    .Y(_09268_));
 sky130_fd_sc_hd__mux4_2 _11938_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07473_));
 sky130_fd_sc_hd__mux4_2 _11939_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07474_));
 sky130_fd_sc_hd__mux4_2 _11940_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07475_));
 sky130_fd_sc_hd__mux4_2 _11941_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07476_));
 sky130_fd_sc_hd__mux4_2 _11942_ (.A0(_07473_),
    .A1(_07474_),
    .A2(_07475_),
    .A3(_07476_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07477_));
 sky130_fd_sc_hd__mux4_2 _11943_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07478_));
 sky130_fd_sc_hd__mux4_2 _11944_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07479_));
 sky130_fd_sc_hd__mux4_2 _11945_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07480_));
 sky130_fd_sc_hd__mux4_2 _11946_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07481_));
 sky130_fd_sc_hd__mux4_2 _11947_ (.A0(_07478_),
    .A1(_07479_),
    .A2(_07480_),
    .A3(_07481_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07482_));
 sky130_fd_sc_hd__mux2i_1 _11948_ (.A0(_07477_),
    .A1(_07482_),
    .S(\count7_2[5] ),
    .Y(_09277_));
 sky130_fd_sc_hd__mux4_2 _11949_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07483_));
 sky130_fd_sc_hd__mux4_2 _11950_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07484_));
 sky130_fd_sc_hd__mux4_2 _11951_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07485_));
 sky130_fd_sc_hd__mux4_2 _11952_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07486_));
 sky130_fd_sc_hd__mux4_2 _11953_ (.A0(_07483_),
    .A1(_07484_),
    .A2(_07485_),
    .A3(_07486_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07487_));
 sky130_fd_sc_hd__mux4_2 _11954_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07488_));
 sky130_fd_sc_hd__mux4_2 _11955_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07489_));
 sky130_fd_sc_hd__mux4_2 _11956_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07490_));
 sky130_fd_sc_hd__mux4_2 _11957_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07491_));
 sky130_fd_sc_hd__mux4_2 _11958_ (.A0(_07488_),
    .A1(_07489_),
    .A2(_07490_),
    .A3(_07491_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07492_));
 sky130_fd_sc_hd__mux2i_1 _11959_ (.A0(_07487_),
    .A1(_07492_),
    .S(\count7_2[5] ),
    .Y(_09286_));
 sky130_fd_sc_hd__mux4_2 _11960_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07493_));
 sky130_fd_sc_hd__mux4_2 _11961_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07494_));
 sky130_fd_sc_hd__mux4_2 _11962_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07495_));
 sky130_fd_sc_hd__mux4_2 _11963_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07496_));
 sky130_fd_sc_hd__mux4_2 _11964_ (.A0(_07493_),
    .A1(_07494_),
    .A2(_07495_),
    .A3(_07496_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07497_));
 sky130_fd_sc_hd__mux4_2 _11965_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07498_));
 sky130_fd_sc_hd__mux4_2 _11967_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07500_));
 sky130_fd_sc_hd__mux4_2 _11968_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07501_));
 sky130_fd_sc_hd__mux4_2 _11969_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07502_));
 sky130_fd_sc_hd__mux4_2 _11970_ (.A0(_07498_),
    .A1(_07500_),
    .A2(_07501_),
    .A3(_07502_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07503_));
 sky130_fd_sc_hd__mux2i_1 _11971_ (.A0(_07497_),
    .A1(_07503_),
    .S(\count7_2[5] ),
    .Y(_09295_));
 sky130_fd_sc_hd__mux4_2 _11972_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07504_));
 sky130_fd_sc_hd__mux4_2 _11973_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07505_));
 sky130_fd_sc_hd__mux4_2 _11974_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07506_));
 sky130_fd_sc_hd__mux4_2 _11975_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07507_));
 sky130_fd_sc_hd__mux4_2 _11976_ (.A0(_07504_),
    .A1(_07505_),
    .A2(_07506_),
    .A3(_07507_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07508_));
 sky130_fd_sc_hd__mux4_2 _11977_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07509_));
 sky130_fd_sc_hd__mux4_2 _11979_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07511_));
 sky130_fd_sc_hd__mux4_2 _11980_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07512_));
 sky130_fd_sc_hd__mux4_2 _11981_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07513_));
 sky130_fd_sc_hd__mux4_2 _11982_ (.A0(_07509_),
    .A1(_07511_),
    .A2(_07512_),
    .A3(_07513_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07514_));
 sky130_fd_sc_hd__mux2i_1 _11983_ (.A0(_07508_),
    .A1(_07514_),
    .S(\count7_2[5] ),
    .Y(_09304_));
 sky130_fd_sc_hd__mux4_2 _11984_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07515_));
 sky130_fd_sc_hd__mux4_2 _11985_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07516_));
 sky130_fd_sc_hd__mux4_2 _11986_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07517_));
 sky130_fd_sc_hd__mux4_2 _11987_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07518_));
 sky130_fd_sc_hd__mux4_2 _11988_ (.A0(_07515_),
    .A1(_07516_),
    .A2(_07517_),
    .A3(_07518_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07519_));
 sky130_fd_sc_hd__mux4_2 _11989_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07520_));
 sky130_fd_sc_hd__mux4_2 _11990_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07521_));
 sky130_fd_sc_hd__mux4_2 _11991_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07522_));
 sky130_fd_sc_hd__mux4_2 _11992_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07523_));
 sky130_fd_sc_hd__mux4_2 _11993_ (.A0(_07520_),
    .A1(_07521_),
    .A2(_07522_),
    .A3(_07523_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07524_));
 sky130_fd_sc_hd__mux2i_1 _11994_ (.A0(_07519_),
    .A1(_07524_),
    .S(\count7_2[5] ),
    .Y(_09313_));
 sky130_fd_sc_hd__mux4_2 _12000_ (.A0(\w[1][28] ),
    .A1(\w[3][28] ),
    .A2(\w[5][28] ),
    .A3(\w[7][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07530_));
 sky130_fd_sc_hd__mux4_2 _12002_ (.A0(\w[9][28] ),
    .A1(\w[11][28] ),
    .A2(\w[13][28] ),
    .A3(\w[15][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07532_));
 sky130_fd_sc_hd__mux4_2 _12003_ (.A0(\w[17][28] ),
    .A1(\w[19][28] ),
    .A2(\w[21][28] ),
    .A3(\w[23][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07533_));
 sky130_fd_sc_hd__mux4_2 _12005_ (.A0(\w[25][28] ),
    .A1(\w[27][28] ),
    .A2(\w[29][28] ),
    .A3(\w[31][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07535_));
 sky130_fd_sc_hd__mux4_2 _12009_ (.A0(_07530_),
    .A1(_07532_),
    .A2(_07533_),
    .A3(_07535_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_07539_));
 sky130_fd_sc_hd__mux4_2 _12010_ (.A0(\w[33][28] ),
    .A1(\w[35][28] ),
    .A2(\w[37][28] ),
    .A3(\w[39][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07540_));
 sky130_fd_sc_hd__mux4_2 _12011_ (.A0(\w[41][28] ),
    .A1(\w[43][28] ),
    .A2(\w[45][28] ),
    .A3(\w[47][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07541_));
 sky130_fd_sc_hd__mux4_2 _12012_ (.A0(\w[49][28] ),
    .A1(\w[51][28] ),
    .A2(\w[53][28] ),
    .A3(\w[55][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07542_));
 sky130_fd_sc_hd__mux4_2 _12013_ (.A0(\w[57][28] ),
    .A1(\w[59][28] ),
    .A2(\w[61][28] ),
    .A3(\w[63][28] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07543_));
 sky130_fd_sc_hd__mux4_2 _12014_ (.A0(_07540_),
    .A1(_07541_),
    .A2(_07542_),
    .A3(_07543_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_07544_));
 sky130_fd_sc_hd__mux2_2 _12016_ (.A0(_07539_),
    .A1(_07544_),
    .S(\count16_2[5] ),
    .X(_09322_));
 sky130_fd_sc_hd__mux4_2 _12017_ (.A0(\w[1][29] ),
    .A1(\w[3][29] ),
    .A2(\w[5][29] ),
    .A3(\w[7][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07546_));
 sky130_fd_sc_hd__mux4_2 _12018_ (.A0(\w[9][29] ),
    .A1(\w[11][29] ),
    .A2(\w[13][29] ),
    .A3(\w[15][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07547_));
 sky130_fd_sc_hd__mux4_2 _12019_ (.A0(\w[17][29] ),
    .A1(\w[19][29] ),
    .A2(\w[21][29] ),
    .A3(\w[23][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07548_));
 sky130_fd_sc_hd__mux4_2 _12020_ (.A0(\w[25][29] ),
    .A1(\w[27][29] ),
    .A2(\w[29][29] ),
    .A3(\w[31][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07549_));
 sky130_fd_sc_hd__mux4_2 _12021_ (.A0(_07546_),
    .A1(_07547_),
    .A2(_07548_),
    .A3(_07549_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_07550_));
 sky130_fd_sc_hd__mux4_2 _12022_ (.A0(\w[33][29] ),
    .A1(\w[35][29] ),
    .A2(\w[37][29] ),
    .A3(\w[39][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07551_));
 sky130_fd_sc_hd__mux4_2 _12023_ (.A0(\w[41][29] ),
    .A1(\w[43][29] ),
    .A2(\w[45][29] ),
    .A3(\w[47][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07552_));
 sky130_fd_sc_hd__mux4_2 _12024_ (.A0(\w[49][29] ),
    .A1(\w[51][29] ),
    .A2(\w[53][29] ),
    .A3(\w[55][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07553_));
 sky130_fd_sc_hd__mux4_2 _12025_ (.A0(\w[57][29] ),
    .A1(\w[59][29] ),
    .A2(\w[61][29] ),
    .A3(\w[63][29] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_07554_));
 sky130_fd_sc_hd__mux4_2 _12026_ (.A0(_07551_),
    .A1(_07552_),
    .A2(_07553_),
    .A3(_07554_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_07555_));
 sky130_fd_sc_hd__mux2_2 _12027_ (.A0(_07550_),
    .A1(_07555_),
    .S(\count16_2[5] ),
    .X(_09330_));
 sky130_fd_sc_hd__mux4_2 _12028_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07556_));
 sky130_fd_sc_hd__mux4_2 _12029_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07557_));
 sky130_fd_sc_hd__mux4_2 _12030_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07558_));
 sky130_fd_sc_hd__mux4_2 _12031_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07559_));
 sky130_fd_sc_hd__mux4_2 _12032_ (.A0(_07556_),
    .A1(_07557_),
    .A2(_07558_),
    .A3(_07559_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07560_));
 sky130_fd_sc_hd__mux4_2 _12033_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07561_));
 sky130_fd_sc_hd__mux4_2 _12034_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07562_));
 sky130_fd_sc_hd__mux4_2 _12035_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07563_));
 sky130_fd_sc_hd__mux4_2 _12036_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_07564_));
 sky130_fd_sc_hd__mux4_2 _12037_ (.A0(_07561_),
    .A1(_07562_),
    .A2(_07563_),
    .A3(_07564_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_07565_));
 sky130_fd_sc_hd__mux2i_1 _12038_ (.A0(_07560_),
    .A1(_07565_),
    .S(\count7_2[5] ),
    .Y(_09339_));
 sky130_fd_sc_hd__nor2b_1 _12039_ (.A(reset),
    .B_N(_09554_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_1 _12041_ (.A(_05338_),
    .B(_07566_),
    .Y(_07568_));
 sky130_fd_sc_hd__mux2i_2 _12045_ (.A0(_09370_),
    .A1(\w[62][0] ),
    .S(done),
    .Y(_07572_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(message[31]),
    .B(_07568_),
    .Y(_07576_));
 sky130_fd_sc_hd__o21ai_0 _12050_ (.A1(_07568_),
    .A2(_07572_),
    .B1(_07576_),
    .Y(_00129_));
 sky130_fd_sc_hd__mux2i_2 _12051_ (.A0(_09372_),
    .A1(\w[62][1] ),
    .S(done),
    .Y(_07577_));
 sky130_fd_sc_hd__nand2_1 _12053_ (.A(message[30]),
    .B(_07568_),
    .Y(_07579_));
 sky130_fd_sc_hd__o21ai_0 _12054_ (.A1(_07568_),
    .A2(_07577_),
    .B1(_07579_),
    .Y(_00140_));
 sky130_fd_sc_hd__mux2i_2 _12056_ (.A0(_08845_),
    .A1(\w[62][2] ),
    .S(done),
    .Y(_07581_));
 sky130_fd_sc_hd__nand2_1 _12058_ (.A(message[29]),
    .B(_07568_),
    .Y(_07583_));
 sky130_fd_sc_hd__o21ai_0 _12059_ (.A1(_07568_),
    .A2(_07581_),
    .B1(_07583_),
    .Y(_00151_));
 sky130_fd_sc_hd__xnor2_1 _12062_ (.A(_08844_),
    .B(_09378_),
    .Y(_07586_));
 sky130_fd_sc_hd__nor2_1 _12063_ (.A(done),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__a21oi_1 _12064_ (.A1(\w[62][3] ),
    .A2(done),
    .B1(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__nand2_1 _12066_ (.A(message[28]),
    .B(_07568_),
    .Y(_07590_));
 sky130_fd_sc_hd__o21ai_0 _12067_ (.A1(_07568_),
    .A2(_07588_),
    .B1(_07590_),
    .Y(_00154_));
 sky130_fd_sc_hd__inv_2 _12068_ (.A(done),
    .Y(_07591_));
 sky130_fd_sc_hd__a21o_1 _12071_ (.A1(_08841_),
    .A2(_09374_),
    .B1(_09373_),
    .X(_07594_));
 sky130_fd_sc_hd__a211oi_1 _12072_ (.A1(_09378_),
    .A2(_07594_),
    .B1(_09377_),
    .C1(_09382_),
    .Y(_07595_));
 sky130_fd_sc_hd__a211oi_1 _12073_ (.A1(_08841_),
    .A2(_09374_),
    .B1(_09373_),
    .C1(_09377_),
    .Y(_07596_));
 sky130_fd_sc_hd__o21ai_0 _12074_ (.A1(_09378_),
    .A2(_09377_),
    .B1(_09382_),
    .Y(_07597_));
 sky130_fd_sc_hd__nor2_1 _12075_ (.A(_07596_),
    .B(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__o21ai_0 _12077_ (.A1(_07595_),
    .A2(_07598_),
    .B1(_07591_),
    .Y(_07600_));
 sky130_fd_sc_hd__o21ai_1 _12078_ (.A1(\w[62][4] ),
    .A2(_07591_),
    .B1(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__nand2_1 _12080_ (.A(message[27]),
    .B(_07568_),
    .Y(_07603_));
 sky130_fd_sc_hd__o21ai_0 _12081_ (.A1(_07568_),
    .A2(_07601_),
    .B1(_07603_),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_1 _12083_ (.A(_09390_),
    .Y(_07605_));
 sky130_fd_sc_hd__a21o_1 _12084_ (.A1(_08844_),
    .A2(_09378_),
    .B1(_09377_),
    .X(_07606_));
 sky130_fd_sc_hd__a21oi_1 _12085_ (.A1(_09382_),
    .A2(_07606_),
    .B1(_09381_),
    .Y(_07607_));
 sky130_fd_sc_hd__xnor2_1 _12086_ (.A(_07605_),
    .B(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__nand2_1 _12087_ (.A(_07591_),
    .B(_07608_),
    .Y(_07609_));
 sky130_fd_sc_hd__o21ai_1 _12088_ (.A1(\w[62][5] ),
    .A2(_07591_),
    .B1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__nand2_1 _12090_ (.A(message[26]),
    .B(_07568_),
    .Y(_07612_));
 sky130_fd_sc_hd__o21ai_0 _12091_ (.A1(_07568_),
    .A2(_07610_),
    .B1(_07612_),
    .Y(_00156_));
 sky130_fd_sc_hd__nor2_1 _12092_ (.A(_09381_),
    .B(_09389_),
    .Y(_07613_));
 sky130_fd_sc_hd__o21ai_0 _12093_ (.A1(_07596_),
    .A2(_07597_),
    .B1(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__o21a_1 _12094_ (.A1(_09390_),
    .A2(_09389_),
    .B1(_09386_),
    .X(_07615_));
 sky130_fd_sc_hd__nor2_1 _12095_ (.A(_09386_),
    .B(_09389_),
    .Y(_07616_));
 sky130_fd_sc_hd__o21ai_0 _12096_ (.A1(_09381_),
    .A2(_07598_),
    .B1(_09390_),
    .Y(_07617_));
 sky130_fd_sc_hd__a221oi_1 _12098_ (.A1(_07614_),
    .A2(_07615_),
    .B1(_07616_),
    .B2(_07617_),
    .C1(done),
    .Y(_07619_));
 sky130_fd_sc_hd__a21oi_1 _12099_ (.A1(\w[62][6] ),
    .A2(done),
    .B1(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__nand2_1 _12101_ (.A(message[25]),
    .B(_07568_),
    .Y(_07622_));
 sky130_fd_sc_hd__o21ai_0 _12102_ (.A1(_07568_),
    .A2(_07620_),
    .B1(_07622_),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_1 _12103_ (.A(_09394_),
    .Y(_07623_));
 sky130_fd_sc_hd__o21bai_1 _12104_ (.A1(_07605_),
    .A2(_07607_),
    .B1_N(_09389_),
    .Y(_07624_));
 sky130_fd_sc_hd__a21oi_1 _12105_ (.A1(_09386_),
    .A2(_07624_),
    .B1(_09385_),
    .Y(_07625_));
 sky130_fd_sc_hd__xnor2_1 _12106_ (.A(_07623_),
    .B(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__nor2_1 _12107_ (.A(done),
    .B(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__a21oi_1 _12108_ (.A1(\w[62][7] ),
    .A2(done),
    .B1(_07627_),
    .Y(_07628_));
 sky130_fd_sc_hd__nand2_1 _12110_ (.A(message[24]),
    .B(_07568_),
    .Y(_07630_));
 sky130_fd_sc_hd__o21ai_0 _12111_ (.A1(_07568_),
    .A2(_07628_),
    .B1(_07630_),
    .Y(_00158_));
 sky130_fd_sc_hd__a21oi_1 _12112_ (.A1(_07614_),
    .A2(_07615_),
    .B1(_09385_),
    .Y(_07631_));
 sky130_fd_sc_hd__o21bai_1 _12113_ (.A1(_07623_),
    .A2(_07631_),
    .B1_N(_09393_),
    .Y(_07632_));
 sky130_fd_sc_hd__xnor2_1 _12114_ (.A(_09398_),
    .B(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__nor2_1 _12115_ (.A(done),
    .B(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__a21oi_1 _12116_ (.A1(\w[62][8] ),
    .A2(done),
    .B1(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__nand2_1 _12118_ (.A(message[23]),
    .B(_07568_),
    .Y(_07637_));
 sky130_fd_sc_hd__o21ai_0 _12119_ (.A1(_07568_),
    .A2(_07635_),
    .B1(_07637_),
    .Y(_00159_));
 sky130_fd_sc_hd__o21a_1 _12120_ (.A1(_09386_),
    .A2(_09385_),
    .B1(_09394_),
    .X(_07638_));
 sky130_fd_sc_hd__o21ai_0 _12121_ (.A1(_09393_),
    .A2(_07638_),
    .B1(_09398_),
    .Y(_07639_));
 sky130_fd_sc_hd__nand2b_1 _12122_ (.A_N(_09397_),
    .B(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__a2111oi_0 _12123_ (.A1(_09398_),
    .A2(_09393_),
    .B1(_09397_),
    .C1(_09385_),
    .D1(_09389_),
    .Y(_07641_));
 sky130_fd_sc_hd__o21ai_1 _12124_ (.A1(_07605_),
    .A2(_07607_),
    .B1(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__nand2_1 _12125_ (.A(_07640_),
    .B(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__xor2_1 _12126_ (.A(_09402_),
    .B(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__nor2_1 _12127_ (.A(done),
    .B(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__a21oi_1 _12128_ (.A1(\w[62][9] ),
    .A2(done),
    .B1(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__nand2_1 _12130_ (.A(message[22]),
    .B(_07568_),
    .Y(_07648_));
 sky130_fd_sc_hd__o21ai_0 _12131_ (.A1(_07568_),
    .A2(_07646_),
    .B1(_07648_),
    .Y(_00160_));
 sky130_fd_sc_hd__a21oi_1 _12132_ (.A1(_09394_),
    .A2(_09385_),
    .B1(_09393_),
    .Y(_07649_));
 sky130_fd_sc_hd__nand2_1 _12133_ (.A(_09398_),
    .B(_09402_),
    .Y(_07650_));
 sky130_fd_sc_hd__a21oi_1 _12134_ (.A1(_09402_),
    .A2(_09397_),
    .B1(_09401_),
    .Y(_07651_));
 sky130_fd_sc_hd__o21a_1 _12135_ (.A1(_07649_),
    .A2(_07650_),
    .B1(_07651_),
    .X(_07652_));
 sky130_fd_sc_hd__nor2_1 _12136_ (.A(_07623_),
    .B(_07650_),
    .Y(_07653_));
 sky130_fd_sc_hd__nand3_1 _12137_ (.A(_07614_),
    .B(_07615_),
    .C(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__a21boi_0 _12138_ (.A1(_07652_),
    .A2(_07654_),
    .B1_N(_09406_),
    .Y(_07655_));
 sky130_fd_sc_hd__nand2_1 _12139_ (.A(_07652_),
    .B(_07654_),
    .Y(_07656_));
 sky130_fd_sc_hd__nor2_1 _12140_ (.A(_09406_),
    .B(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__o21ai_0 _12142_ (.A1(_07655_),
    .A2(_07657_),
    .B1(_07591_),
    .Y(_07659_));
 sky130_fd_sc_hd__o21ai_1 _12143_ (.A1(\w[62][10] ),
    .A2(_07591_),
    .B1(_07659_),
    .Y(_07660_));
 sky130_fd_sc_hd__nand2_1 _12146_ (.A(message[21]),
    .B(_07568_),
    .Y(_07663_));
 sky130_fd_sc_hd__o21ai_0 _12147_ (.A1(_07568_),
    .A2(_07660_),
    .B1(_07663_),
    .Y(_00130_));
 sky130_fd_sc_hd__a31o_2 _12149_ (.A1(_09402_),
    .A2(_07640_),
    .A3(_07642_),
    .B1(_09401_),
    .X(_07665_));
 sky130_fd_sc_hd__a21oi_1 _12150_ (.A1(_09406_),
    .A2(_07665_),
    .B1(_09405_),
    .Y(_07666_));
 sky130_fd_sc_hd__xor2_1 _12151_ (.A(_09410_),
    .B(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__nor2_1 _12152_ (.A(done),
    .B(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__a21oi_1 _12153_ (.A1(\w[62][11] ),
    .A2(done),
    .B1(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__nand2_1 _12155_ (.A(message[20]),
    .B(_07568_),
    .Y(_07671_));
 sky130_fd_sc_hd__o21ai_0 _12156_ (.A1(_07568_),
    .A2(_07669_),
    .B1(_07671_),
    .Y(_00131_));
 sky130_fd_sc_hd__o21a_1 _12158_ (.A1(_09405_),
    .A2(_07655_),
    .B1(_09410_),
    .X(_07673_));
 sky130_fd_sc_hd__nor2_1 _12159_ (.A(_09409_),
    .B(_07673_),
    .Y(_07674_));
 sky130_fd_sc_hd__xnor2_1 _12160_ (.A(_09414_),
    .B(_07674_),
    .Y(_07675_));
 sky130_fd_sc_hd__mux2i_2 _12162_ (.A0(\w[62][12] ),
    .A1(_07675_),
    .S(_07591_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand2_1 _12164_ (.A(message[19]),
    .B(_07568_),
    .Y(_07679_));
 sky130_fd_sc_hd__o21ai_0 _12165_ (.A1(_07568_),
    .A2(_07677_),
    .B1(_07679_),
    .Y(_00132_));
 sky130_fd_sc_hd__inv_1 _12166_ (.A(_09418_),
    .Y(_07680_));
 sky130_fd_sc_hd__and3_1 _12167_ (.A(_09406_),
    .B(_09410_),
    .C(_09414_),
    .X(_07681_));
 sky130_fd_sc_hd__and2_1 _12168_ (.A(_09402_),
    .B(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__a21o_1 _12169_ (.A1(_09406_),
    .A2(_09401_),
    .B1(_09405_),
    .X(_07683_));
 sky130_fd_sc_hd__a21o_1 _12170_ (.A1(_09410_),
    .A2(_07683_),
    .B1(_09409_),
    .X(_07684_));
 sky130_fd_sc_hd__a21o_1 _12171_ (.A1(_09414_),
    .A2(_07684_),
    .B1(_09413_),
    .X(_07685_));
 sky130_fd_sc_hd__a31oi_1 _12172_ (.A1(_07640_),
    .A2(_07642_),
    .A3(_07682_),
    .B1(_07685_),
    .Y(_07686_));
 sky130_fd_sc_hd__xnor2_1 _12173_ (.A(_07680_),
    .B(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__nand2_1 _12174_ (.A(_07591_),
    .B(_07687_),
    .Y(_07688_));
 sky130_fd_sc_hd__o21ai_1 _12175_ (.A1(\w[62][13] ),
    .A2(_07591_),
    .B1(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__nand2_1 _12177_ (.A(message[18]),
    .B(_07568_),
    .Y(_07691_));
 sky130_fd_sc_hd__o21ai_0 _12178_ (.A1(_07568_),
    .A2(_07689_),
    .B1(_07691_),
    .Y(_00133_));
 sky130_fd_sc_hd__o21ai_0 _12179_ (.A1(_07649_),
    .A2(_07650_),
    .B1(_07651_),
    .Y(_07692_));
 sky130_fd_sc_hd__and2_1 _12180_ (.A(_09418_),
    .B(_07681_),
    .X(_07693_));
 sky130_fd_sc_hd__a21oi_1 _12181_ (.A1(_09410_),
    .A2(_09405_),
    .B1(_09409_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand2_1 _12182_ (.A(_09414_),
    .B(_09418_),
    .Y(_07695_));
 sky130_fd_sc_hd__a21oi_1 _12183_ (.A1(_09418_),
    .A2(_09413_),
    .B1(_09417_),
    .Y(_07696_));
 sky130_fd_sc_hd__o21ai_0 _12184_ (.A1(_07694_),
    .A2(_07695_),
    .B1(_07696_),
    .Y(_07697_));
 sky130_fd_sc_hd__a21oi_1 _12185_ (.A1(_07692_),
    .A2(_07693_),
    .B1(_07697_),
    .Y(_07698_));
 sky130_fd_sc_hd__nand4_1 _12186_ (.A(_07614_),
    .B(_07615_),
    .C(_07653_),
    .D(_07693_),
    .Y(_07699_));
 sky130_fd_sc_hd__nand2_1 _12187_ (.A(_07698_),
    .B(_07699_),
    .Y(_07700_));
 sky130_fd_sc_hd__xnor2_1 _12188_ (.A(_09422_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__nor2_1 _12189_ (.A(done),
    .B(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__a21oi_1 _12190_ (.A1(\w[62][14] ),
    .A2(done),
    .B1(_07702_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand2_1 _12192_ (.A(message[17]),
    .B(_07568_),
    .Y(_07705_));
 sky130_fd_sc_hd__o21ai_0 _12193_ (.A1(_07568_),
    .A2(_07703_),
    .B1(_07705_),
    .Y(_00134_));
 sky130_fd_sc_hd__o21bai_1 _12194_ (.A1(_07680_),
    .A2(_07686_),
    .B1_N(_09417_),
    .Y(_07706_));
 sky130_fd_sc_hd__a21oi_1 _12195_ (.A1(_09422_),
    .A2(_07706_),
    .B1(_09421_),
    .Y(_07707_));
 sky130_fd_sc_hd__xnor2_1 _12196_ (.A(_09430_),
    .B(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__mux2i_2 _12197_ (.A0(\w[62][15] ),
    .A1(_07708_),
    .S(_07591_),
    .Y(_07709_));
 sky130_fd_sc_hd__nand2_1 _12199_ (.A(message[16]),
    .B(_07568_),
    .Y(_07711_));
 sky130_fd_sc_hd__o21ai_0 _12200_ (.A1(_07568_),
    .A2(_07709_),
    .B1(_07711_),
    .Y(_00135_));
 sky130_fd_sc_hd__a21o_1 _12201_ (.A1(_09422_),
    .A2(_07700_),
    .B1(_09421_),
    .X(_07712_));
 sky130_fd_sc_hd__a21oi_1 _12202_ (.A1(_09430_),
    .A2(_07712_),
    .B1(_09429_),
    .Y(_07713_));
 sky130_fd_sc_hd__xnor2_1 _12203_ (.A(_09426_),
    .B(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__mux2i_2 _12204_ (.A0(\w[62][16] ),
    .A1(_07714_),
    .S(_07591_),
    .Y(_07715_));
 sky130_fd_sc_hd__nand2_1 _12206_ (.A(message[15]),
    .B(_07568_),
    .Y(_07717_));
 sky130_fd_sc_hd__o21ai_0 _12207_ (.A1(_07568_),
    .A2(_07715_),
    .B1(_07717_),
    .Y(_00136_));
 sky130_fd_sc_hd__inv_1 _12208_ (.A(_09421_),
    .Y(_07718_));
 sky130_fd_sc_hd__o21ai_0 _12209_ (.A1(_09418_),
    .A2(_09417_),
    .B1(_09422_),
    .Y(_07719_));
 sky130_fd_sc_hd__nand2_1 _12210_ (.A(_09430_),
    .B(_09426_),
    .Y(_07720_));
 sky130_fd_sc_hd__a21oi_1 _12211_ (.A1(_07718_),
    .A2(_07719_),
    .B1(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__nand2_1 _12212_ (.A(_09422_),
    .B(_09417_),
    .Y(_07722_));
 sky130_fd_sc_hd__nand2_1 _12213_ (.A(_07718_),
    .B(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__a311o_1 _12214_ (.A1(_07640_),
    .A2(_07642_),
    .A3(_07682_),
    .B1(_07685_),
    .C1(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__a21o_1 _12215_ (.A1(_09426_),
    .A2(_09429_),
    .B1(_09425_),
    .X(_07725_));
 sky130_fd_sc_hd__a211oi_1 _12216_ (.A1(_07721_),
    .A2(_07724_),
    .B1(_09434_),
    .C1(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__nor2_1 _12217_ (.A(_07725_),
    .B(_07723_),
    .Y(_07727_));
 sky130_fd_sc_hd__o21ai_0 _12218_ (.A1(_07725_),
    .A2(_07721_),
    .B1(_09434_),
    .Y(_07728_));
 sky130_fd_sc_hd__a21oi_1 _12219_ (.A1(_07686_),
    .A2(_07727_),
    .B1(_07728_),
    .Y(_07729_));
 sky130_fd_sc_hd__nor3_1 _12220_ (.A(done),
    .B(_07726_),
    .C(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__a21oi_1 _12221_ (.A1(\w[62][17] ),
    .A2(done),
    .B1(_07730_),
    .Y(_07731_));
 sky130_fd_sc_hd__nand2_1 _12223_ (.A(message[14]),
    .B(_07568_),
    .Y(_07733_));
 sky130_fd_sc_hd__o21ai_0 _12224_ (.A1(_07568_),
    .A2(_07731_),
    .B1(_07733_),
    .Y(_00137_));
 sky130_fd_sc_hd__o21ai_0 _12225_ (.A1(_09422_),
    .A2(_09421_),
    .B1(_09430_),
    .Y(_07734_));
 sky130_fd_sc_hd__nor2_1 _12226_ (.A(_09425_),
    .B(_09429_),
    .Y(_07735_));
 sky130_fd_sc_hd__nor2_1 _12227_ (.A(_09426_),
    .B(_09425_),
    .Y(_07736_));
 sky130_fd_sc_hd__a21oi_1 _12228_ (.A1(_07734_),
    .A2(_07735_),
    .B1(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__a21oi_1 _12229_ (.A1(_09434_),
    .A2(_07737_),
    .B1(_09433_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand2_1 _12230_ (.A(_09434_),
    .B(_09425_),
    .Y(_07739_));
 sky130_fd_sc_hd__a211oi_1 _12231_ (.A1(_09430_),
    .A2(_09421_),
    .B1(_09429_),
    .C1(_09433_),
    .Y(_07740_));
 sky130_fd_sc_hd__nand2_1 _12232_ (.A(_07739_),
    .B(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__nor2_1 _12233_ (.A(_07700_),
    .B(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__nor2_1 _12234_ (.A(_07738_),
    .B(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__xor2_1 _12235_ (.A(_09438_),
    .B(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__mux2i_2 _12236_ (.A0(\w[62][18] ),
    .A1(_07744_),
    .S(_07591_),
    .Y(_07745_));
 sky130_fd_sc_hd__nand2_1 _12238_ (.A(message[13]),
    .B(_07568_),
    .Y(_07747_));
 sky130_fd_sc_hd__o21ai_0 _12239_ (.A1(_07568_),
    .A2(_07745_),
    .B1(_07747_),
    .Y(_00138_));
 sky130_fd_sc_hd__inv_1 _12240_ (.A(_09437_),
    .Y(_07748_));
 sky130_fd_sc_hd__o21ai_0 _12241_ (.A1(_09433_),
    .A2(_07729_),
    .B1(_09438_),
    .Y(_07749_));
 sky130_fd_sc_hd__a211oi_1 _12242_ (.A1(_07748_),
    .A2(_07749_),
    .B1(done),
    .C1(_09442_),
    .Y(_07750_));
 sky130_fd_sc_hd__and4_1 _12243_ (.A(_09442_),
    .B(_07748_),
    .C(_07591_),
    .D(_07749_),
    .X(_07751_));
 sky130_fd_sc_hd__a211oi_2 _12244_ (.A1(\w[62][19] ),
    .A2(done),
    .B1(_07750_),
    .C1(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__nand2_1 _12246_ (.A(message[12]),
    .B(_07568_),
    .Y(_07754_));
 sky130_fd_sc_hd__o21ai_0 _12247_ (.A1(_07568_),
    .A2(_07752_),
    .B1(_07754_),
    .Y(_00139_));
 sky130_fd_sc_hd__a21oi_1 _12249_ (.A1(_09442_),
    .A2(_09437_),
    .B1(_09441_),
    .Y(_07756_));
 sky130_fd_sc_hd__nand3_1 _12250_ (.A(_07739_),
    .B(_07740_),
    .C(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__a211oi_1 _12251_ (.A1(_07692_),
    .A2(_07693_),
    .B1(_07757_),
    .C1(_07697_),
    .Y(_07758_));
 sky130_fd_sc_hd__and3_1 _12252_ (.A(_09434_),
    .B(_09438_),
    .C(_09442_),
    .X(_07759_));
 sky130_fd_sc_hd__nand3_1 _12253_ (.A(_09438_),
    .B(_09442_),
    .C(_09433_),
    .Y(_07760_));
 sky130_fd_sc_hd__nand2_1 _12254_ (.A(_07756_),
    .B(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__a21oi_1 _12255_ (.A1(_07737_),
    .A2(_07759_),
    .B1(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__a21oi_1 _12256_ (.A1(_07699_),
    .A2(_07758_),
    .B1(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__xnor2_1 _12257_ (.A(_09446_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__nand2_1 _12258_ (.A(_07591_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__o21ai_1 _12259_ (.A1(\w[62][20] ),
    .A2(_07591_),
    .B1(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__nand2_1 _12261_ (.A(message[11]),
    .B(_07568_),
    .Y(_07768_));
 sky130_fd_sc_hd__o21ai_0 _12262_ (.A1(_07568_),
    .A2(_07766_),
    .B1(_07768_),
    .Y(_00141_));
 sky130_fd_sc_hd__nand4_1 _12263_ (.A(_09434_),
    .B(_09438_),
    .C(_09442_),
    .D(_09446_),
    .Y(_07769_));
 sky130_fd_sc_hd__a211oi_1 _12264_ (.A1(_07718_),
    .A2(_07719_),
    .B1(_07769_),
    .C1(_07720_),
    .Y(_07770_));
 sky130_fd_sc_hd__a21o_1 _12265_ (.A1(_09434_),
    .A2(_07725_),
    .B1(_09433_),
    .X(_07771_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(_09438_),
    .A2(_07771_),
    .B1(_09437_),
    .X(_07772_));
 sky130_fd_sc_hd__a21o_1 _12267_ (.A1(_09442_),
    .A2(_07772_),
    .B1(_09441_),
    .X(_07773_));
 sky130_fd_sc_hd__a221oi_1 _12268_ (.A1(_07724_),
    .A2(_07770_),
    .B1(_07773_),
    .B2(_09446_),
    .C1(_09445_),
    .Y(_07774_));
 sky130_fd_sc_hd__xor2_1 _12269_ (.A(_09450_),
    .B(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__nor2_1 _12270_ (.A(done),
    .B(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__a21oi_1 _12271_ (.A1(\w[62][21] ),
    .A2(done),
    .B1(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__nand2_1 _12273_ (.A(message[10]),
    .B(_07568_),
    .Y(_07779_));
 sky130_fd_sc_hd__o21ai_0 _12274_ (.A1(_07568_),
    .A2(_07777_),
    .B1(_07779_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _12275_ (.A(_09446_),
    .B(_09450_),
    .Y(_07780_));
 sky130_fd_sc_hd__a211oi_1 _12276_ (.A1(_07699_),
    .A2(_07758_),
    .B1(_07762_),
    .C1(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__a21o_1 _12277_ (.A1(_09450_),
    .A2(_09445_),
    .B1(_09449_),
    .X(_07782_));
 sky130_fd_sc_hd__o21a_1 _12278_ (.A1(_07781_),
    .A2(_07782_),
    .B1(_09454_),
    .X(_07783_));
 sky130_fd_sc_hd__nor3_1 _12279_ (.A(_09454_),
    .B(_07781_),
    .C(_07782_),
    .Y(_07784_));
 sky130_fd_sc_hd__o21ai_0 _12280_ (.A1(_07783_),
    .A2(_07784_),
    .B1(_07591_),
    .Y(_07785_));
 sky130_fd_sc_hd__o21ai_1 _12281_ (.A1(\w[62][22] ),
    .A2(_07591_),
    .B1(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__nand2_1 _12283_ (.A(message[9]),
    .B(_07568_),
    .Y(_07788_));
 sky130_fd_sc_hd__o21ai_0 _12284_ (.A1(_07568_),
    .A2(_07786_),
    .B1(_07788_),
    .Y(_00143_));
 sky130_fd_sc_hd__nand2_1 _12285_ (.A(_09450_),
    .B(_09454_),
    .Y(_07789_));
 sky130_fd_sc_hd__a21oi_1 _12286_ (.A1(_09446_),
    .A2(_09441_),
    .B1(_09445_),
    .Y(_07790_));
 sky130_fd_sc_hd__a21o_1 _12287_ (.A1(_09454_),
    .A2(_09449_),
    .B1(_09453_),
    .X(_07791_));
 sky130_fd_sc_hd__nor3_1 _12288_ (.A(_09433_),
    .B(_09437_),
    .C(_07791_),
    .Y(_07792_));
 sky130_fd_sc_hd__o21ai_0 _12289_ (.A1(_07789_),
    .A2(_07790_),
    .B1(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__o21ai_0 _12290_ (.A1(_09438_),
    .A2(_09437_),
    .B1(_09442_),
    .Y(_07794_));
 sky130_fd_sc_hd__nand2b_1 _12291_ (.A_N(_09441_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__a21oi_1 _12292_ (.A1(_09446_),
    .A2(_07795_),
    .B1(_09445_),
    .Y(_07796_));
 sky130_fd_sc_hd__o21bai_1 _12293_ (.A1(_07789_),
    .A2(_07796_),
    .B1_N(_07791_),
    .Y(_07797_));
 sky130_fd_sc_hd__o21ai_0 _12294_ (.A1(_07729_),
    .A2(_07793_),
    .B1(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__xnor2_1 _12295_ (.A(_09458_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__mux2i_2 _12296_ (.A0(\w[62][23] ),
    .A1(_07799_),
    .S(_07591_),
    .Y(_07800_));
 sky130_fd_sc_hd__nand2_1 _12298_ (.A(message[8]),
    .B(_07568_),
    .Y(_07802_));
 sky130_fd_sc_hd__o21ai_0 _12299_ (.A1(_07568_),
    .A2(_07800_),
    .B1(_07802_),
    .Y(_00144_));
 sky130_fd_sc_hd__and2_1 _12300_ (.A(_05338_),
    .B(_07566_),
    .X(_07803_));
 sky130_fd_sc_hd__o21a_1 _12302_ (.A1(_09453_),
    .A2(_07783_),
    .B1(_09458_),
    .X(_07805_));
 sky130_fd_sc_hd__nor3_1 _12303_ (.A(_09462_),
    .B(_09457_),
    .C(_07805_),
    .Y(_07806_));
 sky130_fd_sc_hd__o21a_1 _12304_ (.A1(_09457_),
    .A2(_07805_),
    .B1(_09462_),
    .X(_07807_));
 sky130_fd_sc_hd__nand2_1 _12305_ (.A(\w[62][24] ),
    .B(done),
    .Y(_07808_));
 sky130_fd_sc_hd__o31a_1 _12306_ (.A1(done),
    .A2(_07806_),
    .A3(_07807_),
    .B1(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__nor2_1 _12307_ (.A(message[7]),
    .B(_07803_),
    .Y(_07810_));
 sky130_fd_sc_hd__a21oi_1 _12308_ (.A1(_07803_),
    .A2(_07809_),
    .B1(_07810_),
    .Y(_00145_));
 sky130_fd_sc_hd__nand4_1 _12309_ (.A(_09450_),
    .B(_09454_),
    .C(_09458_),
    .D(_09462_),
    .Y(_07811_));
 sky130_fd_sc_hd__a21o_1 _12310_ (.A1(_09458_),
    .A2(_07791_),
    .B1(_09457_),
    .X(_07812_));
 sky130_fd_sc_hd__a21oi_1 _12311_ (.A1(_09462_),
    .A2(_07812_),
    .B1(_09461_),
    .Y(_07813_));
 sky130_fd_sc_hd__o21ai_0 _12312_ (.A1(_07774_),
    .A2(_07811_),
    .B1(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__or2_2 _12313_ (.A(_09466_),
    .B(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__nand2_1 _12314_ (.A(_09466_),
    .B(_07814_),
    .Y(_07816_));
 sky130_fd_sc_hd__and2_1 _12315_ (.A(\w[62][25] ),
    .B(done),
    .X(_07817_));
 sky130_fd_sc_hd__a31oi_2 _12316_ (.A1(_07591_),
    .A2(_07815_),
    .A3(_07816_),
    .B1(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__nand2_1 _12318_ (.A(message[6]),
    .B(_07568_),
    .Y(_07820_));
 sky130_fd_sc_hd__o21ai_0 _12319_ (.A1(_07568_),
    .A2(_07818_),
    .B1(_07820_),
    .Y(_00146_));
 sky130_fd_sc_hd__and3_1 _12320_ (.A(_09458_),
    .B(_09462_),
    .C(_09466_),
    .X(_07821_));
 sky130_fd_sc_hd__nand3_1 _12321_ (.A(_09454_),
    .B(_07782_),
    .C(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__nand4_1 _12322_ (.A(_09446_),
    .B(_09450_),
    .C(_09454_),
    .D(_07821_),
    .Y(_07823_));
 sky130_fd_sc_hd__a211o_1 _12323_ (.A1(_07699_),
    .A2(_07758_),
    .B1(_07762_),
    .C1(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__a21o_1 _12324_ (.A1(_09458_),
    .A2(_09453_),
    .B1(_09457_),
    .X(_07825_));
 sky130_fd_sc_hd__a21o_1 _12325_ (.A1(_09462_),
    .A2(_07825_),
    .B1(_09461_),
    .X(_07826_));
 sky130_fd_sc_hd__a21oi_1 _12326_ (.A1(_09466_),
    .A2(_07826_),
    .B1(_09465_),
    .Y(_07827_));
 sky130_fd_sc_hd__and3_1 _12327_ (.A(_07822_),
    .B(_07824_),
    .C(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__xor2_1 _12328_ (.A(_09470_),
    .B(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__nand2_1 _12329_ (.A(_07591_),
    .B(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__o21ai_1 _12330_ (.A1(\w[62][26] ),
    .A2(_07591_),
    .B1(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__nand2_1 _12332_ (.A(message[5]),
    .B(_07568_),
    .Y(_07833_));
 sky130_fd_sc_hd__o21ai_0 _12333_ (.A1(_07568_),
    .A2(_07831_),
    .B1(_07833_),
    .Y(_00147_));
 sky130_fd_sc_hd__and3_1 _12334_ (.A(_09470_),
    .B(_07797_),
    .C(_07821_),
    .X(_07834_));
 sky130_fd_sc_hd__o21ai_0 _12335_ (.A1(_07729_),
    .A2(_07793_),
    .B1(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__a21o_1 _12336_ (.A1(_09462_),
    .A2(_09457_),
    .B1(_09461_),
    .X(_07836_));
 sky130_fd_sc_hd__a21o_1 _12337_ (.A1(_09466_),
    .A2(_07836_),
    .B1(_09465_),
    .X(_07837_));
 sky130_fd_sc_hd__a21oi_1 _12338_ (.A1(_09470_),
    .A2(_07837_),
    .B1(_09469_),
    .Y(_07838_));
 sky130_fd_sc_hd__a21boi_0 _12339_ (.A1(_07835_),
    .A2(_07838_),
    .B1_N(_09474_),
    .Y(_07839_));
 sky130_fd_sc_hd__a21o_1 _12340_ (.A1(_09470_),
    .A2(_07837_),
    .B1(_09469_),
    .X(_07840_));
 sky130_fd_sc_hd__nor3b_1 _12341_ (.A(_09474_),
    .B(_07840_),
    .C_N(_07835_),
    .Y(_07841_));
 sky130_fd_sc_hd__nand2_1 _12342_ (.A(\w[62][27] ),
    .B(done),
    .Y(_07842_));
 sky130_fd_sc_hd__o31a_1 _12343_ (.A1(done),
    .A2(_07839_),
    .A3(_07841_),
    .B1(_07842_),
    .X(_07843_));
 sky130_fd_sc_hd__nand2_1 _12345_ (.A(message[4]),
    .B(_07568_),
    .Y(_07845_));
 sky130_fd_sc_hd__o21ai_0 _12346_ (.A1(_07568_),
    .A2(_07843_),
    .B1(_07845_),
    .Y(_00148_));
 sky130_fd_sc_hd__nand2_1 _12347_ (.A(_09470_),
    .B(_09474_),
    .Y(_07846_));
 sky130_fd_sc_hd__a21oi_1 _12348_ (.A1(_09474_),
    .A2(_09469_),
    .B1(_09473_),
    .Y(_07847_));
 sky130_fd_sc_hd__o21ai_0 _12349_ (.A1(_07828_),
    .A2(_07846_),
    .B1(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__xor2_1 _12350_ (.A(_09478_),
    .B(_07848_),
    .X(_07849_));
 sky130_fd_sc_hd__mux2i_2 _12351_ (.A0(\w[62][28] ),
    .A1(_07849_),
    .S(_07591_),
    .Y(_07850_));
 sky130_fd_sc_hd__nor2_1 _12352_ (.A(message[3]),
    .B(_07803_),
    .Y(_07851_));
 sky130_fd_sc_hd__a21oi_1 _12353_ (.A1(_07803_),
    .A2(_07850_),
    .B1(_07851_),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_1 _12354_ (.A(_09482_),
    .Y(_07852_));
 sky130_fd_sc_hd__a21oi_1 _12355_ (.A1(_09478_),
    .A2(_09473_),
    .B1(_09477_),
    .Y(_07853_));
 sky130_fd_sc_hd__nand3_1 _12356_ (.A(_07852_),
    .B(_07591_),
    .C(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__nand2_1 _12357_ (.A(_09482_),
    .B(_07591_),
    .Y(_07855_));
 sky130_fd_sc_hd__nand3_1 _12358_ (.A(_09474_),
    .B(_09478_),
    .C(_07840_),
    .Y(_07856_));
 sky130_fd_sc_hd__o2111ai_1 _12359_ (.A1(_07729_),
    .A2(_07793_),
    .B1(_07834_),
    .C1(_09478_),
    .D1(_09474_),
    .Y(_07857_));
 sky130_fd_sc_hd__nand2_1 _12360_ (.A(_07856_),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__mux2i_1 _12361_ (.A0(_07854_),
    .A1(_07855_),
    .S(_07858_),
    .Y(_07859_));
 sky130_fd_sc_hd__o22ai_1 _12362_ (.A1(\w[62][29] ),
    .A2(_07591_),
    .B1(_07853_),
    .B2(_07855_),
    .Y(_07860_));
 sky130_fd_sc_hd__nor2_1 _12363_ (.A(_07568_),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__a21oi_1 _12364_ (.A1(message[2]),
    .A2(_07568_),
    .B1(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__a21oi_1 _12365_ (.A1(_07803_),
    .A2(_07859_),
    .B1(_07862_),
    .Y(_00150_));
 sky130_fd_sc_hd__inv_1 _12366_ (.A(_09486_),
    .Y(_07863_));
 sky130_fd_sc_hd__inv_1 _12367_ (.A(_09477_),
    .Y(_07864_));
 sky130_fd_sc_hd__nand2_1 _12368_ (.A(_07847_),
    .B(_07846_),
    .Y(_07865_));
 sky130_fd_sc_hd__a21oi_1 _12369_ (.A1(_09478_),
    .A2(_07865_),
    .B1(_09477_),
    .Y(_07866_));
 sky130_fd_sc_hd__a31oi_1 _12370_ (.A1(_07864_),
    .A2(_07828_),
    .A3(_07847_),
    .B1(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__nor2_1 _12371_ (.A(_09486_),
    .B(_07855_),
    .Y(_07868_));
 sky130_fd_sc_hd__nor3_1 _12372_ (.A(_09482_),
    .B(_07863_),
    .C(_09481_),
    .Y(_07869_));
 sky130_fd_sc_hd__a21oi_1 _12373_ (.A1(_07863_),
    .A2(_09481_),
    .B1(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__nor2_1 _12374_ (.A(done),
    .B(_07870_),
    .Y(_07871_));
 sky130_fd_sc_hd__a221oi_1 _12375_ (.A1(\w[62][30] ),
    .A2(done),
    .B1(_07867_),
    .B2(_07868_),
    .C1(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__o41a_1 _12376_ (.A1(_07863_),
    .A2(_09481_),
    .A3(done),
    .A4(_07867_),
    .B1(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__nand2_1 _12378_ (.A(message[1]),
    .B(_07568_),
    .Y(_07875_));
 sky130_fd_sc_hd__o21ai_0 _12379_ (.A1(_07568_),
    .A2(_07873_),
    .B1(_07875_),
    .Y(_00152_));
 sky130_fd_sc_hd__nand2_1 _12380_ (.A(_09474_),
    .B(_09478_),
    .Y(_07876_));
 sky130_fd_sc_hd__nor3_1 _12381_ (.A(_07852_),
    .B(_07863_),
    .C(_07876_),
    .Y(_07877_));
 sky130_fd_sc_hd__o211ai_1 _12382_ (.A1(_07729_),
    .A2(_07793_),
    .B1(_07834_),
    .C1(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__o21bai_1 _12383_ (.A1(_07852_),
    .A2(_07853_),
    .B1_N(_09481_),
    .Y(_07879_));
 sky130_fd_sc_hd__a221oi_1 _12384_ (.A1(_09486_),
    .A2(_07879_),
    .B1(_07877_),
    .B2(_07840_),
    .C1(_09485_),
    .Y(_07880_));
 sky130_fd_sc_hd__mux4_2 _12385_ (.A0(\w[4][31] ),
    .A1(\w[12][31] ),
    .A2(\w[6][31] ),
    .A3(\w[14][31] ),
    .S0(\count16_1[3] ),
    .S1(\count16_1[1] ),
    .X(_07881_));
 sky130_fd_sc_hd__mux4_2 _12386_ (.A0(\w[36][31] ),
    .A1(\w[44][31] ),
    .A2(\w[38][31] ),
    .A3(\w[46][31] ),
    .S0(\count16_1[3] ),
    .S1(\count16_1[1] ),
    .X(_07882_));
 sky130_fd_sc_hd__mux2i_1 _12387_ (.A0(_07881_),
    .A1(_07882_),
    .S(\count16_1[5] ),
    .Y(_07883_));
 sky130_fd_sc_hd__nor3b_1 _12388_ (.A(\count16_1[4] ),
    .B(_07883_),
    .C_N(\count16_1[2] ),
    .Y(_07884_));
 sky130_fd_sc_hd__mux4_2 _12389_ (.A0(\w[0][31] ),
    .A1(\w[8][31] ),
    .A2(\w[32][31] ),
    .A3(\w[40][31] ),
    .S0(\count16_1[3] ),
    .S1(\count16_1[5] ),
    .X(_07885_));
 sky130_fd_sc_hd__mux4_2 _12390_ (.A0(\w[2][31] ),
    .A1(\w[10][31] ),
    .A2(\w[34][31] ),
    .A3(\w[42][31] ),
    .S0(\count16_1[3] ),
    .S1(\count16_1[5] ),
    .X(_07886_));
 sky130_fd_sc_hd__mux2i_1 _12391_ (.A0(_07885_),
    .A1(_07886_),
    .S(\count16_1[1] ),
    .Y(_07887_));
 sky130_fd_sc_hd__nor3_1 _12392_ (.A(\count16_1[2] ),
    .B(\count16_1[4] ),
    .C(_07887_),
    .Y(_07888_));
 sky130_fd_sc_hd__mux4_2 _12393_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07889_));
 sky130_fd_sc_hd__mux4_2 _12394_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07890_));
 sky130_fd_sc_hd__mux2i_1 _12395_ (.A0(_07889_),
    .A1(_07890_),
    .S(\count16_1[5] ),
    .Y(_07891_));
 sky130_fd_sc_hd__nand2_1 _12396_ (.A(\count16_1[3] ),
    .B(\count16_1[4] ),
    .Y(_07892_));
 sky130_fd_sc_hd__nand2b_1 _12397_ (.A_N(\count16_1[3] ),
    .B(\count16_1[4] ),
    .Y(_07893_));
 sky130_fd_sc_hd__mux4_2 _12398_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[48][31] ),
    .A3(\w[52][31] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[5] ),
    .X(_07894_));
 sky130_fd_sc_hd__mux4_2 _12399_ (.A0(\w[18][31] ),
    .A1(\w[22][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[5] ),
    .X(_07895_));
 sky130_fd_sc_hd__mux2i_1 _12400_ (.A0(_07894_),
    .A1(_07895_),
    .S(\count16_1[1] ),
    .Y(_07896_));
 sky130_fd_sc_hd__o22ai_1 _12401_ (.A1(_07891_),
    .A2(_07892_),
    .B1(_07893_),
    .B2(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__nor3_1 _12402_ (.A(_07884_),
    .B(_07888_),
    .C(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__xnor2_1 _12403_ (.A(_09068_),
    .B(_09063_),
    .Y(_07899_));
 sky130_fd_sc_hd__xnor2_1 _12404_ (.A(\w_new_calc1.temp2[31] ),
    .B(\w_new_calc1.temp1[31] ),
    .Y(_07900_));
 sky130_fd_sc_hd__xnor2_1 _12405_ (.A(_07899_),
    .B(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__xnor2_1 _12406_ (.A(_07898_),
    .B(_07901_),
    .Y(_07902_));
 sky130_fd_sc_hd__mux4_2 _12407_ (.A0(\w[9][31] ),
    .A1(\w[11][31] ),
    .A2(\w[13][31] ),
    .A3(\w[15][31] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07903_));
 sky130_fd_sc_hd__mux4_2 _12408_ (.A0(\w[25][31] ),
    .A1(\w[27][31] ),
    .A2(\w[29][31] ),
    .A3(\w[31][31] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07904_));
 sky130_fd_sc_hd__mux4_2 _12409_ (.A0(\w[41][31] ),
    .A1(\w[43][31] ),
    .A2(\w[45][31] ),
    .A3(\w[47][31] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07905_));
 sky130_fd_sc_hd__mux4_2 _12410_ (.A0(\w[57][31] ),
    .A1(\w[59][31] ),
    .A2(\w[61][31] ),
    .A3(\w[63][31] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_07906_));
 sky130_fd_sc_hd__mux4_2 _12411_ (.A0(_07903_),
    .A1(_07904_),
    .A2(_07905_),
    .A3(_07906_),
    .S0(\count7_1[4] ),
    .S1(\count7_1[5] ),
    .X(_07907_));
 sky130_fd_sc_hd__inv_1 _12412_ (.A(\count7_1[1] ),
    .Y(_07908_));
 sky130_fd_sc_hd__mux4_2 _12413_ (.A0(\w[3][31] ),
    .A1(\w[7][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[4] ),
    .X(_07909_));
 sky130_fd_sc_hd__nor2_1 _12414_ (.A(\count7_1[3] ),
    .B(\count7_1[5] ),
    .Y(_07910_));
 sky130_fd_sc_hd__o21ai_0 _12415_ (.A1(_07908_),
    .A2(_07909_),
    .B1(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__mux4_2 _12416_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[17][31] ),
    .A3(\w[21][31] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[4] ),
    .X(_07912_));
 sky130_fd_sc_hd__nor2b_1 _12417_ (.A(_07911_),
    .B_N(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__nor2b_1 _12418_ (.A(\count7_1[3] ),
    .B_N(\count7_1[5] ),
    .Y(_07914_));
 sky130_fd_sc_hd__mux4_2 _12419_ (.A0(\w[35][31] ),
    .A1(\w[39][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[4] ),
    .X(_07915_));
 sky130_fd_sc_hd__nand2_1 _12420_ (.A(_07914_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__mux4_2 _12421_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[49][31] ),
    .A3(\w[53][31] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[4] ),
    .X(_07917_));
 sky130_fd_sc_hd__a21oi_1 _12422_ (.A1(_07914_),
    .A2(_07917_),
    .B1(\count7_1[1] ),
    .Y(_07918_));
 sky130_fd_sc_hd__a31oi_1 _12423_ (.A1(\count7_1[1] ),
    .A2(_07911_),
    .A3(_07916_),
    .B1(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__a211o_1 _12424_ (.A1(\count7_1[3] ),
    .A2(_07907_),
    .B1(_07913_),
    .C1(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__xnor2_1 _12425_ (.A(_07902_),
    .B(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__a21oi_1 _12426_ (.A1(_07878_),
    .A2(_07880_),
    .B1(_07921_),
    .Y(_07922_));
 sky130_fd_sc_hd__and3_1 _12427_ (.A(_07921_),
    .B(_07878_),
    .C(_07880_),
    .X(_07923_));
 sky130_fd_sc_hd__nand2_1 _12428_ (.A(\w[62][31] ),
    .B(done),
    .Y(_07924_));
 sky130_fd_sc_hd__o31a_1 _12429_ (.A1(done),
    .A2(_07922_),
    .A3(_07923_),
    .B1(_07924_),
    .X(_07925_));
 sky130_fd_sc_hd__nor2_1 _12430_ (.A(message[0]),
    .B(_07803_),
    .Y(_07926_));
 sky130_fd_sc_hd__a21oi_1 _12431_ (.A1(_07803_),
    .A2(_07925_),
    .B1(_07926_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2b_1 _12432_ (.A(reset),
    .B_N(_09562_),
    .Y(_07927_));
 sky130_fd_sc_hd__nand2_1 _12433_ (.A(_05403_),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__mux2i_2 _12435_ (.A0(_09489_),
    .A1(\w[63][0] ),
    .S(done),
    .Y(_07930_));
 sky130_fd_sc_hd__nand2_1 _12438_ (.A(message[63]),
    .B(_07928_),
    .Y(_07933_));
 sky130_fd_sc_hd__o21ai_0 _12439_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_07933_),
    .Y(_00353_));
 sky130_fd_sc_hd__mux2i_2 _12440_ (.A0(_09490_),
    .A1(\w[63][1] ),
    .S(done),
    .Y(_07934_));
 sky130_fd_sc_hd__nand2_1 _12442_ (.A(message[62]),
    .B(_07928_),
    .Y(_07936_));
 sky130_fd_sc_hd__o21ai_0 _12443_ (.A1(_07928_),
    .A2(_07934_),
    .B1(_07936_),
    .Y(_00364_));
 sky130_fd_sc_hd__mux2i_2 _12444_ (.A0(_09095_),
    .A1(\w[63][2] ),
    .S(done),
    .Y(_07937_));
 sky130_fd_sc_hd__nand2_1 _12446_ (.A(message[61]),
    .B(_07928_),
    .Y(_07939_));
 sky130_fd_sc_hd__o21ai_0 _12447_ (.A1(_07928_),
    .A2(_07937_),
    .B1(_07939_),
    .Y(_00375_));
 sky130_fd_sc_hd__xnor2_1 _12448_ (.A(_09094_),
    .B(_09494_),
    .Y(_07940_));
 sky130_fd_sc_hd__nor2_1 _12449_ (.A(done),
    .B(_07940_),
    .Y(_07941_));
 sky130_fd_sc_hd__a21oi_1 _12450_ (.A1(\w[63][3] ),
    .A2(done),
    .B1(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__nand2_1 _12452_ (.A(message[60]),
    .B(_07928_),
    .Y(_07944_));
 sky130_fd_sc_hd__o21ai_0 _12453_ (.A1(_07928_),
    .A2(_07942_),
    .B1(_07944_),
    .Y(_00378_));
 sky130_fd_sc_hd__a21o_1 _12454_ (.A1(_09093_),
    .A2(_09492_),
    .B1(_09491_),
    .X(_07945_));
 sky130_fd_sc_hd__a21oi_1 _12455_ (.A1(_09494_),
    .A2(_07945_),
    .B1(_09493_),
    .Y(_07946_));
 sky130_fd_sc_hd__xor2_1 _12456_ (.A(_09496_),
    .B(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__nor2_1 _12457_ (.A(done),
    .B(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__a21oi_1 _12458_ (.A1(\w[63][4] ),
    .A2(done),
    .B1(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__nand2_1 _12460_ (.A(message[59]),
    .B(_07928_),
    .Y(_07951_));
 sky130_fd_sc_hd__o21ai_0 _12461_ (.A1(_07928_),
    .A2(_07949_),
    .B1(_07951_),
    .Y(_00379_));
 sky130_fd_sc_hd__a21o_1 _12462_ (.A1(_09094_),
    .A2(_09494_),
    .B1(_09493_),
    .X(_07952_));
 sky130_fd_sc_hd__a21oi_1 _12463_ (.A1(_09496_),
    .A2(_07952_),
    .B1(_09495_),
    .Y(_07953_));
 sky130_fd_sc_hd__xor2_1 _12464_ (.A(_09498_),
    .B(_07953_),
    .X(_07954_));
 sky130_fd_sc_hd__nor2_1 _12465_ (.A(done),
    .B(_07954_),
    .Y(_07955_));
 sky130_fd_sc_hd__a21oi_1 _12466_ (.A1(\w[63][5] ),
    .A2(done),
    .B1(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__nand2_1 _12468_ (.A(message[58]),
    .B(_07928_),
    .Y(_07958_));
 sky130_fd_sc_hd__o21ai_0 _12469_ (.A1(_07928_),
    .A2(_07956_),
    .B1(_07958_),
    .Y(_00380_));
 sky130_fd_sc_hd__a21o_1 _12470_ (.A1(_09496_),
    .A2(_09493_),
    .B1(_09495_),
    .X(_07959_));
 sky130_fd_sc_hd__a21oi_1 _12471_ (.A1(_09498_),
    .A2(_07959_),
    .B1(_09497_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand4_1 _12472_ (.A(_09494_),
    .B(_09496_),
    .C(_09498_),
    .D(_07945_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand2_1 _12473_ (.A(_07960_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__xnor2_1 _12474_ (.A(_09500_),
    .B(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__nand2_1 _12475_ (.A(_07591_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__o21ai_1 _12476_ (.A1(\w[63][6] ),
    .A2(_07591_),
    .B1(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__nand2_1 _12478_ (.A(message[57]),
    .B(_07928_),
    .Y(_07967_));
 sky130_fd_sc_hd__o21ai_0 _12479_ (.A1(_07928_),
    .A2(_07965_),
    .B1(_07967_),
    .Y(_00381_));
 sky130_fd_sc_hd__and2_1 _12480_ (.A(_09498_),
    .B(_09500_),
    .X(_07968_));
 sky130_fd_sc_hd__a221oi_1 _12481_ (.A1(_09500_),
    .A2(_09497_),
    .B1(_07968_),
    .B2(_09495_),
    .C1(_09499_),
    .Y(_07969_));
 sky130_fd_sc_hd__nand3_1 _12482_ (.A(_09496_),
    .B(_07952_),
    .C(_07968_),
    .Y(_07970_));
 sky130_fd_sc_hd__nand2_1 _12483_ (.A(_07969_),
    .B(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__xnor2_1 _12484_ (.A(_09502_),
    .B(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__nand2_1 _12485_ (.A(_07591_),
    .B(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__o21ai_1 _12486_ (.A1(\w[63][7] ),
    .A2(_07591_),
    .B1(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(message[56]),
    .B(_07928_),
    .Y(_07976_));
 sky130_fd_sc_hd__o21ai_0 _12489_ (.A1(_07928_),
    .A2(_07974_),
    .B1(_07976_),
    .Y(_00382_));
 sky130_fd_sc_hd__a21o_1 _12490_ (.A1(_09500_),
    .A2(_07962_),
    .B1(_09499_),
    .X(_07977_));
 sky130_fd_sc_hd__a21oi_1 _12491_ (.A1(_09502_),
    .A2(_07977_),
    .B1(_09501_),
    .Y(_07978_));
 sky130_fd_sc_hd__xor2_1 _12492_ (.A(_09504_),
    .B(_07978_),
    .X(_07979_));
 sky130_fd_sc_hd__nor2_1 _12493_ (.A(done),
    .B(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__a21oi_1 _12494_ (.A1(\w[63][8] ),
    .A2(done),
    .B1(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__nand2_1 _12496_ (.A(message[55]),
    .B(_07928_),
    .Y(_07983_));
 sky130_fd_sc_hd__o21ai_0 _12497_ (.A1(_07928_),
    .A2(_07981_),
    .B1(_07983_),
    .Y(_00383_));
 sky130_fd_sc_hd__a21o_1 _12499_ (.A1(_09504_),
    .A2(_09501_),
    .B1(_09503_),
    .X(_07985_));
 sky130_fd_sc_hd__a31oi_1 _12500_ (.A1(_09502_),
    .A2(_09504_),
    .A3(_07971_),
    .B1(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__xor2_1 _12501_ (.A(_09506_),
    .B(_07986_),
    .X(_07987_));
 sky130_fd_sc_hd__nand2_1 _12502_ (.A(_07591_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__o21ai_1 _12503_ (.A1(\w[63][9] ),
    .A2(_07591_),
    .B1(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__nand2_1 _12505_ (.A(message[54]),
    .B(_07928_),
    .Y(_07991_));
 sky130_fd_sc_hd__o21ai_0 _12506_ (.A1(_07928_),
    .A2(_07989_),
    .B1(_07991_),
    .Y(_00384_));
 sky130_fd_sc_hd__a21oi_1 _12507_ (.A1(_09502_),
    .A2(_09499_),
    .B1(_09501_),
    .Y(_07992_));
 sky130_fd_sc_hd__nand2_1 _12508_ (.A(_09504_),
    .B(_09506_),
    .Y(_07993_));
 sky130_fd_sc_hd__a21oi_1 _12509_ (.A1(_09506_),
    .A2(_09503_),
    .B1(_09505_),
    .Y(_07994_));
 sky130_fd_sc_hd__o21ai_0 _12510_ (.A1(_07992_),
    .A2(_07993_),
    .B1(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__and2_1 _12511_ (.A(_09508_),
    .B(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__nand3_1 _12512_ (.A(_09502_),
    .B(_09504_),
    .C(_09506_),
    .Y(_07997_));
 sky130_fd_sc_hd__inv_1 _12513_ (.A(_09508_),
    .Y(_07998_));
 sky130_fd_sc_hd__inv_1 _12514_ (.A(_09500_),
    .Y(_07999_));
 sky130_fd_sc_hd__a2111oi_1 _12515_ (.A1(_07960_),
    .A2(_07961_),
    .B1(_07997_),
    .C1(_07998_),
    .D1(_07999_),
    .Y(_08000_));
 sky130_fd_sc_hd__nor2_1 _12516_ (.A(_07996_),
    .B(_08000_),
    .Y(_08001_));
 sky130_fd_sc_hd__nand2_1 _12517_ (.A(_09500_),
    .B(_07962_),
    .Y(_08002_));
 sky130_fd_sc_hd__nor2_1 _12518_ (.A(_08002_),
    .B(_07997_),
    .Y(_08003_));
 sky130_fd_sc_hd__or3_1 _12519_ (.A(_09508_),
    .B(_07995_),
    .C(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__and2_1 _12520_ (.A(\w[63][10] ),
    .B(done),
    .X(_08005_));
 sky130_fd_sc_hd__a31oi_2 _12521_ (.A1(_07591_),
    .A2(_08001_),
    .A3(_08004_),
    .B1(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__nand2_1 _12524_ (.A(message[53]),
    .B(_07928_),
    .Y(_08009_));
 sky130_fd_sc_hd__o21ai_0 _12525_ (.A1(_07928_),
    .A2(_08006_),
    .B1(_08009_),
    .Y(_00354_));
 sky130_fd_sc_hd__a21o_1 _12526_ (.A1(_09508_),
    .A2(_09505_),
    .B1(_09507_),
    .X(_08010_));
 sky130_fd_sc_hd__a31oi_1 _12527_ (.A1(_09496_),
    .A2(_07952_),
    .A3(_07968_),
    .B1(_07985_),
    .Y(_08011_));
 sky130_fd_sc_hd__o21a_1 _12528_ (.A1(_09502_),
    .A2(_09501_),
    .B1(_09504_),
    .X(_08012_));
 sky130_fd_sc_hd__o211ai_1 _12529_ (.A1(_09503_),
    .A2(_08012_),
    .B1(_09506_),
    .C1(_09508_),
    .Y(_08013_));
 sky130_fd_sc_hd__a21oi_1 _12530_ (.A1(_07969_),
    .A2(_08011_),
    .B1(_08013_),
    .Y(_08014_));
 sky130_fd_sc_hd__or2_2 _12531_ (.A(_08010_),
    .B(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__xnor2_1 _12532_ (.A(_09510_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand2_1 _12533_ (.A(_07591_),
    .B(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__o21ai_1 _12534_ (.A1(\w[63][11] ),
    .A2(_07591_),
    .B1(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand2_1 _12536_ (.A(message[52]),
    .B(_07928_),
    .Y(_08020_));
 sky130_fd_sc_hd__o21ai_0 _12537_ (.A1(_07928_),
    .A2(_08018_),
    .B1(_08020_),
    .Y(_00355_));
 sky130_fd_sc_hd__o31ai_1 _12538_ (.A1(_09507_),
    .A2(_07996_),
    .A3(_08000_),
    .B1(_09510_),
    .Y(_08021_));
 sky130_fd_sc_hd__nand2b_1 _12539_ (.A_N(_09509_),
    .B(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__xnor2_1 _12540_ (.A(_09512_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__nor2_1 _12541_ (.A(done),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__a21oi_1 _12542_ (.A1(\w[63][12] ),
    .A2(done),
    .B1(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__nand2_1 _12544_ (.A(message[51]),
    .B(_07928_),
    .Y(_08027_));
 sky130_fd_sc_hd__o21ai_0 _12545_ (.A1(_07928_),
    .A2(_08025_),
    .B1(_08027_),
    .Y(_00356_));
 sky130_fd_sc_hd__a21o_1 _12546_ (.A1(_09510_),
    .A2(_08015_),
    .B1(_09509_),
    .X(_08028_));
 sky130_fd_sc_hd__a21oi_1 _12547_ (.A1(_09512_),
    .A2(_08028_),
    .B1(_09511_),
    .Y(_08029_));
 sky130_fd_sc_hd__xnor2_1 _12548_ (.A(_09514_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__mux2i_2 _12549_ (.A0(\w[63][13] ),
    .A1(_08030_),
    .S(_07591_),
    .Y(_08031_));
 sky130_fd_sc_hd__nand2_1 _12551_ (.A(message[50]),
    .B(_07928_),
    .Y(_08033_));
 sky130_fd_sc_hd__o21ai_0 _12552_ (.A1(_07928_),
    .A2(_08031_),
    .B1(_08033_),
    .Y(_00357_));
 sky130_fd_sc_hd__nor2_1 _12553_ (.A(_09509_),
    .B(_09511_),
    .Y(_08034_));
 sky130_fd_sc_hd__nor2_1 _12554_ (.A(_09512_),
    .B(_09511_),
    .Y(_08035_));
 sky130_fd_sc_hd__a21oi_1 _12555_ (.A1(_08021_),
    .A2(_08034_),
    .B1(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__a21oi_1 _12556_ (.A1(_09514_),
    .A2(_08036_),
    .B1(_09513_),
    .Y(_08037_));
 sky130_fd_sc_hd__xnor2_1 _12557_ (.A(_09516_),
    .B(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__mux2i_2 _12558_ (.A0(\w[63][14] ),
    .A1(_08038_),
    .S(_07591_),
    .Y(_08039_));
 sky130_fd_sc_hd__nand2_1 _12560_ (.A(message[49]),
    .B(_07928_),
    .Y(_08041_));
 sky130_fd_sc_hd__o21ai_0 _12561_ (.A1(_07928_),
    .A2(_08039_),
    .B1(_08041_),
    .Y(_00358_));
 sky130_fd_sc_hd__a21o_1 _12562_ (.A1(_09512_),
    .A2(_09509_),
    .B1(_09511_),
    .X(_08042_));
 sky130_fd_sc_hd__a21o_1 _12563_ (.A1(_09514_),
    .A2(_08042_),
    .B1(_09513_),
    .X(_08043_));
 sky130_fd_sc_hd__and4_1 _12564_ (.A(_09510_),
    .B(_09512_),
    .C(_09514_),
    .D(_09516_),
    .X(_08044_));
 sky130_fd_sc_hd__a221o_1 _12565_ (.A1(_09516_),
    .A2(_08043_),
    .B1(_08044_),
    .B2(_08010_),
    .C1(_09515_),
    .X(_08045_));
 sky130_fd_sc_hd__o2111ai_1 _12566_ (.A1(_09503_),
    .A2(_08012_),
    .B1(_08044_),
    .C1(_09508_),
    .D1(_09506_),
    .Y(_08046_));
 sky130_fd_sc_hd__a21oi_1 _12567_ (.A1(_07969_),
    .A2(_08011_),
    .B1(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__o21a_1 _12568_ (.A1(_08045_),
    .A2(_08047_),
    .B1(_09518_),
    .X(_08048_));
 sky130_fd_sc_hd__nor3_1 _12569_ (.A(_09518_),
    .B(_08045_),
    .C(_08047_),
    .Y(_08049_));
 sky130_fd_sc_hd__o21ai_0 _12570_ (.A1(_08048_),
    .A2(_08049_),
    .B1(_07591_),
    .Y(_08050_));
 sky130_fd_sc_hd__o21ai_1 _12571_ (.A1(\w[63][15] ),
    .A2(_07591_),
    .B1(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__nand2_1 _12573_ (.A(message[48]),
    .B(_07928_),
    .Y(_08053_));
 sky130_fd_sc_hd__o21ai_0 _12574_ (.A1(_07928_),
    .A2(_08051_),
    .B1(_08053_),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_1 _12575_ (.A(_09518_),
    .B(_08044_),
    .Y(_08054_));
 sky130_fd_sc_hd__o21a_1 _12576_ (.A1(_09516_),
    .A2(_09515_),
    .B1(_09518_),
    .X(_08055_));
 sky130_fd_sc_hd__nand2_1 _12577_ (.A(_09512_),
    .B(_09514_),
    .Y(_08056_));
 sky130_fd_sc_hd__a21oi_1 _12578_ (.A1(_09510_),
    .A2(_09507_),
    .B1(_09509_),
    .Y(_08057_));
 sky130_fd_sc_hd__a2111oi_0 _12579_ (.A1(_09514_),
    .A2(_09511_),
    .B1(_09513_),
    .C1(_09515_),
    .D1(_09517_),
    .Y(_08058_));
 sky130_fd_sc_hd__o21ai_0 _12580_ (.A1(_08056_),
    .A2(_08057_),
    .B1(_08058_),
    .Y(_08059_));
 sky130_fd_sc_hd__o21ai_0 _12581_ (.A1(_09517_),
    .A2(_08055_),
    .B1(_08059_),
    .Y(_08060_));
 sky130_fd_sc_hd__o21ai_0 _12582_ (.A1(_08001_),
    .A2(_08054_),
    .B1(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__xnor2_1 _12583_ (.A(_09520_),
    .B(_08061_),
    .Y(_08062_));
 sky130_fd_sc_hd__nand2_1 _12584_ (.A(_07591_),
    .B(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__o21ai_1 _12585_ (.A1(\w[63][16] ),
    .A2(_07591_),
    .B1(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__nand2_1 _12587_ (.A(message[47]),
    .B(_07928_),
    .Y(_08066_));
 sky130_fd_sc_hd__o21ai_0 _12588_ (.A1(_07928_),
    .A2(_08064_),
    .B1(_08066_),
    .Y(_00360_));
 sky130_fd_sc_hd__inv_1 _12589_ (.A(_09519_),
    .Y(_08067_));
 sky130_fd_sc_hd__o21ai_0 _12590_ (.A1(_09517_),
    .A2(_08048_),
    .B1(_09520_),
    .Y(_08068_));
 sky130_fd_sc_hd__nand2_1 _12591_ (.A(_08067_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__xor2_1 _12592_ (.A(_09522_),
    .B(_08069_),
    .X(_08070_));
 sky130_fd_sc_hd__mux2i_2 _12593_ (.A0(\w[63][17] ),
    .A1(_08070_),
    .S(_07591_),
    .Y(_08071_));
 sky130_fd_sc_hd__nand2_1 _12595_ (.A(message[46]),
    .B(_07928_),
    .Y(_08073_));
 sky130_fd_sc_hd__o21ai_0 _12596_ (.A1(_07928_),
    .A2(_08071_),
    .B1(_08073_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_1 _12597_ (.A(_09520_),
    .B(_09522_),
    .Y(_08074_));
 sky130_fd_sc_hd__nor2_1 _12598_ (.A(_08054_),
    .B(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__o21ai_0 _12599_ (.A1(_07996_),
    .A2(_08000_),
    .B1(_08075_),
    .Y(_08076_));
 sky130_fd_sc_hd__a21o_1 _12600_ (.A1(_09522_),
    .A2(_09519_),
    .B1(_09521_),
    .X(_08077_));
 sky130_fd_sc_hd__o21ba_2 _12601_ (.A1(_08060_),
    .A2(_08074_),
    .B1_N(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__nand2_1 _12602_ (.A(_08076_),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__xnor2_1 _12603_ (.A(_09524_),
    .B(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__nor2_1 _12604_ (.A(done),
    .B(_08080_),
    .Y(_08081_));
 sky130_fd_sc_hd__a21oi_1 _12605_ (.A1(\w[63][18] ),
    .A2(done),
    .B1(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__nand2_1 _12607_ (.A(message[45]),
    .B(_07928_),
    .Y(_08084_));
 sky130_fd_sc_hd__o21ai_0 _12608_ (.A1(_07928_),
    .A2(_08082_),
    .B1(_08084_),
    .Y(_00362_));
 sky130_fd_sc_hd__nor3_1 _12610_ (.A(_09519_),
    .B(_09521_),
    .C(_09523_),
    .Y(_08086_));
 sky130_fd_sc_hd__or2_2 _12611_ (.A(_09522_),
    .B(_09521_),
    .X(_08087_));
 sky130_fd_sc_hd__a21oi_1 _12612_ (.A1(_09524_),
    .A2(_08087_),
    .B1(_09523_),
    .Y(_08088_));
 sky130_fd_sc_hd__a21oi_1 _12613_ (.A1(_08068_),
    .A2(_08086_),
    .B1(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__xor2_1 _12614_ (.A(_09526_),
    .B(_08089_),
    .X(_08090_));
 sky130_fd_sc_hd__mux2i_2 _12615_ (.A0(\w[63][19] ),
    .A1(_08090_),
    .S(_07591_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand2_1 _12617_ (.A(message[44]),
    .B(_07928_),
    .Y(_08093_));
 sky130_fd_sc_hd__o21ai_0 _12618_ (.A1(_07928_),
    .A2(_08091_),
    .B1(_08093_),
    .Y(_00363_));
 sky130_fd_sc_hd__and3_1 _12619_ (.A(_09522_),
    .B(_09524_),
    .C(_09526_),
    .X(_08094_));
 sky130_fd_sc_hd__nand2_1 _12620_ (.A(_09520_),
    .B(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__a21o_1 _12621_ (.A1(_09524_),
    .A2(_08077_),
    .B1(_09523_),
    .X(_08096_));
 sky130_fd_sc_hd__a21oi_1 _12622_ (.A1(_09526_),
    .A2(_08096_),
    .B1(_09525_),
    .Y(_08097_));
 sky130_fd_sc_hd__o21a_1 _12623_ (.A1(_08060_),
    .A2(_08095_),
    .B1(_08097_),
    .X(_08098_));
 sky130_fd_sc_hd__o31ai_1 _12624_ (.A1(_08001_),
    .A2(_08054_),
    .A3(_08095_),
    .B1(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__xnor2_1 _12625_ (.A(_09528_),
    .B(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__nand2_1 _12626_ (.A(_07591_),
    .B(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__o21ai_1 _12627_ (.A1(\w[63][20] ),
    .A2(_07591_),
    .B1(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__nand2_1 _12630_ (.A(message[43]),
    .B(_07928_),
    .Y(_08105_));
 sky130_fd_sc_hd__o21ai_0 _12631_ (.A1(_07928_),
    .A2(_08102_),
    .B1(_08105_),
    .Y(_00365_));
 sky130_fd_sc_hd__a21o_1 _12632_ (.A1(_09524_),
    .A2(_09521_),
    .B1(_09523_),
    .X(_08106_));
 sky130_fd_sc_hd__a21oi_1 _12633_ (.A1(_09526_),
    .A2(_08106_),
    .B1(_09525_),
    .Y(_08107_));
 sky130_fd_sc_hd__nor2_1 _12634_ (.A(_09519_),
    .B(_09527_),
    .Y(_08108_));
 sky130_fd_sc_hd__nor2_1 _12635_ (.A(_09527_),
    .B(_08094_),
    .Y(_08109_));
 sky130_fd_sc_hd__nand2_1 _12636_ (.A(_08107_),
    .B(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__o21ai_0 _12637_ (.A1(_09528_),
    .A2(_09527_),
    .B1(_08110_),
    .Y(_08111_));
 sky130_fd_sc_hd__a31oi_1 _12638_ (.A1(_08068_),
    .A2(_08107_),
    .A3(_08108_),
    .B1(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__xor2_1 _12639_ (.A(_09530_),
    .B(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__mux2i_2 _12640_ (.A0(\w[63][21] ),
    .A1(_08113_),
    .S(_07591_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_1 _12642_ (.A(message[42]),
    .B(_07928_),
    .Y(_08116_));
 sky130_fd_sc_hd__o21ai_0 _12643_ (.A1(_07928_),
    .A2(_08114_),
    .B1(_08116_),
    .Y(_00366_));
 sky130_fd_sc_hd__a21o_1 _12645_ (.A1(_09526_),
    .A2(_09523_),
    .B1(_09525_),
    .X(_08118_));
 sky130_fd_sc_hd__a21o_1 _12646_ (.A1(_09528_),
    .A2(_08118_),
    .B1(_09527_),
    .X(_08119_));
 sky130_fd_sc_hd__a21o_1 _12647_ (.A1(_09530_),
    .A2(_08119_),
    .B1(_09529_),
    .X(_08120_));
 sky130_fd_sc_hd__nand4_1 _12648_ (.A(_09524_),
    .B(_09526_),
    .C(_09528_),
    .D(_09530_),
    .Y(_08121_));
 sky130_fd_sc_hd__a21oi_1 _12649_ (.A1(_08076_),
    .A2(_08078_),
    .B1(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__nor2_1 _12650_ (.A(_08120_),
    .B(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__xnor2_1 _12651_ (.A(_09532_),
    .B(_08123_),
    .Y(_08124_));
 sky130_fd_sc_hd__mux2i_2 _12652_ (.A0(\w[63][22] ),
    .A1(_08124_),
    .S(_07591_),
    .Y(_08125_));
 sky130_fd_sc_hd__nand2_1 _12654_ (.A(message[41]),
    .B(_07928_),
    .Y(_08127_));
 sky130_fd_sc_hd__o21ai_0 _12655_ (.A1(_07928_),
    .A2(_08125_),
    .B1(_08127_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand3_1 _12656_ (.A(_09528_),
    .B(_09530_),
    .C(_09532_),
    .Y(_08128_));
 sky130_fd_sc_hd__a21o_1 _12657_ (.A1(_09530_),
    .A2(_09527_),
    .B1(_09529_),
    .X(_08129_));
 sky130_fd_sc_hd__a21oi_1 _12658_ (.A1(_09532_),
    .A2(_08129_),
    .B1(_09531_),
    .Y(_08130_));
 sky130_fd_sc_hd__o21ai_0 _12659_ (.A1(_08107_),
    .A2(_08128_),
    .B1(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__nand2_1 _12660_ (.A(_09520_),
    .B(_09517_),
    .Y(_08132_));
 sky130_fd_sc_hd__nand2_1 _12661_ (.A(_08067_),
    .B(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__o21ai_0 _12662_ (.A1(_09518_),
    .A2(_09517_),
    .B1(_09520_),
    .Y(_08134_));
 sky130_fd_sc_hd__and3_1 _12663_ (.A(_09528_),
    .B(_09530_),
    .C(_09532_),
    .X(_08135_));
 sky130_fd_sc_hd__nand2_1 _12664_ (.A(_08094_),
    .B(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__a21oi_1 _12665_ (.A1(_08067_),
    .A2(_08134_),
    .B1(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__o31ai_1 _12666_ (.A1(_08045_),
    .A2(_08047_),
    .A3(_08133_),
    .B1(_08137_),
    .Y(_08138_));
 sky130_fd_sc_hd__nor2b_1 _12667_ (.A(_08131_),
    .B_N(_08138_),
    .Y(_08139_));
 sky130_fd_sc_hd__xor2_1 _12668_ (.A(_09534_),
    .B(_08139_),
    .X(_08140_));
 sky130_fd_sc_hd__nand2_1 _12669_ (.A(_07591_),
    .B(_08140_),
    .Y(_08141_));
 sky130_fd_sc_hd__o21ai_1 _12670_ (.A1(\w[63][23] ),
    .A2(_07591_),
    .B1(_08141_),
    .Y(_08142_));
 sky130_fd_sc_hd__nand2_1 _12672_ (.A(message[40]),
    .B(_07928_),
    .Y(_08144_));
 sky130_fd_sc_hd__o21ai_0 _12673_ (.A1(_07928_),
    .A2(_08142_),
    .B1(_08144_),
    .Y(_00368_));
 sky130_fd_sc_hd__a21boi_1 _12675_ (.A1(_08099_),
    .A2(_08135_),
    .B1_N(_08130_),
    .Y(_08146_));
 sky130_fd_sc_hd__nor4b_1 _12676_ (.A(_09536_),
    .B(done),
    .C(_08146_),
    .D_N(_09534_),
    .Y(_08147_));
 sky130_fd_sc_hd__and4b_1 _12677_ (.A_N(_09533_),
    .B(_07591_),
    .C(_08146_),
    .D(_09536_),
    .X(_08148_));
 sky130_fd_sc_hd__nor4b_1 _12678_ (.A(_09534_),
    .B(_09533_),
    .C(done),
    .D_N(_09536_),
    .Y(_08149_));
 sky130_fd_sc_hd__nor3b_1 _12679_ (.A(_09536_),
    .B(done),
    .C_N(_09533_),
    .Y(_08150_));
 sky130_fd_sc_hd__a211o_1 _12680_ (.A1(\w[63][24] ),
    .A2(done),
    .B1(_08149_),
    .C1(_08150_),
    .X(_08151_));
 sky130_fd_sc_hd__nor3_2 _12681_ (.A(_08147_),
    .B(_08148_),
    .C(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__nand2_1 _12683_ (.A(message[39]),
    .B(_07928_),
    .Y(_08154_));
 sky130_fd_sc_hd__o21ai_1 _12684_ (.A1(_07928_),
    .A2(_08152_),
    .B1(_08154_),
    .Y(_00369_));
 sky130_fd_sc_hd__inv_1 _12685_ (.A(_09538_),
    .Y(_08155_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(_09534_),
    .B(_09536_),
    .Y(_08156_));
 sky130_fd_sc_hd__a21oi_1 _12687_ (.A1(_09536_),
    .A2(_09533_),
    .B1(_09535_),
    .Y(_08157_));
 sky130_fd_sc_hd__o21ai_0 _12688_ (.A1(_08139_),
    .A2(_08156_),
    .B1(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__xnor2_1 _12689_ (.A(_08155_),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__mux2i_2 _12690_ (.A0(\w[63][25] ),
    .A1(_08159_),
    .S(_07591_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand2_1 _12692_ (.A(message[38]),
    .B(_07928_),
    .Y(_08162_));
 sky130_fd_sc_hd__o21ai_0 _12693_ (.A1(_07928_),
    .A2(_08160_),
    .B1(_08162_),
    .Y(_00370_));
 sky130_fd_sc_hd__nor2_1 _12694_ (.A(_08155_),
    .B(_08156_),
    .Y(_08163_));
 sky130_fd_sc_hd__nand2_1 _12695_ (.A(_09536_),
    .B(_09538_),
    .Y(_08164_));
 sky130_fd_sc_hd__a21oi_1 _12696_ (.A1(_09534_),
    .A2(_09531_),
    .B1(_09533_),
    .Y(_08165_));
 sky130_fd_sc_hd__a21oi_1 _12697_ (.A1(_09538_),
    .A2(_09535_),
    .B1(_09537_),
    .Y(_08166_));
 sky130_fd_sc_hd__o21ai_0 _12698_ (.A1(_08164_),
    .A2(_08165_),
    .B1(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__a31o_2 _12699_ (.A1(_09532_),
    .A2(_08120_),
    .A3(_08163_),
    .B1(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__a31oi_1 _12700_ (.A1(_09532_),
    .A2(_08122_),
    .A3(_08163_),
    .B1(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__xnor2_1 _12701_ (.A(_09540_),
    .B(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__mux2i_2 _12702_ (.A0(\w[63][26] ),
    .A1(_08170_),
    .S(_07591_),
    .Y(_08171_));
 sky130_fd_sc_hd__nand2_1 _12704_ (.A(message[37]),
    .B(_07928_),
    .Y(_08173_));
 sky130_fd_sc_hd__o21ai_0 _12705_ (.A1(_07928_),
    .A2(_08171_),
    .B1(_08173_),
    .Y(_00371_));
 sky130_fd_sc_hd__nand2_1 _12706_ (.A(_09540_),
    .B(_08163_),
    .Y(_08174_));
 sky130_fd_sc_hd__o21bai_1 _12707_ (.A1(_08155_),
    .A2(_08157_),
    .B1_N(_09537_),
    .Y(_08175_));
 sky130_fd_sc_hd__a21o_1 _12708_ (.A1(_09540_),
    .A2(_08175_),
    .B1(_09539_),
    .X(_08176_));
 sky130_fd_sc_hd__nor2_1 _12709_ (.A(_09542_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__o21ai_0 _12710_ (.A1(_08139_),
    .A2(_08174_),
    .B1(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__and2_1 _12711_ (.A(_09540_),
    .B(_09542_),
    .X(_08179_));
 sky130_fd_sc_hd__nand2_1 _12712_ (.A(_08163_),
    .B(_08179_),
    .Y(_08180_));
 sky130_fd_sc_hd__a32oi_1 _12713_ (.A1(_08131_),
    .A2(_08163_),
    .A3(_08179_),
    .B1(_08176_),
    .B2(_09542_),
    .Y(_08181_));
 sky130_fd_sc_hd__o21ai_0 _12714_ (.A1(_08138_),
    .A2(_08180_),
    .B1(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__nor2_1 _12715_ (.A(done),
    .B(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__a22oi_1 _12716_ (.A1(\w[63][27] ),
    .A2(done),
    .B1(_08178_),
    .B2(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__nand2_1 _12718_ (.A(message[36]),
    .B(_07928_),
    .Y(_08186_));
 sky130_fd_sc_hd__o21ai_0 _12719_ (.A1(_07928_),
    .A2(_08184_),
    .B1(_08186_),
    .Y(_00372_));
 sky130_fd_sc_hd__nand2b_1 _12721_ (.A_N(_08146_),
    .B(_08163_),
    .Y(_08188_));
 sky130_fd_sc_hd__a21oi_1 _12722_ (.A1(_09542_),
    .A2(_09539_),
    .B1(_09541_),
    .Y(_08189_));
 sky130_fd_sc_hd__nand4_1 _12723_ (.A(_09545_),
    .B(_07591_),
    .C(_08166_),
    .D(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__a31oi_1 _12724_ (.A1(_09536_),
    .A2(_09538_),
    .A3(_09533_),
    .B1(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__inv_1 _12725_ (.A(_09541_),
    .Y(_08192_));
 sky130_fd_sc_hd__o21ai_0 _12726_ (.A1(_09540_),
    .A2(_09539_),
    .B1(_09542_),
    .Y(_08193_));
 sky130_fd_sc_hd__nor2b_1 _12727_ (.A(_08166_),
    .B_N(_09540_),
    .Y(_08194_));
 sky130_fd_sc_hd__o21ai_0 _12728_ (.A1(_09539_),
    .A2(_08194_),
    .B1(_09542_),
    .Y(_08195_));
 sky130_fd_sc_hd__a21oi_1 _12729_ (.A1(_08192_),
    .A2(_08195_),
    .B1(_09545_),
    .Y(_08196_));
 sky130_fd_sc_hd__a311o_1 _12730_ (.A1(_09545_),
    .A2(_08192_),
    .A3(_08193_),
    .B1(_08196_),
    .C1(done),
    .X(_08197_));
 sky130_fd_sc_hd__o21a_1 _12731_ (.A1(\w[63][28] ),
    .A2(_07591_),
    .B1(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__nand2_1 _12732_ (.A(_09540_),
    .B(_09542_),
    .Y(_08199_));
 sky130_fd_sc_hd__nor3_1 _12733_ (.A(_09545_),
    .B(done),
    .C(_08199_),
    .Y(_08200_));
 sky130_fd_sc_hd__nand2_1 _12734_ (.A(_08163_),
    .B(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__nand4_1 _12735_ (.A(_09536_),
    .B(_09538_),
    .C(_09533_),
    .D(_08200_),
    .Y(_08202_));
 sky130_fd_sc_hd__o21ai_0 _12736_ (.A1(_08146_),
    .A2(_08201_),
    .B1(_08202_),
    .Y(_08203_));
 sky130_fd_sc_hd__a211oi_2 _12737_ (.A1(_08188_),
    .A2(_08191_),
    .B1(_08198_),
    .C1(_08203_),
    .Y(_08204_));
 sky130_fd_sc_hd__a21oi_1 _12738_ (.A1(_05403_),
    .A2(_07927_),
    .B1(message[35]),
    .Y(_08205_));
 sky130_fd_sc_hd__a31oi_1 _12739_ (.A1(_05403_),
    .A2(_07927_),
    .A3(_08204_),
    .B1(_08205_),
    .Y(_00373_));
 sky130_fd_sc_hd__o211ai_1 _12740_ (.A1(_08138_),
    .A2(_08180_),
    .B1(_08181_),
    .C1(_08192_),
    .Y(_08206_));
 sky130_fd_sc_hd__a21oi_1 _12741_ (.A1(_09545_),
    .A2(_08206_),
    .B1(_09544_),
    .Y(_08207_));
 sky130_fd_sc_hd__xnor2_1 _12742_ (.A(_09549_),
    .B(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__mux2i_2 _12743_ (.A0(\w[63][29] ),
    .A1(_08208_),
    .S(_07591_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand2_1 _12745_ (.A(message[34]),
    .B(_07928_),
    .Y(_08211_));
 sky130_fd_sc_hd__o21ai_0 _12746_ (.A1(_07928_),
    .A2(_08209_),
    .B1(_08211_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _12747_ (.A(_09532_),
    .B(_08163_),
    .Y(_08212_));
 sky130_fd_sc_hd__a2111oi_0 _12748_ (.A1(_08076_),
    .A2(_08078_),
    .B1(_08121_),
    .C1(_08212_),
    .D1(_08199_),
    .Y(_08213_));
 sky130_fd_sc_hd__nor2_1 _12749_ (.A(_09544_),
    .B(_09548_),
    .Y(_08214_));
 sky130_fd_sc_hd__nand2_1 _12750_ (.A(_08189_),
    .B(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__a21o_1 _12751_ (.A1(_08168_),
    .A2(_08179_),
    .B1(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__o21ai_0 _12752_ (.A1(_09545_),
    .A2(_09544_),
    .B1(_09549_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2b_1 _12753_ (.A_N(_09548_),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__o21ai_0 _12754_ (.A1(_08213_),
    .A2(_08216_),
    .B1(_08218_),
    .Y(_08219_));
 sky130_fd_sc_hd__xnor2_1 _12755_ (.A(_09552_),
    .B(_08219_),
    .Y(_08220_));
 sky130_fd_sc_hd__mux2i_2 _12756_ (.A0(\w[63][30] ),
    .A1(_08220_),
    .S(_07591_),
    .Y(_08221_));
 sky130_fd_sc_hd__nand2_1 _12758_ (.A(message[33]),
    .B(_07928_),
    .Y(_08223_));
 sky130_fd_sc_hd__o21ai_0 _12759_ (.A1(_07928_),
    .A2(_08221_),
    .B1(_08223_),
    .Y(_00376_));
 sky130_fd_sc_hd__xnor2_1 _12760_ (.A(\w_new_calc2.temp1[31] ),
    .B(_09344_),
    .Y(_08224_));
 sky130_fd_sc_hd__xnor2_1 _12761_ (.A(\w_new_calc2.temp2[31] ),
    .B(_09341_),
    .Y(_08225_));
 sky130_fd_sc_hd__xnor2_1 _12762_ (.A(_08224_),
    .B(_08225_),
    .Y(_08226_));
 sky130_fd_sc_hd__mux4_2 _12763_ (.A0(\w[1][31] ),
    .A1(\w[3][31] ),
    .A2(\w[9][31] ),
    .A3(\w[11][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[3] ),
    .X(_08227_));
 sky130_fd_sc_hd__mux4_2 _12764_ (.A0(\w[5][31] ),
    .A1(\w[7][31] ),
    .A2(\w[13][31] ),
    .A3(\w[15][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[3] ),
    .X(_08228_));
 sky130_fd_sc_hd__mux4_2 _12765_ (.A0(\w[33][31] ),
    .A1(\w[35][31] ),
    .A2(\w[41][31] ),
    .A3(\w[43][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[3] ),
    .X(_08229_));
 sky130_fd_sc_hd__mux4_2 _12766_ (.A0(\w[37][31] ),
    .A1(\w[39][31] ),
    .A2(\w[45][31] ),
    .A3(\w[47][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[3] ),
    .X(_08230_));
 sky130_fd_sc_hd__mux4_2 _12767_ (.A0(_08227_),
    .A1(_08228_),
    .A2(_08229_),
    .A3(_08230_),
    .S0(\count16_2[2] ),
    .S1(\count16_2[5] ),
    .X(_08231_));
 sky130_fd_sc_hd__mux4_2 _12768_ (.A0(\w[17][31] ),
    .A1(\w[19][31] ),
    .A2(\w[21][31] ),
    .A3(\w[23][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_08232_));
 sky130_fd_sc_hd__mux4_2 _12769_ (.A0(\w[25][31] ),
    .A1(\w[27][31] ),
    .A2(\w[29][31] ),
    .A3(\w[31][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_08233_));
 sky130_fd_sc_hd__mux4_2 _12770_ (.A0(\w[49][31] ),
    .A1(\w[51][31] ),
    .A2(\w[53][31] ),
    .A3(\w[55][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_08234_));
 sky130_fd_sc_hd__mux4_2 _12771_ (.A0(\w[57][31] ),
    .A1(\w[59][31] ),
    .A2(\w[61][31] ),
    .A3(\w[63][31] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_08235_));
 sky130_fd_sc_hd__mux4_2 _12772_ (.A0(_08232_),
    .A1(_08233_),
    .A2(_08234_),
    .A3(_08235_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[5] ),
    .X(_08236_));
 sky130_fd_sc_hd__mux2i_1 _12773_ (.A0(_08231_),
    .A1(_08236_),
    .S(\count16_2[4] ),
    .Y(_08237_));
 sky130_fd_sc_hd__mux4_2 _12774_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[16][31] ),
    .A3(\w[20][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[4] ),
    .X(_08238_));
 sky130_fd_sc_hd__mux4_2 _12775_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[48][31] ),
    .A3(\w[52][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[4] ),
    .X(_08239_));
 sky130_fd_sc_hd__mux4_2 _12776_ (.A0(\w[2][31] ),
    .A1(\w[6][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[4] ),
    .X(_08240_));
 sky130_fd_sc_hd__mux4_2 _12777_ (.A0(\w[34][31] ),
    .A1(\w[38][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[4] ),
    .X(_08241_));
 sky130_fd_sc_hd__mux4_2 _12778_ (.A0(_08238_),
    .A1(_08239_),
    .A2(_08240_),
    .A3(_08241_),
    .S0(\count7_2[5] ),
    .S1(\count7_2[1] ),
    .X(_08242_));
 sky130_fd_sc_hd__mux4_2 _12779_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_08243_));
 sky130_fd_sc_hd__mux4_2 _12780_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_08244_));
 sky130_fd_sc_hd__mux4_2 _12781_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_08245_));
 sky130_fd_sc_hd__mux4_2 _12782_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_08246_));
 sky130_fd_sc_hd__mux4_2 _12783_ (.A0(_08243_),
    .A1(_08244_),
    .A2(_08245_),
    .A3(_08246_),
    .S0(\count7_2[5] ),
    .S1(\count7_2[4] ),
    .X(_08247_));
 sky130_fd_sc_hd__mux2i_1 _12784_ (.A0(_08242_),
    .A1(_08247_),
    .S(\count7_2[3] ),
    .Y(_08248_));
 sky130_fd_sc_hd__xnor2_1 _12785_ (.A(_08237_),
    .B(_08248_),
    .Y(_08249_));
 sky130_fd_sc_hd__xnor2_1 _12786_ (.A(_08226_),
    .B(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__o2111ai_1 _12787_ (.A1(_08138_),
    .A2(_08180_),
    .B1(_08181_),
    .C1(_08214_),
    .D1(_08192_),
    .Y(_08251_));
 sky130_fd_sc_hd__a31oi_1 _12788_ (.A1(_09552_),
    .A2(_08218_),
    .A3(_08251_),
    .B1(_09551_),
    .Y(_08252_));
 sky130_fd_sc_hd__xnor2_1 _12789_ (.A(_08250_),
    .B(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__mux2i_4 _12790_ (.A0(\w[63][31] ),
    .A1(_08253_),
    .S(_07591_),
    .Y(_08254_));
 sky130_fd_sc_hd__nand2_1 _12792_ (.A(message[32]),
    .B(_07928_),
    .Y(_08256_));
 sky130_fd_sc_hd__o21ai_1 _12793_ (.A1(_07928_),
    .A2(_08254_),
    .B1(_08256_),
    .Y(_00377_));
 sky130_fd_sc_hd__nor2b_1 _12794_ (.A(reset),
    .B_N(_09557_),
    .Y(_08257_));
 sky130_fd_sc_hd__nand2_1 _12796_ (.A(_05338_),
    .B(_08257_),
    .Y(_08259_));
 sky130_fd_sc_hd__nand2_1 _12800_ (.A(message[95]),
    .B(_08259_),
    .Y(_08263_));
 sky130_fd_sc_hd__o21ai_0 _12801_ (.A1(_07572_),
    .A2(_08259_),
    .B1(_08263_),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(message[94]),
    .B(_08259_),
    .Y(_08264_));
 sky130_fd_sc_hd__o21ai_0 _12803_ (.A1(_07577_),
    .A2(_08259_),
    .B1(_08264_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _12804_ (.A(message[93]),
    .B(_08259_),
    .Y(_08265_));
 sky130_fd_sc_hd__o21ai_0 _12805_ (.A1(_07581_),
    .A2(_08259_),
    .B1(_08265_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand2_1 _12807_ (.A(message[92]),
    .B(_08259_),
    .Y(_08267_));
 sky130_fd_sc_hd__o21ai_0 _12808_ (.A1(_07588_),
    .A2(_08259_),
    .B1(_08267_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _12809_ (.A(message[91]),
    .B(_08259_),
    .Y(_08268_));
 sky130_fd_sc_hd__o21ai_0 _12810_ (.A1(_07601_),
    .A2(_08259_),
    .B1(_08268_),
    .Y(_00411_));
 sky130_fd_sc_hd__nand2_1 _12811_ (.A(message[90]),
    .B(_08259_),
    .Y(_08269_));
 sky130_fd_sc_hd__o21ai_0 _12812_ (.A1(_07610_),
    .A2(_08259_),
    .B1(_08269_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _12813_ (.A(message[89]),
    .B(_08259_),
    .Y(_08270_));
 sky130_fd_sc_hd__o21ai_0 _12814_ (.A1(_07620_),
    .A2(_08259_),
    .B1(_08270_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _12815_ (.A(message[88]),
    .B(_08259_),
    .Y(_08271_));
 sky130_fd_sc_hd__o21ai_0 _12816_ (.A1(_07628_),
    .A2(_08259_),
    .B1(_08271_),
    .Y(_00414_));
 sky130_fd_sc_hd__nand2_1 _12817_ (.A(message[87]),
    .B(_08259_),
    .Y(_08272_));
 sky130_fd_sc_hd__o21ai_0 _12818_ (.A1(_07635_),
    .A2(_08259_),
    .B1(_08272_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _12819_ (.A(message[86]),
    .B(_08259_),
    .Y(_08273_));
 sky130_fd_sc_hd__o21ai_0 _12820_ (.A1(_07646_),
    .A2(_08259_),
    .B1(_08273_),
    .Y(_00416_));
 sky130_fd_sc_hd__nand2_1 _12822_ (.A(message[85]),
    .B(_08259_),
    .Y(_08275_));
 sky130_fd_sc_hd__o21ai_0 _12823_ (.A1(_07660_),
    .A2(_08259_),
    .B1(_08275_),
    .Y(_00386_));
 sky130_fd_sc_hd__and2_1 _12824_ (.A(_05338_),
    .B(_08257_),
    .X(_08276_));
 sky130_fd_sc_hd__nor2_1 _12826_ (.A(message[84]),
    .B(_08276_),
    .Y(_08278_));
 sky130_fd_sc_hd__a21oi_1 _12827_ (.A1(_07669_),
    .A2(_08276_),
    .B1(_08278_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _12828_ (.A(message[83]),
    .B(_08259_),
    .Y(_08279_));
 sky130_fd_sc_hd__o21ai_0 _12829_ (.A1(_07677_),
    .A2(_08259_),
    .B1(_08279_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _12830_ (.A(message[82]),
    .B(_08259_),
    .Y(_08280_));
 sky130_fd_sc_hd__o21ai_0 _12831_ (.A1(_07689_),
    .A2(_08259_),
    .B1(_08280_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _12833_ (.A(message[81]),
    .B(_08259_),
    .Y(_08282_));
 sky130_fd_sc_hd__o21ai_0 _12834_ (.A1(_07703_),
    .A2(_08259_),
    .B1(_08282_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _12835_ (.A(message[80]),
    .B(_08259_),
    .Y(_08283_));
 sky130_fd_sc_hd__o21ai_0 _12836_ (.A1(_07709_),
    .A2(_08259_),
    .B1(_08283_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_1 _12837_ (.A(message[79]),
    .B(_08259_),
    .Y(_08284_));
 sky130_fd_sc_hd__o21ai_0 _12838_ (.A1(_07715_),
    .A2(_08259_),
    .B1(_08284_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand2_1 _12839_ (.A(message[78]),
    .B(_08259_),
    .Y(_08285_));
 sky130_fd_sc_hd__o21ai_0 _12840_ (.A1(_07731_),
    .A2(_08259_),
    .B1(_08285_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _12841_ (.A(message[77]),
    .B(_08259_),
    .Y(_08286_));
 sky130_fd_sc_hd__o21ai_0 _12842_ (.A1(_07745_),
    .A2(_08259_),
    .B1(_08286_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _12843_ (.A(message[76]),
    .B(_08259_),
    .Y(_08287_));
 sky130_fd_sc_hd__o21ai_0 _12844_ (.A1(_07752_),
    .A2(_08259_),
    .B1(_08287_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _12845_ (.A(message[75]),
    .B(_08259_),
    .Y(_08288_));
 sky130_fd_sc_hd__o21ai_0 _12846_ (.A1(_07766_),
    .A2(_08259_),
    .B1(_08288_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _12847_ (.A(message[74]),
    .B(_08259_),
    .Y(_08289_));
 sky130_fd_sc_hd__o21ai_0 _12848_ (.A1(_07777_),
    .A2(_08259_),
    .B1(_08289_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _12849_ (.A(message[73]),
    .B(_08259_),
    .Y(_08290_));
 sky130_fd_sc_hd__o21ai_0 _12850_ (.A1(_07786_),
    .A2(_08259_),
    .B1(_08290_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _12851_ (.A(message[72]),
    .B(_08259_),
    .Y(_08291_));
 sky130_fd_sc_hd__o21ai_0 _12852_ (.A1(_07800_),
    .A2(_08259_),
    .B1(_08291_),
    .Y(_00400_));
 sky130_fd_sc_hd__nor2_1 _12854_ (.A(message[71]),
    .B(_08276_),
    .Y(_08293_));
 sky130_fd_sc_hd__a21oi_1 _12855_ (.A1(_07809_),
    .A2(_08276_),
    .B1(_08293_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _12856_ (.A(message[70]),
    .B(_08259_),
    .Y(_08294_));
 sky130_fd_sc_hd__o21ai_0 _12857_ (.A1(_07818_),
    .A2(_08259_),
    .B1(_08294_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _12858_ (.A(message[69]),
    .B(_08259_),
    .Y(_08295_));
 sky130_fd_sc_hd__o21ai_0 _12859_ (.A1(_07831_),
    .A2(_08259_),
    .B1(_08295_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _12860_ (.A(message[68]),
    .B(_08259_),
    .Y(_08296_));
 sky130_fd_sc_hd__o21ai_0 _12861_ (.A1(_07843_),
    .A2(_08259_),
    .B1(_08296_),
    .Y(_00404_));
 sky130_fd_sc_hd__nor2_1 _12863_ (.A(message[67]),
    .B(_08276_),
    .Y(_08298_));
 sky130_fd_sc_hd__a21oi_1 _12864_ (.A1(_07850_),
    .A2(_08276_),
    .B1(_08298_),
    .Y(_00405_));
 sky130_fd_sc_hd__nor2_1 _12865_ (.A(_07860_),
    .B(_08259_),
    .Y(_08299_));
 sky130_fd_sc_hd__a21oi_1 _12866_ (.A1(message[66]),
    .A2(_08259_),
    .B1(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__a21oi_1 _12867_ (.A1(_07859_),
    .A2(_08276_),
    .B1(_08300_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _12868_ (.A(message[65]),
    .B(_08259_),
    .Y(_08301_));
 sky130_fd_sc_hd__o21ai_0 _12869_ (.A1(_07873_),
    .A2(_08259_),
    .B1(_08301_),
    .Y(_00408_));
 sky130_fd_sc_hd__nor2_1 _12871_ (.A(message[64]),
    .B(_08276_),
    .Y(_08303_));
 sky130_fd_sc_hd__a21oi_1 _12872_ (.A1(_07925_),
    .A2(_08276_),
    .B1(_08303_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2b_1 _12873_ (.A(reset),
    .B_N(_09565_),
    .Y(_08304_));
 sky130_fd_sc_hd__nand2_1 _12874_ (.A(_05403_),
    .B(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _12877_ (.A(message[127]),
    .B(_08305_),
    .Y(_08308_));
 sky130_fd_sc_hd__o21ai_0 _12878_ (.A1(_07930_),
    .A2(_08305_),
    .B1(_08308_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _12879_ (.A(message[126]),
    .B(_08305_),
    .Y(_08309_));
 sky130_fd_sc_hd__o21ai_0 _12880_ (.A1(_07934_),
    .A2(_08305_),
    .B1(_08309_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _12881_ (.A(message[125]),
    .B(_08305_),
    .Y(_08310_));
 sky130_fd_sc_hd__o21ai_0 _12882_ (.A1(_07937_),
    .A2(_08305_),
    .B1(_08310_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _12883_ (.A(message[124]),
    .B(_08305_),
    .Y(_08311_));
 sky130_fd_sc_hd__o21ai_0 _12884_ (.A1(_07942_),
    .A2(_08305_),
    .B1(_08311_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _12885_ (.A(message[123]),
    .B(_08305_),
    .Y(_08312_));
 sky130_fd_sc_hd__o21ai_0 _12886_ (.A1(_07949_),
    .A2(_08305_),
    .B1(_08312_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _12887_ (.A(message[122]),
    .B(_08305_),
    .Y(_08313_));
 sky130_fd_sc_hd__o21ai_0 _12888_ (.A1(_07956_),
    .A2(_08305_),
    .B1(_08313_),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _12889_ (.A(message[121]),
    .B(_08305_),
    .Y(_08314_));
 sky130_fd_sc_hd__o21ai_0 _12890_ (.A1(_07965_),
    .A2(_08305_),
    .B1(_08314_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _12891_ (.A(message[120]),
    .B(_08305_),
    .Y(_08315_));
 sky130_fd_sc_hd__o21ai_0 _12892_ (.A1(_07974_),
    .A2(_08305_),
    .B1(_08315_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _12893_ (.A(message[119]),
    .B(_08305_),
    .Y(_08316_));
 sky130_fd_sc_hd__o21ai_0 _12894_ (.A1(_07981_),
    .A2(_08305_),
    .B1(_08316_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand2_1 _12896_ (.A(message[118]),
    .B(_08305_),
    .Y(_08318_));
 sky130_fd_sc_hd__o21ai_0 _12897_ (.A1(_07989_),
    .A2(_08305_),
    .B1(_08318_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _12899_ (.A(message[117]),
    .B(_08305_),
    .Y(_08320_));
 sky130_fd_sc_hd__o21ai_0 _12900_ (.A1(_08006_),
    .A2(_08305_),
    .B1(_08320_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _12901_ (.A(message[116]),
    .B(_08305_),
    .Y(_08321_));
 sky130_fd_sc_hd__o21ai_0 _12902_ (.A1(_08018_),
    .A2(_08305_),
    .B1(_08321_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _12903_ (.A(message[115]),
    .B(_08305_),
    .Y(_08322_));
 sky130_fd_sc_hd__o21ai_0 _12904_ (.A1(_08025_),
    .A2(_08305_),
    .B1(_08322_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _12905_ (.A(message[114]),
    .B(_08305_),
    .Y(_08323_));
 sky130_fd_sc_hd__o21ai_0 _12906_ (.A1(_08031_),
    .A2(_08305_),
    .B1(_08323_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _12907_ (.A(message[113]),
    .B(_08305_),
    .Y(_08324_));
 sky130_fd_sc_hd__o21ai_0 _12908_ (.A1(_08039_),
    .A2(_08305_),
    .B1(_08324_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _12909_ (.A(message[112]),
    .B(_08305_),
    .Y(_08325_));
 sky130_fd_sc_hd__o21ai_0 _12910_ (.A1(_08051_),
    .A2(_08305_),
    .B1(_08325_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _12911_ (.A(message[111]),
    .B(_08305_),
    .Y(_08326_));
 sky130_fd_sc_hd__o21ai_0 _12912_ (.A1(_08064_),
    .A2(_08305_),
    .B1(_08326_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _12913_ (.A(message[110]),
    .B(_08305_),
    .Y(_08327_));
 sky130_fd_sc_hd__o21ai_0 _12914_ (.A1(_08071_),
    .A2(_08305_),
    .B1(_08327_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _12915_ (.A(message[109]),
    .B(_08305_),
    .Y(_08328_));
 sky130_fd_sc_hd__o21ai_0 _12916_ (.A1(_08082_),
    .A2(_08305_),
    .B1(_08328_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _12918_ (.A(message[108]),
    .B(_08305_),
    .Y(_08330_));
 sky130_fd_sc_hd__o21ai_0 _12919_ (.A1(_08091_),
    .A2(_08305_),
    .B1(_08330_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _12921_ (.A(message[107]),
    .B(_08305_),
    .Y(_08332_));
 sky130_fd_sc_hd__o21ai_0 _12922_ (.A1(_08102_),
    .A2(_08305_),
    .B1(_08332_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _12923_ (.A(message[106]),
    .B(_08305_),
    .Y(_08333_));
 sky130_fd_sc_hd__o21ai_0 _12924_ (.A1(_08114_),
    .A2(_08305_),
    .B1(_08333_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _12925_ (.A(message[105]),
    .B(_08305_),
    .Y(_08334_));
 sky130_fd_sc_hd__o21ai_0 _12926_ (.A1(_08125_),
    .A2(_08305_),
    .B1(_08334_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _12927_ (.A(message[104]),
    .B(_08305_),
    .Y(_08335_));
 sky130_fd_sc_hd__o21ai_0 _12928_ (.A1(_08142_),
    .A2(_08305_),
    .B1(_08335_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _12929_ (.A(message[103]),
    .B(_08305_),
    .Y(_08336_));
 sky130_fd_sc_hd__o21ai_1 _12930_ (.A1(_08152_),
    .A2(_08305_),
    .B1(_08336_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _12931_ (.A(message[102]),
    .B(_08305_),
    .Y(_08337_));
 sky130_fd_sc_hd__o21ai_0 _12932_ (.A1(_08160_),
    .A2(_08305_),
    .B1(_08337_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _12933_ (.A(message[101]),
    .B(_08305_),
    .Y(_08338_));
 sky130_fd_sc_hd__o21ai_0 _12934_ (.A1(_08171_),
    .A2(_08305_),
    .B1(_08338_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _12935_ (.A(message[100]),
    .B(_08305_),
    .Y(_08339_));
 sky130_fd_sc_hd__o21ai_0 _12936_ (.A1(_08184_),
    .A2(_08305_),
    .B1(_08339_),
    .Y(_00436_));
 sky130_fd_sc_hd__a21oi_1 _12939_ (.A1(_05403_),
    .A2(_08304_),
    .B1(message[99]),
    .Y(_08342_));
 sky130_fd_sc_hd__a31oi_1 _12940_ (.A1(_05403_),
    .A2(_08204_),
    .A3(_08304_),
    .B1(_08342_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _12941_ (.A(message[98]),
    .B(_08305_),
    .Y(_08343_));
 sky130_fd_sc_hd__o21ai_0 _12942_ (.A1(_08209_),
    .A2(_08305_),
    .B1(_08343_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(message[97]),
    .B(_08305_),
    .Y(_08344_));
 sky130_fd_sc_hd__o21ai_0 _12944_ (.A1(_08221_),
    .A2(_08305_),
    .B1(_08344_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _12945_ (.A(message[96]),
    .B(_08305_),
    .Y(_08345_));
 sky130_fd_sc_hd__o21ai_1 _12946_ (.A1(_08254_),
    .A2(_08305_),
    .B1(_08345_),
    .Y(_00441_));
 sky130_fd_sc_hd__nor2b_1 _12947_ (.A(reset),
    .B_N(_09555_),
    .Y(_08346_));
 sky130_fd_sc_hd__nand2_1 _12949_ (.A(_05338_),
    .B(_08346_),
    .Y(_08348_));
 sky130_fd_sc_hd__nand2_1 _12952_ (.A(message[159]),
    .B(_08348_),
    .Y(_08351_));
 sky130_fd_sc_hd__o21ai_0 _12953_ (.A1(_07572_),
    .A2(_08348_),
    .B1(_08351_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _12954_ (.A(message[158]),
    .B(_08348_),
    .Y(_08352_));
 sky130_fd_sc_hd__o21ai_0 _12955_ (.A1(_07577_),
    .A2(_08348_),
    .B1(_08352_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _12958_ (.A(message[157]),
    .B(_08348_),
    .Y(_08355_));
 sky130_fd_sc_hd__o21ai_0 _12959_ (.A1(_07581_),
    .A2(_08348_),
    .B1(_08355_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _12960_ (.A(message[156]),
    .B(_08348_),
    .Y(_08356_));
 sky130_fd_sc_hd__o21ai_0 _12961_ (.A1(_07588_),
    .A2(_08348_),
    .B1(_08356_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _12962_ (.A(message[155]),
    .B(_08348_),
    .Y(_08357_));
 sky130_fd_sc_hd__o21ai_0 _12963_ (.A1(_07601_),
    .A2(_08348_),
    .B1(_08357_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _12964_ (.A(message[154]),
    .B(_08348_),
    .Y(_08358_));
 sky130_fd_sc_hd__o21ai_0 _12965_ (.A1(_07610_),
    .A2(_08348_),
    .B1(_08358_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _12966_ (.A(message[153]),
    .B(_08348_),
    .Y(_08359_));
 sky130_fd_sc_hd__o21ai_0 _12967_ (.A1(_07620_),
    .A2(_08348_),
    .B1(_08359_),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _12968_ (.A(message[152]),
    .B(_08348_),
    .Y(_08360_));
 sky130_fd_sc_hd__o21ai_0 _12969_ (.A1(_07628_),
    .A2(_08348_),
    .B1(_08360_),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _12970_ (.A(message[151]),
    .B(_08348_),
    .Y(_08361_));
 sky130_fd_sc_hd__o21ai_0 _12971_ (.A1(_07635_),
    .A2(_08348_),
    .B1(_08361_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _12972_ (.A(message[150]),
    .B(_08348_),
    .Y(_08362_));
 sky130_fd_sc_hd__o21ai_0 _12973_ (.A1(_07646_),
    .A2(_08348_),
    .B1(_08362_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_1 _12975_ (.A(message[149]),
    .B(_08348_),
    .Y(_08364_));
 sky130_fd_sc_hd__o21ai_0 _12976_ (.A1(_07660_),
    .A2(_08348_),
    .B1(_08364_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _12977_ (.A(message[148]),
    .B(_08348_),
    .Y(_08365_));
 sky130_fd_sc_hd__o21ai_0 _12978_ (.A1(_07669_),
    .A2(_08348_),
    .B1(_08365_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _12980_ (.A(message[147]),
    .B(_08348_),
    .Y(_08367_));
 sky130_fd_sc_hd__o21ai_0 _12981_ (.A1(_07677_),
    .A2(_08348_),
    .B1(_08367_),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _12982_ (.A(message[146]),
    .B(_08348_),
    .Y(_08368_));
 sky130_fd_sc_hd__o21ai_0 _12983_ (.A1(_07689_),
    .A2(_08348_),
    .B1(_08368_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _12984_ (.A(message[145]),
    .B(_08348_),
    .Y(_08369_));
 sky130_fd_sc_hd__o21ai_0 _12985_ (.A1(_07703_),
    .A2(_08348_),
    .B1(_08369_),
    .Y(_00454_));
 sky130_fd_sc_hd__nand2_1 _12986_ (.A(message[144]),
    .B(_08348_),
    .Y(_08370_));
 sky130_fd_sc_hd__o21ai_0 _12987_ (.A1(_07709_),
    .A2(_08348_),
    .B1(_08370_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _12988_ (.A(message[143]),
    .B(_08348_),
    .Y(_08371_));
 sky130_fd_sc_hd__o21ai_0 _12989_ (.A1(_07715_),
    .A2(_08348_),
    .B1(_08371_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _12990_ (.A(message[142]),
    .B(_08348_),
    .Y(_08372_));
 sky130_fd_sc_hd__o21ai_0 _12991_ (.A1(_07731_),
    .A2(_08348_),
    .B1(_08372_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _12992_ (.A(message[141]),
    .B(_08348_),
    .Y(_08373_));
 sky130_fd_sc_hd__o21ai_0 _12993_ (.A1(_07745_),
    .A2(_08348_),
    .B1(_08373_),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _12994_ (.A(message[140]),
    .B(_08348_),
    .Y(_08374_));
 sky130_fd_sc_hd__o21ai_0 _12995_ (.A1(_07752_),
    .A2(_08348_),
    .B1(_08374_),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _12996_ (.A(message[139]),
    .B(_08348_),
    .Y(_08375_));
 sky130_fd_sc_hd__o21ai_0 _12997_ (.A1(_07766_),
    .A2(_08348_),
    .B1(_08375_),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _12998_ (.A(message[138]),
    .B(_08348_),
    .Y(_08376_));
 sky130_fd_sc_hd__o21ai_0 _12999_ (.A1(_07777_),
    .A2(_08348_),
    .B1(_08376_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _13000_ (.A(message[137]),
    .B(_08348_),
    .Y(_08377_));
 sky130_fd_sc_hd__o21ai_0 _13001_ (.A1(_07786_),
    .A2(_08348_),
    .B1(_08377_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _13002_ (.A(message[136]),
    .B(_08348_),
    .Y(_08378_));
 sky130_fd_sc_hd__o21ai_0 _13003_ (.A1(_07800_),
    .A2(_08348_),
    .B1(_08378_),
    .Y(_00464_));
 sky130_fd_sc_hd__and2_1 _13004_ (.A(_05338_),
    .B(_08346_),
    .X(_08379_));
 sky130_fd_sc_hd__nor2_1 _13006_ (.A(message[135]),
    .B(_08379_),
    .Y(_08381_));
 sky130_fd_sc_hd__a21oi_1 _13007_ (.A1(_07809_),
    .A2(_08379_),
    .B1(_08381_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _13008_ (.A(message[134]),
    .B(_08348_),
    .Y(_08382_));
 sky130_fd_sc_hd__o21ai_0 _13009_ (.A1(_07818_),
    .A2(_08348_),
    .B1(_08382_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(message[133]),
    .B(_08348_),
    .Y(_08383_));
 sky130_fd_sc_hd__o21ai_0 _13011_ (.A1(_07831_),
    .A2(_08348_),
    .B1(_08383_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _13012_ (.A(message[132]),
    .B(_08348_),
    .Y(_08384_));
 sky130_fd_sc_hd__o21ai_0 _13013_ (.A1(_07843_),
    .A2(_08348_),
    .B1(_08384_),
    .Y(_00468_));
 sky130_fd_sc_hd__nor2_1 _13014_ (.A(message[131]),
    .B(_08379_),
    .Y(_08385_));
 sky130_fd_sc_hd__a21oi_1 _13015_ (.A1(_07850_),
    .A2(_08379_),
    .B1(_08385_),
    .Y(_00469_));
 sky130_fd_sc_hd__nor2_1 _13016_ (.A(_07860_),
    .B(_08348_),
    .Y(_08386_));
 sky130_fd_sc_hd__a21oi_1 _13017_ (.A1(message[130]),
    .A2(_08348_),
    .B1(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__a21oi_1 _13018_ (.A1(_07859_),
    .A2(_08379_),
    .B1(_08387_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _13019_ (.A(message[129]),
    .B(_08348_),
    .Y(_08388_));
 sky130_fd_sc_hd__o21ai_0 _13020_ (.A1(_07873_),
    .A2(_08348_),
    .B1(_08388_),
    .Y(_00472_));
 sky130_fd_sc_hd__nor2_1 _13021_ (.A(message[128]),
    .B(_08379_),
    .Y(_08389_));
 sky130_fd_sc_hd__a21oi_1 _13022_ (.A1(_07925_),
    .A2(_08379_),
    .B1(_08389_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2b_1 _13023_ (.A(reset),
    .B_N(_09563_),
    .Y(_08390_));
 sky130_fd_sc_hd__nand2_1 _13024_ (.A(_05403_),
    .B(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__nand2_1 _13027_ (.A(message[191]),
    .B(_08391_),
    .Y(_08394_));
 sky130_fd_sc_hd__o21ai_0 _13028_ (.A1(_07930_),
    .A2(_08391_),
    .B1(_08394_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _13029_ (.A(message[190]),
    .B(_08391_),
    .Y(_08395_));
 sky130_fd_sc_hd__o21ai_0 _13030_ (.A1(_07934_),
    .A2(_08391_),
    .B1(_08395_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _13031_ (.A(message[189]),
    .B(_08391_),
    .Y(_08396_));
 sky130_fd_sc_hd__o21ai_0 _13032_ (.A1(_07937_),
    .A2(_08391_),
    .B1(_08396_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _13033_ (.A(message[188]),
    .B(_08391_),
    .Y(_08397_));
 sky130_fd_sc_hd__o21ai_0 _13034_ (.A1(_07942_),
    .A2(_08391_),
    .B1(_08397_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _13035_ (.A(message[187]),
    .B(_08391_),
    .Y(_08398_));
 sky130_fd_sc_hd__o21ai_0 _13036_ (.A1(_07949_),
    .A2(_08391_),
    .B1(_08398_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _13037_ (.A(message[186]),
    .B(_08391_),
    .Y(_08399_));
 sky130_fd_sc_hd__o21ai_0 _13038_ (.A1(_07956_),
    .A2(_08391_),
    .B1(_08399_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _13039_ (.A(message[185]),
    .B(_08391_),
    .Y(_08400_));
 sky130_fd_sc_hd__o21ai_0 _13040_ (.A1(_07965_),
    .A2(_08391_),
    .B1(_08400_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _13041_ (.A(message[184]),
    .B(_08391_),
    .Y(_08401_));
 sky130_fd_sc_hd__o21ai_0 _13042_ (.A1(_07974_),
    .A2(_08391_),
    .B1(_08401_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _13043_ (.A(message[183]),
    .B(_08391_),
    .Y(_08402_));
 sky130_fd_sc_hd__o21ai_0 _13044_ (.A1(_07981_),
    .A2(_08391_),
    .B1(_08402_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _13046_ (.A(message[182]),
    .B(_08391_),
    .Y(_08404_));
 sky130_fd_sc_hd__o21ai_0 _13047_ (.A1(_07989_),
    .A2(_08391_),
    .B1(_08404_),
    .Y(_00512_));
 sky130_fd_sc_hd__nand2_1 _13049_ (.A(message[181]),
    .B(_08391_),
    .Y(_08406_));
 sky130_fd_sc_hd__o21ai_0 _13050_ (.A1(_08006_),
    .A2(_08391_),
    .B1(_08406_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _13051_ (.A(message[180]),
    .B(_08391_),
    .Y(_08407_));
 sky130_fd_sc_hd__o21ai_0 _13052_ (.A1(_08018_),
    .A2(_08391_),
    .B1(_08407_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _13053_ (.A(message[179]),
    .B(_08391_),
    .Y(_08408_));
 sky130_fd_sc_hd__o21ai_0 _13054_ (.A1(_08025_),
    .A2(_08391_),
    .B1(_08408_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _13055_ (.A(message[178]),
    .B(_08391_),
    .Y(_08409_));
 sky130_fd_sc_hd__o21ai_0 _13056_ (.A1(_08031_),
    .A2(_08391_),
    .B1(_08409_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _13057_ (.A(message[177]),
    .B(_08391_),
    .Y(_08410_));
 sky130_fd_sc_hd__o21ai_0 _13058_ (.A1(_08039_),
    .A2(_08391_),
    .B1(_08410_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _13059_ (.A(message[176]),
    .B(_08391_),
    .Y(_08411_));
 sky130_fd_sc_hd__o21ai_0 _13060_ (.A1(_08051_),
    .A2(_08391_),
    .B1(_08411_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _13061_ (.A(message[175]),
    .B(_08391_),
    .Y(_08412_));
 sky130_fd_sc_hd__o21ai_0 _13062_ (.A1(_08064_),
    .A2(_08391_),
    .B1(_08412_),
    .Y(_00488_));
 sky130_fd_sc_hd__nand2_1 _13063_ (.A(message[174]),
    .B(_08391_),
    .Y(_08413_));
 sky130_fd_sc_hd__o21ai_0 _13064_ (.A1(_08071_),
    .A2(_08391_),
    .B1(_08413_),
    .Y(_00489_));
 sky130_fd_sc_hd__nand2_1 _13065_ (.A(message[173]),
    .B(_08391_),
    .Y(_08414_));
 sky130_fd_sc_hd__o21ai_0 _13066_ (.A1(_08082_),
    .A2(_08391_),
    .B1(_08414_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_1 _13068_ (.A(message[172]),
    .B(_08391_),
    .Y(_08416_));
 sky130_fd_sc_hd__o21ai_0 _13069_ (.A1(_08091_),
    .A2(_08391_),
    .B1(_08416_),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _13071_ (.A(message[171]),
    .B(_08391_),
    .Y(_08418_));
 sky130_fd_sc_hd__o21ai_0 _13072_ (.A1(_08102_),
    .A2(_08391_),
    .B1(_08418_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _13073_ (.A(message[170]),
    .B(_08391_),
    .Y(_08419_));
 sky130_fd_sc_hd__o21ai_0 _13074_ (.A1(_08114_),
    .A2(_08391_),
    .B1(_08419_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _13075_ (.A(message[169]),
    .B(_08391_),
    .Y(_08420_));
 sky130_fd_sc_hd__o21ai_0 _13076_ (.A1(_08125_),
    .A2(_08391_),
    .B1(_08420_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand2_1 _13077_ (.A(message[168]),
    .B(_08391_),
    .Y(_08421_));
 sky130_fd_sc_hd__o21ai_0 _13078_ (.A1(_08142_),
    .A2(_08391_),
    .B1(_08421_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _13079_ (.A(message[167]),
    .B(_08391_),
    .Y(_08422_));
 sky130_fd_sc_hd__o21ai_0 _13080_ (.A1(_08152_),
    .A2(_08391_),
    .B1(_08422_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _13081_ (.A(message[166]),
    .B(_08391_),
    .Y(_08423_));
 sky130_fd_sc_hd__o21ai_0 _13082_ (.A1(_08160_),
    .A2(_08391_),
    .B1(_08423_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _13083_ (.A(message[165]),
    .B(_08391_),
    .Y(_08424_));
 sky130_fd_sc_hd__o21ai_0 _13084_ (.A1(_08171_),
    .A2(_08391_),
    .B1(_08424_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _13085_ (.A(message[164]),
    .B(_08391_),
    .Y(_08425_));
 sky130_fd_sc_hd__o21ai_0 _13086_ (.A1(_08184_),
    .A2(_08391_),
    .B1(_08425_),
    .Y(_00500_));
 sky130_fd_sc_hd__a21oi_1 _13088_ (.A1(_05403_),
    .A2(_08390_),
    .B1(message[163]),
    .Y(_08427_));
 sky130_fd_sc_hd__a31oi_1 _13089_ (.A1(_05403_),
    .A2(_08204_),
    .A3(_08390_),
    .B1(_08427_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _13090_ (.A(message[162]),
    .B(_08391_),
    .Y(_08428_));
 sky130_fd_sc_hd__o21ai_0 _13091_ (.A1(_08209_),
    .A2(_08391_),
    .B1(_08428_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2_1 _13092_ (.A(message[161]),
    .B(_08391_),
    .Y(_08429_));
 sky130_fd_sc_hd__o21ai_0 _13093_ (.A1(_08221_),
    .A2(_08391_),
    .B1(_08429_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _13094_ (.A(message[160]),
    .B(_08391_),
    .Y(_08430_));
 sky130_fd_sc_hd__o21ai_1 _13095_ (.A1(_08254_),
    .A2(_08391_),
    .B1(_08430_),
    .Y(_00505_));
 sky130_fd_sc_hd__nor2b_1 _13096_ (.A(reset),
    .B_N(_09559_),
    .Y(_08431_));
 sky130_fd_sc_hd__nand2_1 _13098_ (.A(_05338_),
    .B(_08431_),
    .Y(_08433_));
 sky130_fd_sc_hd__nand2_1 _13101_ (.A(message[223]),
    .B(_08433_),
    .Y(_08436_));
 sky130_fd_sc_hd__o21ai_0 _13102_ (.A1(_07572_),
    .A2(_08433_),
    .B1(_08436_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _13103_ (.A(message[222]),
    .B(_08433_),
    .Y(_08437_));
 sky130_fd_sc_hd__o21ai_0 _13104_ (.A1(_07577_),
    .A2(_08433_),
    .B1(_08437_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _13107_ (.A(message[221]),
    .B(_08433_),
    .Y(_08440_));
 sky130_fd_sc_hd__o21ai_0 _13108_ (.A1(_07581_),
    .A2(_08433_),
    .B1(_08440_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _13109_ (.A(message[220]),
    .B(_08433_),
    .Y(_08441_));
 sky130_fd_sc_hd__o21ai_0 _13110_ (.A1(_07588_),
    .A2(_08433_),
    .B1(_08441_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _13111_ (.A(message[219]),
    .B(_08433_),
    .Y(_08442_));
 sky130_fd_sc_hd__o21ai_0 _13112_ (.A1(_07601_),
    .A2(_08433_),
    .B1(_08442_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand2_1 _13113_ (.A(message[218]),
    .B(_08433_),
    .Y(_08443_));
 sky130_fd_sc_hd__o21ai_0 _13114_ (.A1(_07610_),
    .A2(_08433_),
    .B1(_08443_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _13115_ (.A(message[217]),
    .B(_08433_),
    .Y(_08444_));
 sky130_fd_sc_hd__o21ai_0 _13116_ (.A1(_07620_),
    .A2(_08433_),
    .B1(_08444_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _13117_ (.A(message[216]),
    .B(_08433_),
    .Y(_08445_));
 sky130_fd_sc_hd__o21ai_0 _13118_ (.A1(_07628_),
    .A2(_08433_),
    .B1(_08445_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _13119_ (.A(message[215]),
    .B(_08433_),
    .Y(_08446_));
 sky130_fd_sc_hd__o21ai_0 _13120_ (.A1(_07635_),
    .A2(_08433_),
    .B1(_08446_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _13121_ (.A(message[214]),
    .B(_08433_),
    .Y(_08447_));
 sky130_fd_sc_hd__o21ai_0 _13122_ (.A1(_07646_),
    .A2(_08433_),
    .B1(_08447_),
    .Y(_00544_));
 sky130_fd_sc_hd__nand2_1 _13124_ (.A(message[213]),
    .B(_08433_),
    .Y(_08449_));
 sky130_fd_sc_hd__o21ai_0 _13125_ (.A1(_07660_),
    .A2(_08433_),
    .B1(_08449_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _13126_ (.A(message[212]),
    .B(_08433_),
    .Y(_08450_));
 sky130_fd_sc_hd__o21ai_0 _13127_ (.A1(_07669_),
    .A2(_08433_),
    .B1(_08450_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _13129_ (.A(message[211]),
    .B(_08433_),
    .Y(_08452_));
 sky130_fd_sc_hd__o21ai_0 _13130_ (.A1(_07677_),
    .A2(_08433_),
    .B1(_08452_),
    .Y(_00516_));
 sky130_fd_sc_hd__nand2_1 _13131_ (.A(message[210]),
    .B(_08433_),
    .Y(_08453_));
 sky130_fd_sc_hd__o21ai_0 _13132_ (.A1(_07689_),
    .A2(_08433_),
    .B1(_08453_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _13133_ (.A(message[209]),
    .B(_08433_),
    .Y(_08454_));
 sky130_fd_sc_hd__o21ai_0 _13134_ (.A1(_07703_),
    .A2(_08433_),
    .B1(_08454_),
    .Y(_00518_));
 sky130_fd_sc_hd__nand2_1 _13135_ (.A(message[208]),
    .B(_08433_),
    .Y(_08455_));
 sky130_fd_sc_hd__o21ai_0 _13136_ (.A1(_07709_),
    .A2(_08433_),
    .B1(_08455_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _13137_ (.A(message[207]),
    .B(_08433_),
    .Y(_08456_));
 sky130_fd_sc_hd__o21ai_0 _13138_ (.A1(_07715_),
    .A2(_08433_),
    .B1(_08456_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _13139_ (.A(message[206]),
    .B(_08433_),
    .Y(_08457_));
 sky130_fd_sc_hd__o21ai_0 _13140_ (.A1(_07731_),
    .A2(_08433_),
    .B1(_08457_),
    .Y(_00521_));
 sky130_fd_sc_hd__nand2_1 _13141_ (.A(message[205]),
    .B(_08433_),
    .Y(_08458_));
 sky130_fd_sc_hd__o21ai_0 _13142_ (.A1(_07745_),
    .A2(_08433_),
    .B1(_08458_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_1 _13143_ (.A(message[204]),
    .B(_08433_),
    .Y(_08459_));
 sky130_fd_sc_hd__o21ai_0 _13144_ (.A1(_07752_),
    .A2(_08433_),
    .B1(_08459_),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2_1 _13145_ (.A(message[203]),
    .B(_08433_),
    .Y(_08460_));
 sky130_fd_sc_hd__o21ai_0 _13146_ (.A1(_07766_),
    .A2(_08433_),
    .B1(_08460_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _13147_ (.A(message[202]),
    .B(_08433_),
    .Y(_08461_));
 sky130_fd_sc_hd__o21ai_0 _13148_ (.A1(_07777_),
    .A2(_08433_),
    .B1(_08461_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _13149_ (.A(message[201]),
    .B(_08433_),
    .Y(_08462_));
 sky130_fd_sc_hd__o21ai_0 _13150_ (.A1(_07786_),
    .A2(_08433_),
    .B1(_08462_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _13151_ (.A(message[200]),
    .B(_08433_),
    .Y(_08463_));
 sky130_fd_sc_hd__o21ai_0 _13152_ (.A1(_07800_),
    .A2(_08433_),
    .B1(_08463_),
    .Y(_00528_));
 sky130_fd_sc_hd__and2_1 _13153_ (.A(_05338_),
    .B(_08431_),
    .X(_08464_));
 sky130_fd_sc_hd__nor2_1 _13155_ (.A(message[199]),
    .B(_08464_),
    .Y(_08466_));
 sky130_fd_sc_hd__a21oi_1 _13156_ (.A1(_07809_),
    .A2(_08464_),
    .B1(_08466_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _13157_ (.A(message[198]),
    .B(_08433_),
    .Y(_08467_));
 sky130_fd_sc_hd__o21ai_0 _13158_ (.A1(_07818_),
    .A2(_08433_),
    .B1(_08467_),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _13159_ (.A(message[197]),
    .B(_08433_),
    .Y(_08468_));
 sky130_fd_sc_hd__o21ai_0 _13160_ (.A1(_07831_),
    .A2(_08433_),
    .B1(_08468_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _13161_ (.A(message[196]),
    .B(_08433_),
    .Y(_08469_));
 sky130_fd_sc_hd__o21ai_0 _13162_ (.A1(_07843_),
    .A2(_08433_),
    .B1(_08469_),
    .Y(_00532_));
 sky130_fd_sc_hd__nor2_1 _13163_ (.A(message[195]),
    .B(_08464_),
    .Y(_08470_));
 sky130_fd_sc_hd__a21oi_1 _13164_ (.A1(_07850_),
    .A2(_08464_),
    .B1(_08470_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_1 _13165_ (.A(_07860_),
    .B(_08433_),
    .Y(_08471_));
 sky130_fd_sc_hd__a21oi_1 _13166_ (.A1(message[194]),
    .A2(_08433_),
    .B1(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__a21oi_1 _13167_ (.A1(_07859_),
    .A2(_08464_),
    .B1(_08472_),
    .Y(_00534_));
 sky130_fd_sc_hd__nand2_1 _13168_ (.A(message[193]),
    .B(_08433_),
    .Y(_08473_));
 sky130_fd_sc_hd__o21ai_0 _13169_ (.A1(_07873_),
    .A2(_08433_),
    .B1(_08473_),
    .Y(_00536_));
 sky130_fd_sc_hd__nor2_1 _13170_ (.A(message[192]),
    .B(_08464_),
    .Y(_08474_));
 sky130_fd_sc_hd__a21oi_1 _13171_ (.A1(_07925_),
    .A2(_08464_),
    .B1(_08474_),
    .Y(_00537_));
 sky130_fd_sc_hd__nor2b_1 _13172_ (.A(\count_2[5] ),
    .B_N(_09567_),
    .Y(_08475_));
 sky130_fd_sc_hd__nor3_1 _13173_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(reset),
    .Y(_08476_));
 sky130_fd_sc_hd__nand2_1 _13174_ (.A(_08475_),
    .B(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__nand2_1 _13178_ (.A(message[255]),
    .B(_08477_),
    .Y(_08481_));
 sky130_fd_sc_hd__o21ai_0 _13179_ (.A1(_07930_),
    .A2(_08477_),
    .B1(_08481_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _13180_ (.A(message[254]),
    .B(_08477_),
    .Y(_08482_));
 sky130_fd_sc_hd__o21ai_0 _13181_ (.A1(_07934_),
    .A2(_08477_),
    .B1(_08482_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand2_1 _13183_ (.A(message[253]),
    .B(_08477_),
    .Y(_08484_));
 sky130_fd_sc_hd__o21ai_0 _13184_ (.A1(_07937_),
    .A2(_08477_),
    .B1(_08484_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand2_1 _13185_ (.A(message[252]),
    .B(_08477_),
    .Y(_08485_));
 sky130_fd_sc_hd__o21ai_0 _13186_ (.A1(_07942_),
    .A2(_08477_),
    .B1(_08485_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _13187_ (.A(message[251]),
    .B(_08477_),
    .Y(_08486_));
 sky130_fd_sc_hd__o21ai_0 _13188_ (.A1(_07949_),
    .A2(_08477_),
    .B1(_08486_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _13189_ (.A(message[250]),
    .B(_08477_),
    .Y(_08487_));
 sky130_fd_sc_hd__o21ai_0 _13190_ (.A1(_07956_),
    .A2(_08477_),
    .B1(_08487_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _13191_ (.A(message[249]),
    .B(_08477_),
    .Y(_08488_));
 sky130_fd_sc_hd__o21ai_0 _13192_ (.A1(_07965_),
    .A2(_08477_),
    .B1(_08488_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _13193_ (.A(message[248]),
    .B(_08477_),
    .Y(_08489_));
 sky130_fd_sc_hd__o21ai_0 _13194_ (.A1(_07974_),
    .A2(_08477_),
    .B1(_08489_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _13195_ (.A(message[247]),
    .B(_08477_),
    .Y(_08490_));
 sky130_fd_sc_hd__o21ai_0 _13196_ (.A1(_07981_),
    .A2(_08477_),
    .B1(_08490_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _13197_ (.A(message[246]),
    .B(_08477_),
    .Y(_08491_));
 sky130_fd_sc_hd__o21ai_0 _13198_ (.A1(_07989_),
    .A2(_08477_),
    .B1(_08491_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _13200_ (.A(message[245]),
    .B(_08477_),
    .Y(_08493_));
 sky130_fd_sc_hd__o21ai_0 _13201_ (.A1(_08006_),
    .A2(_08477_),
    .B1(_08493_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _13202_ (.A(message[244]),
    .B(_08477_),
    .Y(_08494_));
 sky130_fd_sc_hd__o21ai_0 _13203_ (.A1(_08018_),
    .A2(_08477_),
    .B1(_08494_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _13205_ (.A(message[243]),
    .B(_08477_),
    .Y(_08496_));
 sky130_fd_sc_hd__o21ai_0 _13206_ (.A1(_08025_),
    .A2(_08477_),
    .B1(_08496_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _13207_ (.A(message[242]),
    .B(_08477_),
    .Y(_08497_));
 sky130_fd_sc_hd__o21ai_0 _13208_ (.A1(_08031_),
    .A2(_08477_),
    .B1(_08497_),
    .Y(_00549_));
 sky130_fd_sc_hd__and2_1 _13209_ (.A(_08475_),
    .B(_08476_),
    .X(_08498_));
 sky130_fd_sc_hd__nor2_1 _13211_ (.A(message[241]),
    .B(_08498_),
    .Y(_08500_));
 sky130_fd_sc_hd__a21oi_1 _13212_ (.A1(_08039_),
    .A2(_08498_),
    .B1(_08500_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _13213_ (.A(message[240]),
    .B(_08477_),
    .Y(_08501_));
 sky130_fd_sc_hd__o21ai_0 _13214_ (.A1(_08051_),
    .A2(_08477_),
    .B1(_08501_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _13215_ (.A(message[239]),
    .B(_08477_),
    .Y(_08502_));
 sky130_fd_sc_hd__o21ai_0 _13216_ (.A1(_08064_),
    .A2(_08477_),
    .B1(_08502_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _13217_ (.A(message[238]),
    .B(_08477_),
    .Y(_08503_));
 sky130_fd_sc_hd__o21ai_0 _13218_ (.A1(_08071_),
    .A2(_08477_),
    .B1(_08503_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_1 _13219_ (.A(message[237]),
    .B(_08477_),
    .Y(_08504_));
 sky130_fd_sc_hd__o21ai_0 _13220_ (.A1(_08082_),
    .A2(_08477_),
    .B1(_08504_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _13221_ (.A(message[236]),
    .B(_08477_),
    .Y(_08505_));
 sky130_fd_sc_hd__o21ai_0 _13222_ (.A1(_08091_),
    .A2(_08477_),
    .B1(_08505_),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _13223_ (.A(message[235]),
    .B(_08477_),
    .Y(_08506_));
 sky130_fd_sc_hd__o21ai_0 _13224_ (.A1(_08102_),
    .A2(_08477_),
    .B1(_08506_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _13225_ (.A(message[234]),
    .B(_08477_),
    .Y(_08507_));
 sky130_fd_sc_hd__o21ai_0 _13226_ (.A1(_08114_),
    .A2(_08477_),
    .B1(_08507_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_1 _13227_ (.A(message[233]),
    .B(_08477_),
    .Y(_08508_));
 sky130_fd_sc_hd__o21ai_0 _13228_ (.A1(_08125_),
    .A2(_08477_),
    .B1(_08508_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _13229_ (.A(message[232]),
    .B(_08477_),
    .Y(_08509_));
 sky130_fd_sc_hd__o21ai_0 _13230_ (.A1(_08142_),
    .A2(_08477_),
    .B1(_08509_),
    .Y(_00560_));
 sky130_fd_sc_hd__nor2_1 _13231_ (.A(message[231]),
    .B(_08498_),
    .Y(_08510_));
 sky130_fd_sc_hd__a21oi_1 _13232_ (.A1(_08152_),
    .A2(_08498_),
    .B1(_08510_),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_1 _13233_ (.A(message[230]),
    .B(_08477_),
    .Y(_08511_));
 sky130_fd_sc_hd__o21ai_0 _13234_ (.A1(_08160_),
    .A2(_08477_),
    .B1(_08511_),
    .Y(_00562_));
 sky130_fd_sc_hd__nor2_1 _13235_ (.A(message[229]),
    .B(_08498_),
    .Y(_08512_));
 sky130_fd_sc_hd__a21oi_1 _13236_ (.A1(_08171_),
    .A2(_08498_),
    .B1(_08512_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _13237_ (.A(message[228]),
    .B(_08477_),
    .Y(_08513_));
 sky130_fd_sc_hd__o21ai_0 _13238_ (.A1(_08184_),
    .A2(_08477_),
    .B1(_08513_),
    .Y(_00564_));
 sky130_fd_sc_hd__nor2_1 _13239_ (.A(message[227]),
    .B(_08498_),
    .Y(_08514_));
 sky130_fd_sc_hd__a21oi_1 _13240_ (.A1(_08204_),
    .A2(_08498_),
    .B1(_08514_),
    .Y(_00565_));
 sky130_fd_sc_hd__nand2_1 _13241_ (.A(message[226]),
    .B(_08477_),
    .Y(_08515_));
 sky130_fd_sc_hd__o21ai_0 _13242_ (.A1(_08209_),
    .A2(_08477_),
    .B1(_08515_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _13243_ (.A(message[225]),
    .B(_08477_),
    .Y(_08516_));
 sky130_fd_sc_hd__o21ai_0 _13244_ (.A1(_08221_),
    .A2(_08477_),
    .B1(_08516_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _13245_ (.A(message[224]),
    .B(_08477_),
    .Y(_08517_));
 sky130_fd_sc_hd__o21ai_1 _13246_ (.A1(_08254_),
    .A2(_08477_),
    .B1(_08517_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _13247_ (.A(_05343_),
    .B(_07566_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand2_1 _13250_ (.A(message[287]),
    .B(_08518_),
    .Y(_08521_));
 sky130_fd_sc_hd__o21ai_0 _13251_ (.A1(_07572_),
    .A2(_08518_),
    .B1(_08521_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _13252_ (.A(message[286]),
    .B(_08518_),
    .Y(_08522_));
 sky130_fd_sc_hd__o21ai_0 _13253_ (.A1(_07577_),
    .A2(_08518_),
    .B1(_08522_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _13256_ (.A(message[285]),
    .B(_08518_),
    .Y(_08525_));
 sky130_fd_sc_hd__o21ai_0 _13257_ (.A1(_07581_),
    .A2(_08518_),
    .B1(_08525_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _13258_ (.A(message[284]),
    .B(_08518_),
    .Y(_08526_));
 sky130_fd_sc_hd__o21ai_0 _13259_ (.A1(_07588_),
    .A2(_08518_),
    .B1(_08526_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _13260_ (.A(message[283]),
    .B(_08518_),
    .Y(_08527_));
 sky130_fd_sc_hd__o21ai_0 _13261_ (.A1(_07601_),
    .A2(_08518_),
    .B1(_08527_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _13262_ (.A(message[282]),
    .B(_08518_),
    .Y(_08528_));
 sky130_fd_sc_hd__o21ai_0 _13263_ (.A1(_07610_),
    .A2(_08518_),
    .B1(_08528_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _13264_ (.A(message[281]),
    .B(_08518_),
    .Y(_08529_));
 sky130_fd_sc_hd__o21ai_0 _13265_ (.A1(_07620_),
    .A2(_08518_),
    .B1(_08529_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _13266_ (.A(message[280]),
    .B(_08518_),
    .Y(_08530_));
 sky130_fd_sc_hd__o21ai_0 _13267_ (.A1(_07628_),
    .A2(_08518_),
    .B1(_08530_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _13268_ (.A(message[279]),
    .B(_08518_),
    .Y(_08531_));
 sky130_fd_sc_hd__o21ai_0 _13269_ (.A1(_07635_),
    .A2(_08518_),
    .B1(_08531_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _13270_ (.A(message[278]),
    .B(_08518_),
    .Y(_08532_));
 sky130_fd_sc_hd__o21ai_0 _13271_ (.A1(_07646_),
    .A2(_08518_),
    .B1(_08532_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _13273_ (.A(message[277]),
    .B(_08518_),
    .Y(_08534_));
 sky130_fd_sc_hd__o21ai_0 _13274_ (.A1(_07660_),
    .A2(_08518_),
    .B1(_08534_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _13275_ (.A(message[276]),
    .B(_08518_),
    .Y(_08535_));
 sky130_fd_sc_hd__o21ai_0 _13276_ (.A1(_07669_),
    .A2(_08518_),
    .B1(_08535_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _13278_ (.A(message[275]),
    .B(_08518_),
    .Y(_08537_));
 sky130_fd_sc_hd__o21ai_0 _13279_ (.A1(_07677_),
    .A2(_08518_),
    .B1(_08537_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_1 _13280_ (.A(message[274]),
    .B(_08518_),
    .Y(_08538_));
 sky130_fd_sc_hd__o21ai_0 _13281_ (.A1(_07689_),
    .A2(_08518_),
    .B1(_08538_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_1 _13282_ (.A(message[273]),
    .B(_08518_),
    .Y(_08539_));
 sky130_fd_sc_hd__o21ai_0 _13283_ (.A1(_07703_),
    .A2(_08518_),
    .B1(_08539_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _13284_ (.A(message[272]),
    .B(_08518_),
    .Y(_08540_));
 sky130_fd_sc_hd__o21ai_0 _13285_ (.A1(_07709_),
    .A2(_08518_),
    .B1(_08540_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _13286_ (.A(message[271]),
    .B(_08518_),
    .Y(_08541_));
 sky130_fd_sc_hd__o21ai_0 _13287_ (.A1(_07715_),
    .A2(_08518_),
    .B1(_08541_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _13288_ (.A(message[270]),
    .B(_08518_),
    .Y(_08542_));
 sky130_fd_sc_hd__o21ai_0 _13289_ (.A1(_07731_),
    .A2(_08518_),
    .B1(_08542_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_1 _13290_ (.A(message[269]),
    .B(_08518_),
    .Y(_08543_));
 sky130_fd_sc_hd__o21ai_0 _13291_ (.A1(_07745_),
    .A2(_08518_),
    .B1(_08543_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _13292_ (.A(message[268]),
    .B(_08518_),
    .Y(_08544_));
 sky130_fd_sc_hd__o21ai_0 _13293_ (.A1(_07752_),
    .A2(_08518_),
    .B1(_08544_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_1 _13294_ (.A(message[267]),
    .B(_08518_),
    .Y(_08545_));
 sky130_fd_sc_hd__o21ai_0 _13295_ (.A1(_07766_),
    .A2(_08518_),
    .B1(_08545_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _13296_ (.A(message[266]),
    .B(_08518_),
    .Y(_08546_));
 sky130_fd_sc_hd__o21ai_0 _13297_ (.A1(_07777_),
    .A2(_08518_),
    .B1(_08546_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _13298_ (.A(message[265]),
    .B(_08518_),
    .Y(_08547_));
 sky130_fd_sc_hd__o21ai_0 _13299_ (.A1(_07786_),
    .A2(_08518_),
    .B1(_08547_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand2_1 _13300_ (.A(message[264]),
    .B(_08518_),
    .Y(_08548_));
 sky130_fd_sc_hd__o21ai_0 _13301_ (.A1(_07800_),
    .A2(_08518_),
    .B1(_08548_),
    .Y(_00592_));
 sky130_fd_sc_hd__and2_1 _13302_ (.A(_05343_),
    .B(_07566_),
    .X(_08549_));
 sky130_fd_sc_hd__nor2_1 _13304_ (.A(message[263]),
    .B(_08549_),
    .Y(_08551_));
 sky130_fd_sc_hd__a21oi_1 _13305_ (.A1(_07809_),
    .A2(_08549_),
    .B1(_08551_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _13306_ (.A(message[262]),
    .B(_08518_),
    .Y(_08552_));
 sky130_fd_sc_hd__o21ai_0 _13307_ (.A1(_07818_),
    .A2(_08518_),
    .B1(_08552_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _13308_ (.A(message[261]),
    .B(_08518_),
    .Y(_08553_));
 sky130_fd_sc_hd__o21ai_0 _13309_ (.A1(_07831_),
    .A2(_08518_),
    .B1(_08553_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _13310_ (.A(message[260]),
    .B(_08518_),
    .Y(_08554_));
 sky130_fd_sc_hd__o21ai_0 _13311_ (.A1(_07843_),
    .A2(_08518_),
    .B1(_08554_),
    .Y(_00596_));
 sky130_fd_sc_hd__nor2_1 _13312_ (.A(message[259]),
    .B(_08549_),
    .Y(_08555_));
 sky130_fd_sc_hd__a21oi_1 _13313_ (.A1(_07850_),
    .A2(_08549_),
    .B1(_08555_),
    .Y(_00597_));
 sky130_fd_sc_hd__nor2_1 _13314_ (.A(_07860_),
    .B(_08518_),
    .Y(_08556_));
 sky130_fd_sc_hd__a21oi_1 _13315_ (.A1(message[258]),
    .A2(_08518_),
    .B1(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__a21oi_1 _13316_ (.A1(_07859_),
    .A2(_08549_),
    .B1(_08557_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _13317_ (.A(message[257]),
    .B(_08518_),
    .Y(_08558_));
 sky130_fd_sc_hd__o21ai_0 _13318_ (.A1(_07873_),
    .A2(_08518_),
    .B1(_08558_),
    .Y(_00600_));
 sky130_fd_sc_hd__nor2_1 _13319_ (.A(message[256]),
    .B(_08549_),
    .Y(_08559_));
 sky130_fd_sc_hd__a21oi_1 _13320_ (.A1(_07925_),
    .A2(_08549_),
    .B1(_08559_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _13321_ (.A(_05389_),
    .B(_07927_),
    .Y(_08560_));
 sky130_fd_sc_hd__nand2_1 _13324_ (.A(message[319]),
    .B(_08560_),
    .Y(_08563_));
 sky130_fd_sc_hd__o21ai_0 _13325_ (.A1(_07930_),
    .A2(_08560_),
    .B1(_08563_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _13326_ (.A(message[318]),
    .B(_08560_),
    .Y(_08564_));
 sky130_fd_sc_hd__o21ai_0 _13327_ (.A1(_07934_),
    .A2(_08560_),
    .B1(_08564_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _13328_ (.A(message[317]),
    .B(_08560_),
    .Y(_08565_));
 sky130_fd_sc_hd__o21ai_0 _13329_ (.A1(_07937_),
    .A2(_08560_),
    .B1(_08565_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _13330_ (.A(message[316]),
    .B(_08560_),
    .Y(_08566_));
 sky130_fd_sc_hd__o21ai_0 _13331_ (.A1(_07942_),
    .A2(_08560_),
    .B1(_08566_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _13332_ (.A(message[315]),
    .B(_08560_),
    .Y(_08567_));
 sky130_fd_sc_hd__o21ai_0 _13333_ (.A1(_07949_),
    .A2(_08560_),
    .B1(_08567_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _13334_ (.A(message[314]),
    .B(_08560_),
    .Y(_08568_));
 sky130_fd_sc_hd__o21ai_0 _13335_ (.A1(_07956_),
    .A2(_08560_),
    .B1(_08568_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _13336_ (.A(message[313]),
    .B(_08560_),
    .Y(_08569_));
 sky130_fd_sc_hd__o21ai_0 _13337_ (.A1(_07965_),
    .A2(_08560_),
    .B1(_08569_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _13338_ (.A(message[312]),
    .B(_08560_),
    .Y(_08570_));
 sky130_fd_sc_hd__o21ai_0 _13339_ (.A1(_07974_),
    .A2(_08560_),
    .B1(_08570_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(message[311]),
    .B(_08560_),
    .Y(_08571_));
 sky130_fd_sc_hd__o21ai_0 _13341_ (.A1(_07981_),
    .A2(_08560_),
    .B1(_08571_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2_1 _13343_ (.A(message[310]),
    .B(_08560_),
    .Y(_08573_));
 sky130_fd_sc_hd__o21ai_0 _13344_ (.A1(_07989_),
    .A2(_08560_),
    .B1(_08573_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _13346_ (.A(message[309]),
    .B(_08560_),
    .Y(_08575_));
 sky130_fd_sc_hd__o21ai_0 _13347_ (.A1(_08006_),
    .A2(_08560_),
    .B1(_08575_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _13348_ (.A(message[308]),
    .B(_08560_),
    .Y(_08576_));
 sky130_fd_sc_hd__o21ai_0 _13349_ (.A1(_08018_),
    .A2(_08560_),
    .B1(_08576_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _13350_ (.A(message[307]),
    .B(_08560_),
    .Y(_08577_));
 sky130_fd_sc_hd__o21ai_0 _13351_ (.A1(_08025_),
    .A2(_08560_),
    .B1(_08577_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _13352_ (.A(message[306]),
    .B(_08560_),
    .Y(_08578_));
 sky130_fd_sc_hd__o21ai_0 _13353_ (.A1(_08031_),
    .A2(_08560_),
    .B1(_08578_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _13354_ (.A(message[305]),
    .B(_08560_),
    .Y(_08579_));
 sky130_fd_sc_hd__o21ai_0 _13355_ (.A1(_08039_),
    .A2(_08560_),
    .B1(_08579_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _13356_ (.A(message[304]),
    .B(_08560_),
    .Y(_08580_));
 sky130_fd_sc_hd__o21ai_0 _13357_ (.A1(_08051_),
    .A2(_08560_),
    .B1(_08580_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _13358_ (.A(message[303]),
    .B(_08560_),
    .Y(_08581_));
 sky130_fd_sc_hd__o21ai_0 _13359_ (.A1(_08064_),
    .A2(_08560_),
    .B1(_08581_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _13360_ (.A(message[302]),
    .B(_08560_),
    .Y(_08582_));
 sky130_fd_sc_hd__o21ai_0 _13361_ (.A1(_08071_),
    .A2(_08560_),
    .B1(_08582_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _13362_ (.A(message[301]),
    .B(_08560_),
    .Y(_08583_));
 sky130_fd_sc_hd__o21ai_0 _13363_ (.A1(_08082_),
    .A2(_08560_),
    .B1(_08583_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand2_1 _13365_ (.A(message[300]),
    .B(_08560_),
    .Y(_08585_));
 sky130_fd_sc_hd__o21ai_0 _13366_ (.A1(_08091_),
    .A2(_08560_),
    .B1(_08585_),
    .Y(_00619_));
 sky130_fd_sc_hd__nand2_1 _13368_ (.A(message[299]),
    .B(_08560_),
    .Y(_08587_));
 sky130_fd_sc_hd__o21ai_0 _13369_ (.A1(_08102_),
    .A2(_08560_),
    .B1(_08587_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _13370_ (.A(message[298]),
    .B(_08560_),
    .Y(_08588_));
 sky130_fd_sc_hd__o21ai_0 _13371_ (.A1(_08114_),
    .A2(_08560_),
    .B1(_08588_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _13372_ (.A(message[297]),
    .B(_08560_),
    .Y(_08589_));
 sky130_fd_sc_hd__o21ai_0 _13373_ (.A1(_08125_),
    .A2(_08560_),
    .B1(_08589_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _13374_ (.A(message[296]),
    .B(_08560_),
    .Y(_08590_));
 sky130_fd_sc_hd__o21ai_0 _13375_ (.A1(_08142_),
    .A2(_08560_),
    .B1(_08590_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _13376_ (.A(message[295]),
    .B(_08560_),
    .Y(_08591_));
 sky130_fd_sc_hd__o21ai_0 _13377_ (.A1(_08152_),
    .A2(_08560_),
    .B1(_08591_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _13378_ (.A(message[294]),
    .B(_08560_),
    .Y(_08592_));
 sky130_fd_sc_hd__o21ai_0 _13379_ (.A1(_08160_),
    .A2(_08560_),
    .B1(_08592_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _13380_ (.A(message[293]),
    .B(_08560_),
    .Y(_08593_));
 sky130_fd_sc_hd__o21ai_0 _13381_ (.A1(_08171_),
    .A2(_08560_),
    .B1(_08593_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _13382_ (.A(message[292]),
    .B(_08560_),
    .Y(_08594_));
 sky130_fd_sc_hd__o21ai_0 _13383_ (.A1(_08184_),
    .A2(_08560_),
    .B1(_08594_),
    .Y(_00628_));
 sky130_fd_sc_hd__a21oi_1 _13384_ (.A1(_05389_),
    .A2(_07927_),
    .B1(message[291]),
    .Y(_08595_));
 sky130_fd_sc_hd__a31oi_1 _13385_ (.A1(_05389_),
    .A2(_07927_),
    .A3(_08204_),
    .B1(_08595_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _13386_ (.A(message[290]),
    .B(_08560_),
    .Y(_08596_));
 sky130_fd_sc_hd__o21ai_0 _13387_ (.A1(_08209_),
    .A2(_08560_),
    .B1(_08596_),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _13388_ (.A(message[289]),
    .B(_08560_),
    .Y(_08597_));
 sky130_fd_sc_hd__o21ai_0 _13389_ (.A1(_08221_),
    .A2(_08560_),
    .B1(_08597_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _13390_ (.A(message[288]),
    .B(_08560_),
    .Y(_08598_));
 sky130_fd_sc_hd__o21ai_1 _13391_ (.A1(_08254_),
    .A2(_08560_),
    .B1(_08598_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _13392_ (.A(_05343_),
    .B(_08257_),
    .Y(_08599_));
 sky130_fd_sc_hd__nand2_1 _13396_ (.A(message[351]),
    .B(_08599_),
    .Y(_08603_));
 sky130_fd_sc_hd__o21ai_0 _13397_ (.A1(_07572_),
    .A2(_08599_),
    .B1(_08603_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _13398_ (.A(message[350]),
    .B(_08599_),
    .Y(_08604_));
 sky130_fd_sc_hd__o21ai_0 _13399_ (.A1(_07577_),
    .A2(_08599_),
    .B1(_08604_),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _13400_ (.A(message[349]),
    .B(_08599_),
    .Y(_08605_));
 sky130_fd_sc_hd__o21ai_0 _13401_ (.A1(_07581_),
    .A2(_08599_),
    .B1(_08605_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2_1 _13403_ (.A(message[348]),
    .B(_08599_),
    .Y(_08607_));
 sky130_fd_sc_hd__o21ai_0 _13404_ (.A1(_07588_),
    .A2(_08599_),
    .B1(_08607_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _13405_ (.A(message[347]),
    .B(_08599_),
    .Y(_08608_));
 sky130_fd_sc_hd__o21ai_0 _13406_ (.A1(_07601_),
    .A2(_08599_),
    .B1(_08608_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _13407_ (.A(message[346]),
    .B(_08599_),
    .Y(_08609_));
 sky130_fd_sc_hd__o21ai_0 _13408_ (.A1(_07610_),
    .A2(_08599_),
    .B1(_08609_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(message[345]),
    .B(_08599_),
    .Y(_08610_));
 sky130_fd_sc_hd__o21ai_0 _13410_ (.A1(_07620_),
    .A2(_08599_),
    .B1(_08610_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _13411_ (.A(message[344]),
    .B(_08599_),
    .Y(_08611_));
 sky130_fd_sc_hd__o21ai_0 _13412_ (.A1(_07628_),
    .A2(_08599_),
    .B1(_08611_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _13413_ (.A(message[343]),
    .B(_08599_),
    .Y(_08612_));
 sky130_fd_sc_hd__o21ai_0 _13414_ (.A1(_07635_),
    .A2(_08599_),
    .B1(_08612_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _13415_ (.A(message[342]),
    .B(_08599_),
    .Y(_08613_));
 sky130_fd_sc_hd__o21ai_0 _13416_ (.A1(_07646_),
    .A2(_08599_),
    .B1(_08613_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _13418_ (.A(message[341]),
    .B(_08599_),
    .Y(_08615_));
 sky130_fd_sc_hd__o21ai_0 _13419_ (.A1(_07660_),
    .A2(_08599_),
    .B1(_08615_),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _13420_ (.A(message[340]),
    .B(_08599_),
    .Y(_08616_));
 sky130_fd_sc_hd__o21ai_0 _13421_ (.A1(_07669_),
    .A2(_08599_),
    .B1(_08616_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(message[339]),
    .B(_08599_),
    .Y(_08617_));
 sky130_fd_sc_hd__o21ai_0 _13423_ (.A1(_07677_),
    .A2(_08599_),
    .B1(_08617_),
    .Y(_00164_));
 sky130_fd_sc_hd__nand2_1 _13425_ (.A(message[338]),
    .B(_08599_),
    .Y(_08619_));
 sky130_fd_sc_hd__o21ai_0 _13426_ (.A1(_07689_),
    .A2(_08599_),
    .B1(_08619_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _13427_ (.A(message[337]),
    .B(_08599_),
    .Y(_08620_));
 sky130_fd_sc_hd__o21ai_0 _13428_ (.A1(_07703_),
    .A2(_08599_),
    .B1(_08620_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand2_1 _13429_ (.A(message[336]),
    .B(_08599_),
    .Y(_08621_));
 sky130_fd_sc_hd__o21ai_0 _13430_ (.A1(_07709_),
    .A2(_08599_),
    .B1(_08621_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _13431_ (.A(message[335]),
    .B(_08599_),
    .Y(_08622_));
 sky130_fd_sc_hd__o21ai_0 _13432_ (.A1(_07715_),
    .A2(_08599_),
    .B1(_08622_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _13433_ (.A(message[334]),
    .B(_08599_),
    .Y(_08623_));
 sky130_fd_sc_hd__o21ai_0 _13434_ (.A1(_07731_),
    .A2(_08599_),
    .B1(_08623_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand2_1 _13435_ (.A(message[333]),
    .B(_08599_),
    .Y(_08624_));
 sky130_fd_sc_hd__o21ai_0 _13436_ (.A1(_07745_),
    .A2(_08599_),
    .B1(_08624_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_1 _13437_ (.A(message[332]),
    .B(_08599_),
    .Y(_08625_));
 sky130_fd_sc_hd__o21ai_0 _13438_ (.A1(_07752_),
    .A2(_08599_),
    .B1(_08625_),
    .Y(_00171_));
 sky130_fd_sc_hd__nand2_1 _13439_ (.A(message[331]),
    .B(_08599_),
    .Y(_08626_));
 sky130_fd_sc_hd__o21ai_0 _13440_ (.A1(_07766_),
    .A2(_08599_),
    .B1(_08626_),
    .Y(_00173_));
 sky130_fd_sc_hd__and2_1 _13441_ (.A(_05343_),
    .B(_08257_),
    .X(_08627_));
 sky130_fd_sc_hd__nor2_1 _13443_ (.A(message[330]),
    .B(_08627_),
    .Y(_08629_));
 sky130_fd_sc_hd__a21oi_1 _13444_ (.A1(_07777_),
    .A2(_08627_),
    .B1(_08629_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _13445_ (.A(message[329]),
    .B(_08599_),
    .Y(_08630_));
 sky130_fd_sc_hd__o21ai_0 _13446_ (.A1(_07786_),
    .A2(_08599_),
    .B1(_08630_),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _13447_ (.A(message[328]),
    .B(_08599_),
    .Y(_08631_));
 sky130_fd_sc_hd__o21ai_0 _13448_ (.A1(_07800_),
    .A2(_08599_),
    .B1(_08631_),
    .Y(_00176_));
 sky130_fd_sc_hd__nor2_1 _13449_ (.A(message[327]),
    .B(_08627_),
    .Y(_08632_));
 sky130_fd_sc_hd__a21oi_1 _13450_ (.A1(_07809_),
    .A2(_08627_),
    .B1(_08632_),
    .Y(_00177_));
 sky130_fd_sc_hd__nand2_1 _13451_ (.A(message[326]),
    .B(_08599_),
    .Y(_08633_));
 sky130_fd_sc_hd__o21ai_0 _13452_ (.A1(_07818_),
    .A2(_08599_),
    .B1(_08633_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _13453_ (.A(message[325]),
    .B(_08599_),
    .Y(_08634_));
 sky130_fd_sc_hd__o21ai_0 _13454_ (.A1(_07831_),
    .A2(_08599_),
    .B1(_08634_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _13455_ (.A(message[324]),
    .B(_08599_),
    .Y(_08635_));
 sky130_fd_sc_hd__o21ai_0 _13456_ (.A1(_07843_),
    .A2(_08599_),
    .B1(_08635_),
    .Y(_00180_));
 sky130_fd_sc_hd__nor2_1 _13457_ (.A(message[323]),
    .B(_08627_),
    .Y(_08636_));
 sky130_fd_sc_hd__a21oi_1 _13458_ (.A1(_07850_),
    .A2(_08627_),
    .B1(_08636_),
    .Y(_00181_));
 sky130_fd_sc_hd__nor2_1 _13459_ (.A(_07860_),
    .B(_08599_),
    .Y(_08637_));
 sky130_fd_sc_hd__a21oi_1 _13460_ (.A1(message[322]),
    .A2(_08599_),
    .B1(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__a21oi_1 _13461_ (.A1(_07859_),
    .A2(_08627_),
    .B1(_08638_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _13462_ (.A(message[321]),
    .B(_08599_),
    .Y(_08639_));
 sky130_fd_sc_hd__o21ai_0 _13463_ (.A1(_07873_),
    .A2(_08599_),
    .B1(_08639_),
    .Y(_00184_));
 sky130_fd_sc_hd__nor2_1 _13464_ (.A(message[320]),
    .B(_08627_),
    .Y(_08640_));
 sky130_fd_sc_hd__a21oi_1 _13465_ (.A1(_07925_),
    .A2(_08627_),
    .B1(_08640_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_1 _13466_ (.A(_05389_),
    .B(_08304_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand2_1 _13469_ (.A(message[383]),
    .B(_08641_),
    .Y(_08644_));
 sky130_fd_sc_hd__o21ai_0 _13470_ (.A1(_07930_),
    .A2(_08641_),
    .B1(_08644_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _13471_ (.A(message[382]),
    .B(_08641_),
    .Y(_08645_));
 sky130_fd_sc_hd__o21ai_0 _13472_ (.A1(_07934_),
    .A2(_08641_),
    .B1(_08645_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _13473_ (.A(message[381]),
    .B(_08641_),
    .Y(_08646_));
 sky130_fd_sc_hd__o21ai_0 _13474_ (.A1(_07937_),
    .A2(_08641_),
    .B1(_08646_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _13475_ (.A(message[380]),
    .B(_08641_),
    .Y(_08647_));
 sky130_fd_sc_hd__o21ai_0 _13476_ (.A1(_07942_),
    .A2(_08641_),
    .B1(_08647_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _13477_ (.A(message[379]),
    .B(_08641_),
    .Y(_08648_));
 sky130_fd_sc_hd__o21ai_0 _13478_ (.A1(_07949_),
    .A2(_08641_),
    .B1(_08648_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _13479_ (.A(message[378]),
    .B(_08641_),
    .Y(_08649_));
 sky130_fd_sc_hd__o21ai_0 _13480_ (.A1(_07956_),
    .A2(_08641_),
    .B1(_08649_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _13481_ (.A(message[377]),
    .B(_08641_),
    .Y(_08650_));
 sky130_fd_sc_hd__o21ai_0 _13482_ (.A1(_07965_),
    .A2(_08641_),
    .B1(_08650_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _13483_ (.A(message[376]),
    .B(_08641_),
    .Y(_08651_));
 sky130_fd_sc_hd__o21ai_0 _13484_ (.A1(_07974_),
    .A2(_08641_),
    .B1(_08651_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _13485_ (.A(message[375]),
    .B(_08641_),
    .Y(_08652_));
 sky130_fd_sc_hd__o21ai_0 _13486_ (.A1(_07981_),
    .A2(_08641_),
    .B1(_08652_),
    .Y(_00223_));
 sky130_fd_sc_hd__nand2_1 _13488_ (.A(message[374]),
    .B(_08641_),
    .Y(_08654_));
 sky130_fd_sc_hd__o21ai_0 _13489_ (.A1(_07989_),
    .A2(_08641_),
    .B1(_08654_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _13491_ (.A(message[373]),
    .B(_08641_),
    .Y(_08656_));
 sky130_fd_sc_hd__o21ai_0 _13492_ (.A1(_08006_),
    .A2(_08641_),
    .B1(_08656_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _13493_ (.A(message[372]),
    .B(_08641_),
    .Y(_08657_));
 sky130_fd_sc_hd__o21ai_0 _13494_ (.A1(_08018_),
    .A2(_08641_),
    .B1(_08657_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _13495_ (.A(message[371]),
    .B(_08641_),
    .Y(_08658_));
 sky130_fd_sc_hd__o21ai_0 _13496_ (.A1(_08025_),
    .A2(_08641_),
    .B1(_08658_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _13497_ (.A(message[370]),
    .B(_08641_),
    .Y(_08659_));
 sky130_fd_sc_hd__o21ai_0 _13498_ (.A1(_08031_),
    .A2(_08641_),
    .B1(_08659_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand2_1 _13499_ (.A(message[369]),
    .B(_08641_),
    .Y(_08660_));
 sky130_fd_sc_hd__o21ai_0 _13500_ (.A1(_08039_),
    .A2(_08641_),
    .B1(_08660_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _13501_ (.A(message[368]),
    .B(_08641_),
    .Y(_08661_));
 sky130_fd_sc_hd__o21ai_0 _13502_ (.A1(_08051_),
    .A2(_08641_),
    .B1(_08661_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _13503_ (.A(message[367]),
    .B(_08641_),
    .Y(_08662_));
 sky130_fd_sc_hd__o21ai_0 _13504_ (.A1(_08064_),
    .A2(_08641_),
    .B1(_08662_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _13505_ (.A(message[366]),
    .B(_08641_),
    .Y(_08663_));
 sky130_fd_sc_hd__o21ai_0 _13506_ (.A1(_08071_),
    .A2(_08641_),
    .B1(_08663_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _13507_ (.A(message[365]),
    .B(_08641_),
    .Y(_08664_));
 sky130_fd_sc_hd__o21ai_0 _13508_ (.A1(_08082_),
    .A2(_08641_),
    .B1(_08664_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _13510_ (.A(message[364]),
    .B(_08641_),
    .Y(_08666_));
 sky130_fd_sc_hd__o21ai_0 _13511_ (.A1(_08091_),
    .A2(_08641_),
    .B1(_08666_),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _13513_ (.A(message[363]),
    .B(_08641_),
    .Y(_08668_));
 sky130_fd_sc_hd__o21ai_0 _13514_ (.A1(_08102_),
    .A2(_08641_),
    .B1(_08668_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _13515_ (.A(message[362]),
    .B(_08641_),
    .Y(_08669_));
 sky130_fd_sc_hd__o21ai_0 _13516_ (.A1(_08114_),
    .A2(_08641_),
    .B1(_08669_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _13517_ (.A(message[361]),
    .B(_08641_),
    .Y(_08670_));
 sky130_fd_sc_hd__o21ai_0 _13518_ (.A1(_08125_),
    .A2(_08641_),
    .B1(_08670_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_1 _13519_ (.A(message[360]),
    .B(_08641_),
    .Y(_08671_));
 sky130_fd_sc_hd__o21ai_0 _13520_ (.A1(_08142_),
    .A2(_08641_),
    .B1(_08671_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _13521_ (.A(message[359]),
    .B(_08641_),
    .Y(_08672_));
 sky130_fd_sc_hd__o21ai_0 _13522_ (.A1(_08152_),
    .A2(_08641_),
    .B1(_08672_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _13523_ (.A(message[358]),
    .B(_08641_),
    .Y(_08673_));
 sky130_fd_sc_hd__o21ai_0 _13524_ (.A1(_08160_),
    .A2(_08641_),
    .B1(_08673_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _13525_ (.A(message[357]),
    .B(_08641_),
    .Y(_08674_));
 sky130_fd_sc_hd__o21ai_0 _13526_ (.A1(_08171_),
    .A2(_08641_),
    .B1(_08674_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _13527_ (.A(message[356]),
    .B(_08641_),
    .Y(_08675_));
 sky130_fd_sc_hd__o21ai_0 _13528_ (.A1(_08184_),
    .A2(_08641_),
    .B1(_08675_),
    .Y(_00212_));
 sky130_fd_sc_hd__a21oi_1 _13529_ (.A1(_05389_),
    .A2(_08304_),
    .B1(message[355]),
    .Y(_08676_));
 sky130_fd_sc_hd__a31oi_1 _13530_ (.A1(_05389_),
    .A2(_08204_),
    .A3(_08304_),
    .B1(_08676_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _13531_ (.A(message[354]),
    .B(_08641_),
    .Y(_08677_));
 sky130_fd_sc_hd__o21ai_0 _13532_ (.A1(_08209_),
    .A2(_08641_),
    .B1(_08677_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _13533_ (.A(message[353]),
    .B(_08641_),
    .Y(_08678_));
 sky130_fd_sc_hd__o21ai_0 _13534_ (.A1(_08221_),
    .A2(_08641_),
    .B1(_08678_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _13535_ (.A(message[352]),
    .B(_08641_),
    .Y(_08679_));
 sky130_fd_sc_hd__o21ai_1 _13536_ (.A1(_08254_),
    .A2(_08641_),
    .B1(_08679_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _13537_ (.A(_05343_),
    .B(_08346_),
    .Y(_08680_));
 sky130_fd_sc_hd__nand2_1 _13541_ (.A(message[415]),
    .B(_08680_),
    .Y(_08684_));
 sky130_fd_sc_hd__o21ai_0 _13542_ (.A1(_07572_),
    .A2(_08680_),
    .B1(_08684_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _13543_ (.A(message[414]),
    .B(_08680_),
    .Y(_08685_));
 sky130_fd_sc_hd__o21ai_0 _13544_ (.A1(_07577_),
    .A2(_08680_),
    .B1(_08685_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _13545_ (.A(message[413]),
    .B(_08680_),
    .Y(_08686_));
 sky130_fd_sc_hd__o21ai_0 _13546_ (.A1(_07581_),
    .A2(_08680_),
    .B1(_08686_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _13548_ (.A(message[412]),
    .B(_08680_),
    .Y(_08688_));
 sky130_fd_sc_hd__o21ai_0 _13549_ (.A1(_07588_),
    .A2(_08680_),
    .B1(_08688_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _13550_ (.A(message[411]),
    .B(_08680_),
    .Y(_08689_));
 sky130_fd_sc_hd__o21ai_0 _13551_ (.A1(_07601_),
    .A2(_08680_),
    .B1(_08689_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _13552_ (.A(message[410]),
    .B(_08680_),
    .Y(_08690_));
 sky130_fd_sc_hd__o21ai_0 _13553_ (.A1(_07610_),
    .A2(_08680_),
    .B1(_08690_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _13554_ (.A(message[409]),
    .B(_08680_),
    .Y(_08691_));
 sky130_fd_sc_hd__o21ai_0 _13555_ (.A1(_07620_),
    .A2(_08680_),
    .B1(_08691_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _13556_ (.A(message[408]),
    .B(_08680_),
    .Y(_08692_));
 sky130_fd_sc_hd__o21ai_0 _13557_ (.A1(_07628_),
    .A2(_08680_),
    .B1(_08692_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(message[407]),
    .B(_08680_),
    .Y(_08693_));
 sky130_fd_sc_hd__o21ai_0 _13559_ (.A1(_07635_),
    .A2(_08680_),
    .B1(_08693_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _13560_ (.A(message[406]),
    .B(_08680_),
    .Y(_08694_));
 sky130_fd_sc_hd__o21ai_0 _13561_ (.A1(_07646_),
    .A2(_08680_),
    .B1(_08694_),
    .Y(_00256_));
 sky130_fd_sc_hd__nand2_1 _13563_ (.A(message[405]),
    .B(_08680_),
    .Y(_08696_));
 sky130_fd_sc_hd__o21ai_0 _13564_ (.A1(_07660_),
    .A2(_08680_),
    .B1(_08696_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _13565_ (.A(message[404]),
    .B(_08680_),
    .Y(_08697_));
 sky130_fd_sc_hd__o21ai_0 _13566_ (.A1(_07669_),
    .A2(_08680_),
    .B1(_08697_),
    .Y(_00227_));
 sky130_fd_sc_hd__and2_1 _13567_ (.A(_05343_),
    .B(_08346_),
    .X(_08698_));
 sky130_fd_sc_hd__nor2_1 _13569_ (.A(message[403]),
    .B(_08698_),
    .Y(_08700_));
 sky130_fd_sc_hd__a21oi_1 _13570_ (.A1(_07677_),
    .A2(_08698_),
    .B1(_08700_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _13571_ (.A(message[402]),
    .B(_08680_),
    .Y(_08701_));
 sky130_fd_sc_hd__o21ai_0 _13572_ (.A1(_07689_),
    .A2(_08680_),
    .B1(_08701_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _13574_ (.A(message[401]),
    .B(_08680_),
    .Y(_08703_));
 sky130_fd_sc_hd__o21ai_0 _13575_ (.A1(_07703_),
    .A2(_08680_),
    .B1(_08703_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _13576_ (.A(message[400]),
    .B(_08680_),
    .Y(_08704_));
 sky130_fd_sc_hd__o21ai_0 _13577_ (.A1(_07709_),
    .A2(_08680_),
    .B1(_08704_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _13578_ (.A(message[399]),
    .B(_08680_),
    .Y(_08705_));
 sky130_fd_sc_hd__o21ai_0 _13579_ (.A1(_07715_),
    .A2(_08680_),
    .B1(_08705_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _13580_ (.A(message[398]),
    .B(_08680_),
    .Y(_08706_));
 sky130_fd_sc_hd__o21ai_0 _13581_ (.A1(_07731_),
    .A2(_08680_),
    .B1(_08706_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand2_1 _13582_ (.A(message[397]),
    .B(_08680_),
    .Y(_08707_));
 sky130_fd_sc_hd__o21ai_0 _13583_ (.A1(_07745_),
    .A2(_08680_),
    .B1(_08707_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _13584_ (.A(message[396]),
    .B(_08680_),
    .Y(_08708_));
 sky130_fd_sc_hd__o21ai_0 _13585_ (.A1(_07752_),
    .A2(_08680_),
    .B1(_08708_),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_1 _13586_ (.A(message[395]),
    .B(_08680_),
    .Y(_08709_));
 sky130_fd_sc_hd__o21ai_0 _13587_ (.A1(_07766_),
    .A2(_08680_),
    .B1(_08709_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _13588_ (.A(message[394]),
    .B(_08680_),
    .Y(_08710_));
 sky130_fd_sc_hd__o21ai_0 _13589_ (.A1(_07777_),
    .A2(_08680_),
    .B1(_08710_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _13590_ (.A(message[393]),
    .B(_08680_),
    .Y(_08711_));
 sky130_fd_sc_hd__o21ai_0 _13591_ (.A1(_07786_),
    .A2(_08680_),
    .B1(_08711_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _13592_ (.A(message[392]),
    .B(_08680_),
    .Y(_08712_));
 sky130_fd_sc_hd__o21ai_0 _13593_ (.A1(_07800_),
    .A2(_08680_),
    .B1(_08712_),
    .Y(_00240_));
 sky130_fd_sc_hd__nor2_1 _13594_ (.A(message[391]),
    .B(_08698_),
    .Y(_08713_));
 sky130_fd_sc_hd__a21oi_1 _13595_ (.A1(_07809_),
    .A2(_08698_),
    .B1(_08713_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _13596_ (.A(message[390]),
    .B(_08680_),
    .Y(_08714_));
 sky130_fd_sc_hd__o21ai_0 _13597_ (.A1(_07818_),
    .A2(_08680_),
    .B1(_08714_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _13598_ (.A(message[389]),
    .B(_08680_),
    .Y(_08715_));
 sky130_fd_sc_hd__o21ai_0 _13599_ (.A1(_07831_),
    .A2(_08680_),
    .B1(_08715_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _13600_ (.A(message[388]),
    .B(_08680_),
    .Y(_08716_));
 sky130_fd_sc_hd__o21ai_0 _13601_ (.A1(_07843_),
    .A2(_08680_),
    .B1(_08716_),
    .Y(_00244_));
 sky130_fd_sc_hd__nor2_1 _13602_ (.A(message[387]),
    .B(_08698_),
    .Y(_08717_));
 sky130_fd_sc_hd__a21oi_1 _13603_ (.A1(_07850_),
    .A2(_08698_),
    .B1(_08717_),
    .Y(_00245_));
 sky130_fd_sc_hd__nor2_1 _13604_ (.A(_07860_),
    .B(_08680_),
    .Y(_08718_));
 sky130_fd_sc_hd__a21oi_1 _13605_ (.A1(message[386]),
    .A2(_08680_),
    .B1(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__a21oi_1 _13606_ (.A1(_07859_),
    .A2(_08698_),
    .B1(_08719_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _13607_ (.A(message[385]),
    .B(_08680_),
    .Y(_08720_));
 sky130_fd_sc_hd__o21ai_0 _13608_ (.A1(_07873_),
    .A2(_08680_),
    .B1(_08720_),
    .Y(_00248_));
 sky130_fd_sc_hd__nor2_1 _13609_ (.A(message[384]),
    .B(_08698_),
    .Y(_08721_));
 sky130_fd_sc_hd__a21oi_1 _13610_ (.A1(_07925_),
    .A2(_08698_),
    .B1(_08721_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_1 _13611_ (.A(_05389_),
    .B(_08390_),
    .Y(_08722_));
 sky130_fd_sc_hd__nand2_1 _13614_ (.A(message[447]),
    .B(_08722_),
    .Y(_08725_));
 sky130_fd_sc_hd__o21ai_0 _13615_ (.A1(_07930_),
    .A2(_08722_),
    .B1(_08725_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _13616_ (.A(message[446]),
    .B(_08722_),
    .Y(_08726_));
 sky130_fd_sc_hd__o21ai_0 _13617_ (.A1(_07934_),
    .A2(_08722_),
    .B1(_08726_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _13618_ (.A(message[445]),
    .B(_08722_),
    .Y(_08727_));
 sky130_fd_sc_hd__o21ai_0 _13619_ (.A1(_07937_),
    .A2(_08722_),
    .B1(_08727_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _13620_ (.A(message[444]),
    .B(_08722_),
    .Y(_08728_));
 sky130_fd_sc_hd__o21ai_0 _13621_ (.A1(_07942_),
    .A2(_08722_),
    .B1(_08728_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _13622_ (.A(message[443]),
    .B(_08722_),
    .Y(_08729_));
 sky130_fd_sc_hd__o21ai_0 _13623_ (.A1(_07949_),
    .A2(_08722_),
    .B1(_08729_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _13624_ (.A(message[442]),
    .B(_08722_),
    .Y(_08730_));
 sky130_fd_sc_hd__o21ai_0 _13625_ (.A1(_07956_),
    .A2(_08722_),
    .B1(_08730_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _13626_ (.A(message[441]),
    .B(_08722_),
    .Y(_08731_));
 sky130_fd_sc_hd__o21ai_0 _13627_ (.A1(_07965_),
    .A2(_08722_),
    .B1(_08731_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _13628_ (.A(message[440]),
    .B(_08722_),
    .Y(_08732_));
 sky130_fd_sc_hd__o21ai_0 _13629_ (.A1(_07974_),
    .A2(_08722_),
    .B1(_08732_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _13630_ (.A(message[439]),
    .B(_08722_),
    .Y(_08733_));
 sky130_fd_sc_hd__o21ai_0 _13631_ (.A1(_07981_),
    .A2(_08722_),
    .B1(_08733_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _13633_ (.A(message[438]),
    .B(_08722_),
    .Y(_08735_));
 sky130_fd_sc_hd__o21ai_0 _13634_ (.A1(_07989_),
    .A2(_08722_),
    .B1(_08735_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand2_1 _13636_ (.A(message[437]),
    .B(_08722_),
    .Y(_08737_));
 sky130_fd_sc_hd__o21ai_0 _13637_ (.A1(_08006_),
    .A2(_08722_),
    .B1(_08737_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _13638_ (.A(message[436]),
    .B(_08722_),
    .Y(_08738_));
 sky130_fd_sc_hd__o21ai_0 _13639_ (.A1(_08018_),
    .A2(_08722_),
    .B1(_08738_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _13640_ (.A(message[435]),
    .B(_08722_),
    .Y(_08739_));
 sky130_fd_sc_hd__o21ai_0 _13641_ (.A1(_08025_),
    .A2(_08722_),
    .B1(_08739_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _13642_ (.A(message[434]),
    .B(_08722_),
    .Y(_08740_));
 sky130_fd_sc_hd__o21ai_0 _13643_ (.A1(_08031_),
    .A2(_08722_),
    .B1(_08740_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _13644_ (.A(message[433]),
    .B(_08722_),
    .Y(_08741_));
 sky130_fd_sc_hd__o21ai_0 _13645_ (.A1(_08039_),
    .A2(_08722_),
    .B1(_08741_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _13646_ (.A(message[432]),
    .B(_08722_),
    .Y(_08742_));
 sky130_fd_sc_hd__o21ai_0 _13647_ (.A1(_08051_),
    .A2(_08722_),
    .B1(_08742_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _13648_ (.A(message[431]),
    .B(_08722_),
    .Y(_08743_));
 sky130_fd_sc_hd__o21ai_0 _13649_ (.A1(_08064_),
    .A2(_08722_),
    .B1(_08743_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _13650_ (.A(message[430]),
    .B(_08722_),
    .Y(_08744_));
 sky130_fd_sc_hd__o21ai_0 _13651_ (.A1(_08071_),
    .A2(_08722_),
    .B1(_08744_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _13652_ (.A(message[429]),
    .B(_08722_),
    .Y(_08745_));
 sky130_fd_sc_hd__o21ai_0 _13653_ (.A1(_08082_),
    .A2(_08722_),
    .B1(_08745_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_1 _13655_ (.A(message[428]),
    .B(_08722_),
    .Y(_08747_));
 sky130_fd_sc_hd__o21ai_0 _13656_ (.A1(_08091_),
    .A2(_08722_),
    .B1(_08747_),
    .Y(_00267_));
 sky130_fd_sc_hd__nand2_1 _13658_ (.A(message[427]),
    .B(_08722_),
    .Y(_08749_));
 sky130_fd_sc_hd__o21ai_0 _13659_ (.A1(_08102_),
    .A2(_08722_),
    .B1(_08749_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _13660_ (.A(message[426]),
    .B(_08722_),
    .Y(_08750_));
 sky130_fd_sc_hd__o21ai_0 _13661_ (.A1(_08114_),
    .A2(_08722_),
    .B1(_08750_),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _13662_ (.A(message[425]),
    .B(_08722_),
    .Y(_08751_));
 sky130_fd_sc_hd__o21ai_0 _13663_ (.A1(_08125_),
    .A2(_08722_),
    .B1(_08751_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _13664_ (.A(message[424]),
    .B(_08722_),
    .Y(_08752_));
 sky130_fd_sc_hd__o21ai_0 _13665_ (.A1(_08142_),
    .A2(_08722_),
    .B1(_08752_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _13666_ (.A(message[423]),
    .B(_08722_),
    .Y(_08753_));
 sky130_fd_sc_hd__o21ai_0 _13667_ (.A1(_08152_),
    .A2(_08722_),
    .B1(_08753_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _13668_ (.A(message[422]),
    .B(_08722_),
    .Y(_08754_));
 sky130_fd_sc_hd__o21ai_0 _13669_ (.A1(_08160_),
    .A2(_08722_),
    .B1(_08754_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _13670_ (.A(message[421]),
    .B(_08722_),
    .Y(_08755_));
 sky130_fd_sc_hd__o21ai_0 _13671_ (.A1(_08171_),
    .A2(_08722_),
    .B1(_08755_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _13672_ (.A(message[420]),
    .B(_08722_),
    .Y(_08756_));
 sky130_fd_sc_hd__o21ai_0 _13673_ (.A1(_08184_),
    .A2(_08722_),
    .B1(_08756_),
    .Y(_00276_));
 sky130_fd_sc_hd__a21oi_1 _13674_ (.A1(_05389_),
    .A2(_08390_),
    .B1(message[419]),
    .Y(_08757_));
 sky130_fd_sc_hd__a31oi_1 _13675_ (.A1(_05389_),
    .A2(_08204_),
    .A3(_08390_),
    .B1(_08757_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _13676_ (.A(message[418]),
    .B(_08722_),
    .Y(_08758_));
 sky130_fd_sc_hd__o21ai_0 _13677_ (.A1(_08209_),
    .A2(_08722_),
    .B1(_08758_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _13678_ (.A(message[417]),
    .B(_08722_),
    .Y(_08759_));
 sky130_fd_sc_hd__o21ai_0 _13679_ (.A1(_08221_),
    .A2(_08722_),
    .B1(_08759_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _13680_ (.A(message[416]),
    .B(_08722_),
    .Y(_08760_));
 sky130_fd_sc_hd__o21ai_0 _13681_ (.A1(_08254_),
    .A2(_08722_),
    .B1(_08760_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _13682_ (.A(_05343_),
    .B(_08431_),
    .Y(_08761_));
 sky130_fd_sc_hd__nand2_1 _13685_ (.A(message[479]),
    .B(_08761_),
    .Y(_08764_));
 sky130_fd_sc_hd__o21ai_0 _13686_ (.A1(_07572_),
    .A2(_08761_),
    .B1(_08764_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _13687_ (.A(message[478]),
    .B(_08761_),
    .Y(_08765_));
 sky130_fd_sc_hd__o21ai_0 _13688_ (.A1(_07577_),
    .A2(_08761_),
    .B1(_08765_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _13691_ (.A(message[477]),
    .B(_08761_),
    .Y(_08768_));
 sky130_fd_sc_hd__o21ai_0 _13692_ (.A1(_07581_),
    .A2(_08761_),
    .B1(_08768_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _13693_ (.A(message[476]),
    .B(_08761_),
    .Y(_08769_));
 sky130_fd_sc_hd__o21ai_0 _13694_ (.A1(_07588_),
    .A2(_08761_),
    .B1(_08769_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _13695_ (.A(message[475]),
    .B(_08761_),
    .Y(_08770_));
 sky130_fd_sc_hd__o21ai_0 _13696_ (.A1(_07601_),
    .A2(_08761_),
    .B1(_08770_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _13697_ (.A(message[474]),
    .B(_08761_),
    .Y(_08771_));
 sky130_fd_sc_hd__o21ai_0 _13698_ (.A1(_07610_),
    .A2(_08761_),
    .B1(_08771_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _13699_ (.A(message[473]),
    .B(_08761_),
    .Y(_08772_));
 sky130_fd_sc_hd__o21ai_0 _13700_ (.A1(_07620_),
    .A2(_08761_),
    .B1(_08772_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _13701_ (.A(message[472]),
    .B(_08761_),
    .Y(_08773_));
 sky130_fd_sc_hd__o21ai_0 _13702_ (.A1(_07628_),
    .A2(_08761_),
    .B1(_08773_),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_1 _13703_ (.A(message[471]),
    .B(_08761_),
    .Y(_08774_));
 sky130_fd_sc_hd__o21ai_0 _13704_ (.A1(_07635_),
    .A2(_08761_),
    .B1(_08774_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _13705_ (.A(message[470]),
    .B(_08761_),
    .Y(_08775_));
 sky130_fd_sc_hd__o21ai_0 _13706_ (.A1(_07646_),
    .A2(_08761_),
    .B1(_08775_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _13708_ (.A(message[469]),
    .B(_08761_),
    .Y(_08777_));
 sky130_fd_sc_hd__o21ai_0 _13709_ (.A1(_07660_),
    .A2(_08761_),
    .B1(_08777_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _13710_ (.A(message[468]),
    .B(_08761_),
    .Y(_08778_));
 sky130_fd_sc_hd__o21ai_0 _13711_ (.A1(_07669_),
    .A2(_08761_),
    .B1(_08778_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _13713_ (.A(message[467]),
    .B(_08761_),
    .Y(_08780_));
 sky130_fd_sc_hd__o21ai_0 _13714_ (.A1(_07677_),
    .A2(_08761_),
    .B1(_08780_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _13715_ (.A(message[466]),
    .B(_08761_),
    .Y(_08781_));
 sky130_fd_sc_hd__o21ai_0 _13716_ (.A1(_07689_),
    .A2(_08761_),
    .B1(_08781_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _13717_ (.A(message[465]),
    .B(_08761_),
    .Y(_08782_));
 sky130_fd_sc_hd__o21ai_0 _13718_ (.A1(_07703_),
    .A2(_08761_),
    .B1(_08782_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _13719_ (.A(message[464]),
    .B(_08761_),
    .Y(_08783_));
 sky130_fd_sc_hd__o21ai_0 _13720_ (.A1(_07709_),
    .A2(_08761_),
    .B1(_08783_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _13721_ (.A(message[463]),
    .B(_08761_),
    .Y(_08784_));
 sky130_fd_sc_hd__o21ai_0 _13722_ (.A1(_07715_),
    .A2(_08761_),
    .B1(_08784_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _13723_ (.A(message[462]),
    .B(_08761_),
    .Y(_08785_));
 sky130_fd_sc_hd__o21ai_0 _13724_ (.A1(_07731_),
    .A2(_08761_),
    .B1(_08785_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _13725_ (.A(message[461]),
    .B(_08761_),
    .Y(_08786_));
 sky130_fd_sc_hd__o21ai_0 _13726_ (.A1(_07745_),
    .A2(_08761_),
    .B1(_08786_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _13727_ (.A(message[460]),
    .B(_08761_),
    .Y(_08787_));
 sky130_fd_sc_hd__o21ai_0 _13728_ (.A1(_07752_),
    .A2(_08761_),
    .B1(_08787_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _13729_ (.A(message[459]),
    .B(_08761_),
    .Y(_08788_));
 sky130_fd_sc_hd__o21ai_0 _13730_ (.A1(_07766_),
    .A2(_08761_),
    .B1(_08788_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _13731_ (.A(message[458]),
    .B(_08761_),
    .Y(_08789_));
 sky130_fd_sc_hd__o21ai_0 _13732_ (.A1(_07777_),
    .A2(_08761_),
    .B1(_08789_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _13733_ (.A(message[457]),
    .B(_08761_),
    .Y(_08790_));
 sky130_fd_sc_hd__o21ai_0 _13734_ (.A1(_07786_),
    .A2(_08761_),
    .B1(_08790_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _13735_ (.A(message[456]),
    .B(_08761_),
    .Y(_08791_));
 sky130_fd_sc_hd__o21ai_0 _13736_ (.A1(_07800_),
    .A2(_08761_),
    .B1(_08791_),
    .Y(_00304_));
 sky130_fd_sc_hd__and2_1 _13737_ (.A(_05343_),
    .B(_08431_),
    .X(_08792_));
 sky130_fd_sc_hd__nor2_1 _13739_ (.A(message[455]),
    .B(_08792_),
    .Y(_08794_));
 sky130_fd_sc_hd__a21oi_1 _13740_ (.A1(_07809_),
    .A2(_08792_),
    .B1(_08794_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _13741_ (.A(message[454]),
    .B(_08761_),
    .Y(_08795_));
 sky130_fd_sc_hd__o21ai_0 _13742_ (.A1(_07818_),
    .A2(_08761_),
    .B1(_08795_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _13743_ (.A(message[453]),
    .B(_08761_),
    .Y(_08796_));
 sky130_fd_sc_hd__o21ai_0 _13744_ (.A1(_07831_),
    .A2(_08761_),
    .B1(_08796_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _13745_ (.A(message[452]),
    .B(_08761_),
    .Y(_08797_));
 sky130_fd_sc_hd__o21ai_0 _13746_ (.A1(_07843_),
    .A2(_08761_),
    .B1(_08797_),
    .Y(_00308_));
 sky130_fd_sc_hd__nor2_1 _13747_ (.A(message[451]),
    .B(_08792_),
    .Y(_08798_));
 sky130_fd_sc_hd__a21oi_1 _13748_ (.A1(_07850_),
    .A2(_08792_),
    .B1(_08798_),
    .Y(_00309_));
 sky130_fd_sc_hd__nor2_1 _13749_ (.A(_07860_),
    .B(_08761_),
    .Y(_08799_));
 sky130_fd_sc_hd__a21oi_1 _13750_ (.A1(message[450]),
    .A2(_08761_),
    .B1(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__a21oi_1 _13751_ (.A1(_07859_),
    .A2(_08792_),
    .B1(_08800_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _13752_ (.A(message[449]),
    .B(_08761_),
    .Y(_08801_));
 sky130_fd_sc_hd__o21ai_0 _13753_ (.A1(_07873_),
    .A2(_08761_),
    .B1(_08801_),
    .Y(_00312_));
 sky130_fd_sc_hd__nor2_1 _13754_ (.A(message[448]),
    .B(_08792_),
    .Y(_08802_));
 sky130_fd_sc_hd__a21oi_1 _13755_ (.A1(_07925_),
    .A2(_08792_),
    .B1(_08802_),
    .Y(_00313_));
 sky130_fd_sc_hd__nor2b_1 _13756_ (.A(reset),
    .B_N(_09567_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand2_1 _13757_ (.A(_05389_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__nand2_1 _13760_ (.A(message[511]),
    .B(_08804_),
    .Y(_08807_));
 sky130_fd_sc_hd__o21ai_0 _13761_ (.A1(_07930_),
    .A2(_08804_),
    .B1(_08807_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _13762_ (.A(message[510]),
    .B(_08804_),
    .Y(_08808_));
 sky130_fd_sc_hd__o21ai_0 _13763_ (.A1(_07934_),
    .A2(_08804_),
    .B1(_08808_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _13764_ (.A(message[509]),
    .B(_08804_),
    .Y(_08809_));
 sky130_fd_sc_hd__o21ai_0 _13765_ (.A1(_07937_),
    .A2(_08804_),
    .B1(_08809_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _13766_ (.A(message[508]),
    .B(_08804_),
    .Y(_08810_));
 sky130_fd_sc_hd__o21ai_0 _13767_ (.A1(_07942_),
    .A2(_08804_),
    .B1(_08810_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _13768_ (.A(message[507]),
    .B(_08804_),
    .Y(_08811_));
 sky130_fd_sc_hd__o21ai_0 _13769_ (.A1(_07949_),
    .A2(_08804_),
    .B1(_08811_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _13770_ (.A(message[506]),
    .B(_08804_),
    .Y(_08812_));
 sky130_fd_sc_hd__o21ai_0 _13771_ (.A1(_07956_),
    .A2(_08804_),
    .B1(_08812_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _13772_ (.A(message[505]),
    .B(_08804_),
    .Y(_08813_));
 sky130_fd_sc_hd__o21ai_0 _13773_ (.A1(_07965_),
    .A2(_08804_),
    .B1(_08813_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _13774_ (.A(message[504]),
    .B(_08804_),
    .Y(_08814_));
 sky130_fd_sc_hd__o21ai_0 _13775_ (.A1(_07974_),
    .A2(_08804_),
    .B1(_08814_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _13776_ (.A(message[503]),
    .B(_08804_),
    .Y(_08815_));
 sky130_fd_sc_hd__o21ai_0 _13777_ (.A1(_07981_),
    .A2(_08804_),
    .B1(_08815_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _13779_ (.A(message[502]),
    .B(_08804_),
    .Y(_08817_));
 sky130_fd_sc_hd__o21ai_0 _13780_ (.A1(_07989_),
    .A2(_08804_),
    .B1(_08817_),
    .Y(_00352_));
 sky130_fd_sc_hd__nand2_1 _13782_ (.A(message[501]),
    .B(_08804_),
    .Y(_08819_));
 sky130_fd_sc_hd__o21ai_0 _13783_ (.A1(_08006_),
    .A2(_08804_),
    .B1(_08819_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(message[500]),
    .B(_08804_),
    .Y(_08820_));
 sky130_fd_sc_hd__o21ai_0 _13785_ (.A1(_08018_),
    .A2(_08804_),
    .B1(_08820_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _13786_ (.A(message[499]),
    .B(_08804_),
    .Y(_08821_));
 sky130_fd_sc_hd__o21ai_0 _13787_ (.A1(_08025_),
    .A2(_08804_),
    .B1(_08821_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _13788_ (.A(message[498]),
    .B(_08804_),
    .Y(_02321_));
 sky130_fd_sc_hd__o21ai_0 _13789_ (.A1(_08031_),
    .A2(_08804_),
    .B1(_02321_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _13790_ (.A(message[497]),
    .B(_08804_),
    .Y(_02322_));
 sky130_fd_sc_hd__o21ai_0 _13791_ (.A1(_08039_),
    .A2(_08804_),
    .B1(_02322_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _13792_ (.A(message[496]),
    .B(_08804_),
    .Y(_02323_));
 sky130_fd_sc_hd__o21ai_0 _13793_ (.A1(_08051_),
    .A2(_08804_),
    .B1(_02323_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _13794_ (.A(message[495]),
    .B(_08804_),
    .Y(_02324_));
 sky130_fd_sc_hd__o21ai_0 _13795_ (.A1(_08064_),
    .A2(_08804_),
    .B1(_02324_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _13796_ (.A(message[494]),
    .B(_08804_),
    .Y(_02325_));
 sky130_fd_sc_hd__o21ai_0 _13797_ (.A1(_08071_),
    .A2(_08804_),
    .B1(_02325_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _13798_ (.A(message[493]),
    .B(_08804_),
    .Y(_02326_));
 sky130_fd_sc_hd__o21ai_0 _13799_ (.A1(_08082_),
    .A2(_08804_),
    .B1(_02326_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _13801_ (.A(message[492]),
    .B(_08804_),
    .Y(_02328_));
 sky130_fd_sc_hd__o21ai_0 _13802_ (.A1(_08091_),
    .A2(_08804_),
    .B1(_02328_),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _13804_ (.A(message[491]),
    .B(_08804_),
    .Y(_02330_));
 sky130_fd_sc_hd__o21ai_0 _13805_ (.A1(_08102_),
    .A2(_08804_),
    .B1(_02330_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _13806_ (.A(message[490]),
    .B(_08804_),
    .Y(_02331_));
 sky130_fd_sc_hd__o21ai_0 _13807_ (.A1(_08114_),
    .A2(_08804_),
    .B1(_02331_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _13808_ (.A(message[489]),
    .B(_08804_),
    .Y(_02332_));
 sky130_fd_sc_hd__o21ai_0 _13809_ (.A1(_08125_),
    .A2(_08804_),
    .B1(_02332_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _13810_ (.A(message[488]),
    .B(_08804_),
    .Y(_02333_));
 sky130_fd_sc_hd__o21ai_0 _13811_ (.A1(_08142_),
    .A2(_08804_),
    .B1(_02333_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _13812_ (.A(message[487]),
    .B(_08804_),
    .Y(_02334_));
 sky130_fd_sc_hd__o21ai_0 _13813_ (.A1(_08152_),
    .A2(_08804_),
    .B1(_02334_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _13814_ (.A(message[486]),
    .B(_08804_),
    .Y(_02335_));
 sky130_fd_sc_hd__o21ai_0 _13815_ (.A1(_08160_),
    .A2(_08804_),
    .B1(_02335_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _13816_ (.A(message[485]),
    .B(_08804_),
    .Y(_02336_));
 sky130_fd_sc_hd__o21ai_0 _13817_ (.A1(_08171_),
    .A2(_08804_),
    .B1(_02336_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _13818_ (.A(message[484]),
    .B(_08804_),
    .Y(_02337_));
 sky130_fd_sc_hd__o21ai_0 _13819_ (.A1(_08184_),
    .A2(_08804_),
    .B1(_02337_),
    .Y(_00340_));
 sky130_fd_sc_hd__a21oi_1 _13820_ (.A1(_05389_),
    .A2(_08803_),
    .B1(message[483]),
    .Y(_02338_));
 sky130_fd_sc_hd__a31oi_1 _13821_ (.A1(_05389_),
    .A2(_08204_),
    .A3(_08803_),
    .B1(_02338_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _13822_ (.A(message[482]),
    .B(_08804_),
    .Y(_02339_));
 sky130_fd_sc_hd__o21ai_0 _13823_ (.A1(_08209_),
    .A2(_08804_),
    .B1(_02339_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_1 _13824_ (.A(message[481]),
    .B(_08804_),
    .Y(_02340_));
 sky130_fd_sc_hd__o21ai_0 _13825_ (.A1(_08221_),
    .A2(_08804_),
    .B1(_02340_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _13826_ (.A(message[480]),
    .B(_08804_),
    .Y(_02341_));
 sky130_fd_sc_hd__o21ai_0 _13827_ (.A1(_08254_),
    .A2(_08804_),
    .B1(_02341_),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_1 _13828_ (.A(\w_new_calc2.temp2[0] ),
    .Y(_09070_));
 sky130_fd_sc_hd__inv_1 _13829_ (.A(\w_new_calc2.temp2[1] ),
    .Y(_09075_));
 sky130_fd_sc_hd__inv_1 _13830_ (.A(\w_new_calc2.temp2[2] ),
    .Y(_09084_));
 sky130_fd_sc_hd__inv_1 _13831_ (.A(\w_new_calc2.temp2[3] ),
    .Y(_09096_));
 sky130_fd_sc_hd__inv_1 _13832_ (.A(\w_new_calc2.temp2[4] ),
    .Y(_09105_));
 sky130_fd_sc_hd__inv_1 _13833_ (.A(\w_new_calc2.temp2[5] ),
    .Y(_09114_));
 sky130_fd_sc_hd__inv_1 _13834_ (.A(\w_new_calc2.temp2[6] ),
    .Y(_09123_));
 sky130_fd_sc_hd__inv_1 _13835_ (.A(\w_new_calc2.temp2[7] ),
    .Y(_09132_));
 sky130_fd_sc_hd__inv_1 _13836_ (.A(\w_new_calc2.temp2[8] ),
    .Y(_09141_));
 sky130_fd_sc_hd__inv_1 _13837_ (.A(\w_new_calc2.temp2[9] ),
    .Y(_09150_));
 sky130_fd_sc_hd__inv_1 _13838_ (.A(\w_new_calc2.temp2[10] ),
    .Y(_09159_));
 sky130_fd_sc_hd__inv_1 _13839_ (.A(\w_new_calc2.temp2[11] ),
    .Y(_09168_));
 sky130_fd_sc_hd__inv_1 _13840_ (.A(\w_new_calc2.temp2[12] ),
    .Y(_09177_));
 sky130_fd_sc_hd__inv_1 _13841_ (.A(\w_new_calc2.temp2[13] ),
    .Y(_09186_));
 sky130_fd_sc_hd__inv_1 _13842_ (.A(\w_new_calc2.temp2[14] ),
    .Y(_09195_));
 sky130_fd_sc_hd__inv_1 _13843_ (.A(\w_new_calc2.temp2[15] ),
    .Y(_09204_));
 sky130_fd_sc_hd__inv_1 _13844_ (.A(\w_new_calc2.temp2[16] ),
    .Y(_09213_));
 sky130_fd_sc_hd__inv_1 _13845_ (.A(\w_new_calc2.temp2[17] ),
    .Y(_09222_));
 sky130_fd_sc_hd__inv_1 _13846_ (.A(\w_new_calc2.temp2[18] ),
    .Y(_09231_));
 sky130_fd_sc_hd__inv_1 _13847_ (.A(\w_new_calc2.temp2[19] ),
    .Y(_09240_));
 sky130_fd_sc_hd__inv_1 _13848_ (.A(\w_new_calc2.temp2[20] ),
    .Y(_09249_));
 sky130_fd_sc_hd__inv_1 _13849_ (.A(\w_new_calc2.temp2[21] ),
    .Y(_09258_));
 sky130_fd_sc_hd__inv_1 _13850_ (.A(\w_new_calc2.temp2[22] ),
    .Y(_09267_));
 sky130_fd_sc_hd__inv_1 _13851_ (.A(\w_new_calc2.temp2[23] ),
    .Y(_09276_));
 sky130_fd_sc_hd__inv_1 _13852_ (.A(\w_new_calc2.temp2[24] ),
    .Y(_09285_));
 sky130_fd_sc_hd__inv_1 _13853_ (.A(\w_new_calc2.temp2[25] ),
    .Y(_09294_));
 sky130_fd_sc_hd__inv_1 _13854_ (.A(\w_new_calc2.temp2[26] ),
    .Y(_09303_));
 sky130_fd_sc_hd__inv_1 _13855_ (.A(\w_new_calc2.temp2[27] ),
    .Y(_09312_));
 sky130_fd_sc_hd__inv_1 _13856_ (.A(\w_new_calc2.temp1[28] ),
    .Y(_09325_));
 sky130_fd_sc_hd__inv_1 _13857_ (.A(\w_new_calc2.temp1[29] ),
    .Y(_09333_));
 sky130_fd_sc_hd__inv_1 _13858_ (.A(\w_new_calc2.temp2[30] ),
    .Y(_09338_));
 sky130_fd_sc_hd__mux4_2 _13863_ (.A0(\w[1][0] ),
    .A1(\w[3][0] ),
    .A2(\w[5][0] ),
    .A3(\w[7][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02346_));
 sky130_fd_sc_hd__mux4_2 _13868_ (.A0(\w[9][0] ),
    .A1(\w[11][0] ),
    .A2(\w[13][0] ),
    .A3(\w[15][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02351_));
 sky130_fd_sc_hd__mux4_2 _13871_ (.A0(\w[17][0] ),
    .A1(\w[19][0] ),
    .A2(\w[21][0] ),
    .A3(\w[23][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02354_));
 sky130_fd_sc_hd__mux4_2 _13874_ (.A0(\w[25][0] ),
    .A1(\w[27][0] ),
    .A2(\w[29][0] ),
    .A3(\w[31][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02357_));
 sky130_fd_sc_hd__mux4_2 _13877_ (.A0(_02346_),
    .A1(_02351_),
    .A2(_02354_),
    .A3(_02357_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02360_));
 sky130_fd_sc_hd__mux4_2 _13880_ (.A0(\w[33][0] ),
    .A1(\w[35][0] ),
    .A2(\w[37][0] ),
    .A3(\w[39][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02363_));
 sky130_fd_sc_hd__mux4_2 _13883_ (.A0(\w[41][0] ),
    .A1(\w[43][0] ),
    .A2(\w[45][0] ),
    .A3(\w[47][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02366_));
 sky130_fd_sc_hd__mux4_2 _13886_ (.A0(\w[49][0] ),
    .A1(\w[51][0] ),
    .A2(\w[53][0] ),
    .A3(\w[55][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02369_));
 sky130_fd_sc_hd__mux4_2 _13889_ (.A0(\w[57][0] ),
    .A1(\w[59][0] ),
    .A2(\w[61][0] ),
    .A3(\w[63][0] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02372_));
 sky130_fd_sc_hd__mux4_2 _13892_ (.A0(_02363_),
    .A1(_02366_),
    .A2(_02369_),
    .A3(_02372_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02375_));
 sky130_fd_sc_hd__mux2i_1 _13894_ (.A0(_02360_),
    .A1(_02375_),
    .S(\count16_2[5] ),
    .Y(_09072_));
 sky130_fd_sc_hd__mux4_2 _13895_ (.A0(\w[1][1] ),
    .A1(\w[3][1] ),
    .A2(\w[5][1] ),
    .A3(\w[7][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02377_));
 sky130_fd_sc_hd__mux4_2 _13896_ (.A0(\w[9][1] ),
    .A1(\w[11][1] ),
    .A2(\w[13][1] ),
    .A3(\w[15][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02378_));
 sky130_fd_sc_hd__mux4_2 _13898_ (.A0(\w[17][1] ),
    .A1(\w[19][1] ),
    .A2(\w[21][1] ),
    .A3(\w[23][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02380_));
 sky130_fd_sc_hd__mux4_2 _13899_ (.A0(\w[25][1] ),
    .A1(\w[27][1] ),
    .A2(\w[29][1] ),
    .A3(\w[31][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02381_));
 sky130_fd_sc_hd__mux4_2 _13900_ (.A0(_02377_),
    .A1(_02378_),
    .A2(_02380_),
    .A3(_02381_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02382_));
 sky130_fd_sc_hd__mux4_2 _13901_ (.A0(\w[33][1] ),
    .A1(\w[35][1] ),
    .A2(\w[37][1] ),
    .A3(\w[39][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02383_));
 sky130_fd_sc_hd__mux4_2 _13902_ (.A0(\w[41][1] ),
    .A1(\w[43][1] ),
    .A2(\w[45][1] ),
    .A3(\w[47][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02384_));
 sky130_fd_sc_hd__mux4_2 _13903_ (.A0(\w[49][1] ),
    .A1(\w[51][1] ),
    .A2(\w[53][1] ),
    .A3(\w[55][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02385_));
 sky130_fd_sc_hd__mux4_2 _13905_ (.A0(\w[57][1] ),
    .A1(\w[59][1] ),
    .A2(\w[61][1] ),
    .A3(\w[63][1] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02387_));
 sky130_fd_sc_hd__mux4_2 _13906_ (.A0(_02383_),
    .A1(_02384_),
    .A2(_02385_),
    .A3(_02387_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02388_));
 sky130_fd_sc_hd__mux2i_1 _13907_ (.A0(_02382_),
    .A1(_02388_),
    .S(\count16_2[5] ),
    .Y(_09077_));
 sky130_fd_sc_hd__mux4_2 _13908_ (.A0(\w[1][2] ),
    .A1(\w[3][2] ),
    .A2(\w[5][2] ),
    .A3(\w[7][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02389_));
 sky130_fd_sc_hd__mux4_2 _13909_ (.A0(\w[9][2] ),
    .A1(\w[11][2] ),
    .A2(\w[13][2] ),
    .A3(\w[15][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02390_));
 sky130_fd_sc_hd__mux4_2 _13911_ (.A0(\w[17][2] ),
    .A1(\w[19][2] ),
    .A2(\w[21][2] ),
    .A3(\w[23][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02392_));
 sky130_fd_sc_hd__mux4_2 _13912_ (.A0(\w[25][2] ),
    .A1(\w[27][2] ),
    .A2(\w[29][2] ),
    .A3(\w[31][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02393_));
 sky130_fd_sc_hd__mux4_2 _13913_ (.A0(_02389_),
    .A1(_02390_),
    .A2(_02392_),
    .A3(_02393_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02394_));
 sky130_fd_sc_hd__mux4_2 _13915_ (.A0(\w[33][2] ),
    .A1(\w[35][2] ),
    .A2(\w[37][2] ),
    .A3(\w[39][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02396_));
 sky130_fd_sc_hd__mux4_2 _13916_ (.A0(\w[41][2] ),
    .A1(\w[43][2] ),
    .A2(\w[45][2] ),
    .A3(\w[47][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02397_));
 sky130_fd_sc_hd__mux4_2 _13917_ (.A0(\w[49][2] ),
    .A1(\w[51][2] ),
    .A2(\w[53][2] ),
    .A3(\w[55][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02398_));
 sky130_fd_sc_hd__mux4_2 _13918_ (.A0(\w[57][2] ),
    .A1(\w[59][2] ),
    .A2(\w[61][2] ),
    .A3(\w[63][2] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02399_));
 sky130_fd_sc_hd__mux4_2 _13919_ (.A0(_02396_),
    .A1(_02397_),
    .A2(_02398_),
    .A3(_02399_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02400_));
 sky130_fd_sc_hd__mux2i_1 _13920_ (.A0(_02394_),
    .A1(_02400_),
    .S(\count16_2[5] ),
    .Y(_09086_));
 sky130_fd_sc_hd__mux4_2 _13921_ (.A0(\w[1][3] ),
    .A1(\w[3][3] ),
    .A2(\w[5][3] ),
    .A3(\w[7][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02401_));
 sky130_fd_sc_hd__mux4_2 _13922_ (.A0(\w[9][3] ),
    .A1(\w[11][3] ),
    .A2(\w[13][3] ),
    .A3(\w[15][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02402_));
 sky130_fd_sc_hd__mux4_2 _13923_ (.A0(\w[17][3] ),
    .A1(\w[19][3] ),
    .A2(\w[21][3] ),
    .A3(\w[23][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02403_));
 sky130_fd_sc_hd__mux4_2 _13924_ (.A0(\w[25][3] ),
    .A1(\w[27][3] ),
    .A2(\w[29][3] ),
    .A3(\w[31][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02404_));
 sky130_fd_sc_hd__mux4_2 _13925_ (.A0(_02401_),
    .A1(_02402_),
    .A2(_02403_),
    .A3(_02404_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02405_));
 sky130_fd_sc_hd__mux4_2 _13927_ (.A0(\w[33][3] ),
    .A1(\w[35][3] ),
    .A2(\w[37][3] ),
    .A3(\w[39][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02407_));
 sky130_fd_sc_hd__mux4_2 _13928_ (.A0(\w[41][3] ),
    .A1(\w[43][3] ),
    .A2(\w[45][3] ),
    .A3(\w[47][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02408_));
 sky130_fd_sc_hd__mux4_2 _13930_ (.A0(\w[49][3] ),
    .A1(\w[51][3] ),
    .A2(\w[53][3] ),
    .A3(\w[55][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02410_));
 sky130_fd_sc_hd__mux4_2 _13931_ (.A0(\w[57][3] ),
    .A1(\w[59][3] ),
    .A2(\w[61][3] ),
    .A3(\w[63][3] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_2 _13932_ (.A0(_02407_),
    .A1(_02408_),
    .A2(_02410_),
    .A3(_02411_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02412_));
 sky130_fd_sc_hd__mux2i_1 _13933_ (.A0(_02405_),
    .A1(_02412_),
    .S(\count16_2[5] ),
    .Y(_09098_));
 sky130_fd_sc_hd__mux4_2 _13934_ (.A0(\w[1][4] ),
    .A1(\w[3][4] ),
    .A2(\w[5][4] ),
    .A3(\w[7][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02413_));
 sky130_fd_sc_hd__mux4_2 _13936_ (.A0(\w[9][4] ),
    .A1(\w[11][4] ),
    .A2(\w[13][4] ),
    .A3(\w[15][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__mux4_2 _13937_ (.A0(\w[17][4] ),
    .A1(\w[19][4] ),
    .A2(\w[21][4] ),
    .A3(\w[23][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02416_));
 sky130_fd_sc_hd__mux4_2 _13938_ (.A0(\w[25][4] ),
    .A1(\w[27][4] ),
    .A2(\w[29][4] ),
    .A3(\w[31][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02417_));
 sky130_fd_sc_hd__mux4_2 _13939_ (.A0(_02413_),
    .A1(_02415_),
    .A2(_02416_),
    .A3(_02417_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02418_));
 sky130_fd_sc_hd__mux4_2 _13940_ (.A0(\w[33][4] ),
    .A1(\w[35][4] ),
    .A2(\w[37][4] ),
    .A3(\w[39][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02419_));
 sky130_fd_sc_hd__mux4_2 _13941_ (.A0(\w[41][4] ),
    .A1(\w[43][4] ),
    .A2(\w[45][4] ),
    .A3(\w[47][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02420_));
 sky130_fd_sc_hd__mux4_2 _13943_ (.A0(\w[49][4] ),
    .A1(\w[51][4] ),
    .A2(\w[53][4] ),
    .A3(\w[55][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02422_));
 sky130_fd_sc_hd__mux4_2 _13944_ (.A0(\w[57][4] ),
    .A1(\w[59][4] ),
    .A2(\w[61][4] ),
    .A3(\w[63][4] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux4_2 _13945_ (.A0(_02419_),
    .A1(_02420_),
    .A2(_02422_),
    .A3(_02423_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02424_));
 sky130_fd_sc_hd__mux2i_1 _13946_ (.A0(_02418_),
    .A1(_02424_),
    .S(\count16_2[5] ),
    .Y(_09107_));
 sky130_fd_sc_hd__mux4_2 _13947_ (.A0(\w[1][5] ),
    .A1(\w[3][5] ),
    .A2(\w[5][5] ),
    .A3(\w[7][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02425_));
 sky130_fd_sc_hd__mux4_2 _13949_ (.A0(\w[9][5] ),
    .A1(\w[11][5] ),
    .A2(\w[13][5] ),
    .A3(\w[15][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02427_));
 sky130_fd_sc_hd__mux4_2 _13950_ (.A0(\w[17][5] ),
    .A1(\w[19][5] ),
    .A2(\w[21][5] ),
    .A3(\w[23][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02428_));
 sky130_fd_sc_hd__mux4_2 _13951_ (.A0(\w[25][5] ),
    .A1(\w[27][5] ),
    .A2(\w[29][5] ),
    .A3(\w[31][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02429_));
 sky130_fd_sc_hd__mux4_2 _13952_ (.A0(_02425_),
    .A1(_02427_),
    .A2(_02428_),
    .A3(_02429_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02430_));
 sky130_fd_sc_hd__mux4_2 _13953_ (.A0(\w[33][5] ),
    .A1(\w[35][5] ),
    .A2(\w[37][5] ),
    .A3(\w[39][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02431_));
 sky130_fd_sc_hd__mux4_2 _13955_ (.A0(\w[41][5] ),
    .A1(\w[43][5] ),
    .A2(\w[45][5] ),
    .A3(\w[47][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02433_));
 sky130_fd_sc_hd__mux4_2 _13956_ (.A0(\w[49][5] ),
    .A1(\w[51][5] ),
    .A2(\w[53][5] ),
    .A3(\w[55][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02434_));
 sky130_fd_sc_hd__mux4_2 _13957_ (.A0(\w[57][5] ),
    .A1(\w[59][5] ),
    .A2(\w[61][5] ),
    .A3(\w[63][5] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux4_2 _13958_ (.A0(_02431_),
    .A1(_02433_),
    .A2(_02434_),
    .A3(_02435_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02436_));
 sky130_fd_sc_hd__mux2i_1 _13959_ (.A0(_02430_),
    .A1(_02436_),
    .S(\count16_2[5] ),
    .Y(_09116_));
 sky130_fd_sc_hd__mux4_2 _13960_ (.A0(\w[1][6] ),
    .A1(\w[3][6] ),
    .A2(\w[5][6] ),
    .A3(\w[7][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02437_));
 sky130_fd_sc_hd__mux4_2 _13961_ (.A0(\w[9][6] ),
    .A1(\w[11][6] ),
    .A2(\w[13][6] ),
    .A3(\w[15][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02438_));
 sky130_fd_sc_hd__mux4_2 _13962_ (.A0(\w[17][6] ),
    .A1(\w[19][6] ),
    .A2(\w[21][6] ),
    .A3(\w[23][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02439_));
 sky130_fd_sc_hd__mux4_2 _13963_ (.A0(\w[25][6] ),
    .A1(\w[27][6] ),
    .A2(\w[29][6] ),
    .A3(\w[31][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02440_));
 sky130_fd_sc_hd__mux4_2 _13964_ (.A0(_02437_),
    .A1(_02438_),
    .A2(_02439_),
    .A3(_02440_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02441_));
 sky130_fd_sc_hd__mux4_2 _13965_ (.A0(\w[33][6] ),
    .A1(\w[35][6] ),
    .A2(\w[37][6] ),
    .A3(\w[39][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02442_));
 sky130_fd_sc_hd__mux4_2 _13967_ (.A0(\w[41][6] ),
    .A1(\w[43][6] ),
    .A2(\w[45][6] ),
    .A3(\w[47][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02444_));
 sky130_fd_sc_hd__mux4_2 _13968_ (.A0(\w[49][6] ),
    .A1(\w[51][6] ),
    .A2(\w[53][6] ),
    .A3(\w[55][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02445_));
 sky130_fd_sc_hd__mux4_2 _13969_ (.A0(\w[57][6] ),
    .A1(\w[59][6] ),
    .A2(\w[61][6] ),
    .A3(\w[63][6] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02446_));
 sky130_fd_sc_hd__mux4_2 _13970_ (.A0(_02442_),
    .A1(_02444_),
    .A2(_02445_),
    .A3(_02446_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02447_));
 sky130_fd_sc_hd__mux2i_1 _13971_ (.A0(_02441_),
    .A1(_02447_),
    .S(\count16_2[5] ),
    .Y(_09125_));
 sky130_fd_sc_hd__mux4_2 _13972_ (.A0(\w[1][7] ),
    .A1(\w[3][7] ),
    .A2(\w[5][7] ),
    .A3(\w[7][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02448_));
 sky130_fd_sc_hd__mux4_2 _13973_ (.A0(\w[9][7] ),
    .A1(\w[11][7] ),
    .A2(\w[13][7] ),
    .A3(\w[15][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02449_));
 sky130_fd_sc_hd__mux4_2 _13974_ (.A0(\w[17][7] ),
    .A1(\w[19][7] ),
    .A2(\w[21][7] ),
    .A3(\w[23][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02450_));
 sky130_fd_sc_hd__mux4_2 _13975_ (.A0(\w[25][7] ),
    .A1(\w[27][7] ),
    .A2(\w[29][7] ),
    .A3(\w[31][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02451_));
 sky130_fd_sc_hd__mux4_2 _13977_ (.A0(_02448_),
    .A1(_02449_),
    .A2(_02450_),
    .A3(_02451_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02453_));
 sky130_fd_sc_hd__mux4_2 _13978_ (.A0(\w[33][7] ),
    .A1(\w[35][7] ),
    .A2(\w[37][7] ),
    .A3(\w[39][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02454_));
 sky130_fd_sc_hd__mux4_2 _13979_ (.A0(\w[41][7] ),
    .A1(\w[43][7] ),
    .A2(\w[45][7] ),
    .A3(\w[47][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02455_));
 sky130_fd_sc_hd__mux4_2 _13980_ (.A0(\w[49][7] ),
    .A1(\w[51][7] ),
    .A2(\w[53][7] ),
    .A3(\w[55][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02456_));
 sky130_fd_sc_hd__mux4_2 _13981_ (.A0(\w[57][7] ),
    .A1(\w[59][7] ),
    .A2(\w[61][7] ),
    .A3(\w[63][7] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02457_));
 sky130_fd_sc_hd__mux4_2 _13982_ (.A0(_02454_),
    .A1(_02455_),
    .A2(_02456_),
    .A3(_02457_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02458_));
 sky130_fd_sc_hd__mux2i_1 _13983_ (.A0(_02453_),
    .A1(_02458_),
    .S(\count16_2[5] ),
    .Y(_09134_));
 sky130_fd_sc_hd__mux4_2 _13984_ (.A0(\w[1][8] ),
    .A1(\w[3][8] ),
    .A2(\w[5][8] ),
    .A3(\w[7][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02459_));
 sky130_fd_sc_hd__mux4_2 _13985_ (.A0(\w[9][8] ),
    .A1(\w[11][8] ),
    .A2(\w[13][8] ),
    .A3(\w[15][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02460_));
 sky130_fd_sc_hd__mux4_2 _13986_ (.A0(\w[17][8] ),
    .A1(\w[19][8] ),
    .A2(\w[21][8] ),
    .A3(\w[23][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02461_));
 sky130_fd_sc_hd__mux4_2 _13988_ (.A0(\w[25][8] ),
    .A1(\w[27][8] ),
    .A2(\w[29][8] ),
    .A3(\w[31][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02463_));
 sky130_fd_sc_hd__mux4_2 _13990_ (.A0(_02459_),
    .A1(_02460_),
    .A2(_02461_),
    .A3(_02463_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02465_));
 sky130_fd_sc_hd__mux4_2 _13991_ (.A0(\w[33][8] ),
    .A1(\w[35][8] ),
    .A2(\w[37][8] ),
    .A3(\w[39][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02466_));
 sky130_fd_sc_hd__mux4_2 _13992_ (.A0(\w[41][8] ),
    .A1(\w[43][8] ),
    .A2(\w[45][8] ),
    .A3(\w[47][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02467_));
 sky130_fd_sc_hd__mux4_2 _13993_ (.A0(\w[49][8] ),
    .A1(\w[51][8] ),
    .A2(\w[53][8] ),
    .A3(\w[55][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02468_));
 sky130_fd_sc_hd__mux4_2 _13994_ (.A0(\w[57][8] ),
    .A1(\w[59][8] ),
    .A2(\w[61][8] ),
    .A3(\w[63][8] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02469_));
 sky130_fd_sc_hd__mux4_2 _13996_ (.A0(_02466_),
    .A1(_02467_),
    .A2(_02468_),
    .A3(_02469_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02471_));
 sky130_fd_sc_hd__mux2i_1 _13997_ (.A0(_02465_),
    .A1(_02471_),
    .S(\count16_2[5] ),
    .Y(_09143_));
 sky130_fd_sc_hd__mux4_2 _13999_ (.A0(\w[1][9] ),
    .A1(\w[3][9] ),
    .A2(\w[5][9] ),
    .A3(\w[7][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02473_));
 sky130_fd_sc_hd__mux4_2 _14000_ (.A0(\w[9][9] ),
    .A1(\w[11][9] ),
    .A2(\w[13][9] ),
    .A3(\w[15][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02474_));
 sky130_fd_sc_hd__mux4_2 _14001_ (.A0(\w[17][9] ),
    .A1(\w[19][9] ),
    .A2(\w[21][9] ),
    .A3(\w[23][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02475_));
 sky130_fd_sc_hd__mux4_2 _14003_ (.A0(\w[25][9] ),
    .A1(\w[27][9] ),
    .A2(\w[29][9] ),
    .A3(\w[31][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02477_));
 sky130_fd_sc_hd__mux4_2 _14004_ (.A0(_02473_),
    .A1(_02474_),
    .A2(_02475_),
    .A3(_02477_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02478_));
 sky130_fd_sc_hd__mux4_2 _14005_ (.A0(\w[33][9] ),
    .A1(\w[35][9] ),
    .A2(\w[37][9] ),
    .A3(\w[39][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02479_));
 sky130_fd_sc_hd__mux4_2 _14006_ (.A0(\w[41][9] ),
    .A1(\w[43][9] ),
    .A2(\w[45][9] ),
    .A3(\w[47][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02480_));
 sky130_fd_sc_hd__mux4_2 _14007_ (.A0(\w[49][9] ),
    .A1(\w[51][9] ),
    .A2(\w[53][9] ),
    .A3(\w[55][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02481_));
 sky130_fd_sc_hd__mux4_2 _14008_ (.A0(\w[57][9] ),
    .A1(\w[59][9] ),
    .A2(\w[61][9] ),
    .A3(\w[63][9] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02482_));
 sky130_fd_sc_hd__mux4_2 _14010_ (.A0(_02479_),
    .A1(_02480_),
    .A2(_02481_),
    .A3(_02482_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02484_));
 sky130_fd_sc_hd__mux2i_1 _14011_ (.A0(_02478_),
    .A1(_02484_),
    .S(\count16_2[5] ),
    .Y(_09152_));
 sky130_fd_sc_hd__mux4_2 _14013_ (.A0(\w[1][10] ),
    .A1(\w[3][10] ),
    .A2(\w[5][10] ),
    .A3(\w[7][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02486_));
 sky130_fd_sc_hd__mux4_2 _14014_ (.A0(\w[9][10] ),
    .A1(\w[11][10] ),
    .A2(\w[13][10] ),
    .A3(\w[15][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02487_));
 sky130_fd_sc_hd__mux4_2 _14015_ (.A0(\w[17][10] ),
    .A1(\w[19][10] ),
    .A2(\w[21][10] ),
    .A3(\w[23][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02488_));
 sky130_fd_sc_hd__mux4_2 _14016_ (.A0(\w[25][10] ),
    .A1(\w[27][10] ),
    .A2(\w[29][10] ),
    .A3(\w[31][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02489_));
 sky130_fd_sc_hd__mux4_2 _14017_ (.A0(_02486_),
    .A1(_02487_),
    .A2(_02488_),
    .A3(_02489_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02490_));
 sky130_fd_sc_hd__mux4_2 _14018_ (.A0(\w[33][10] ),
    .A1(\w[35][10] ),
    .A2(\w[37][10] ),
    .A3(\w[39][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02491_));
 sky130_fd_sc_hd__mux4_2 _14019_ (.A0(\w[41][10] ),
    .A1(\w[43][10] ),
    .A2(\w[45][10] ),
    .A3(\w[47][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02492_));
 sky130_fd_sc_hd__mux4_2 _14020_ (.A0(\w[49][10] ),
    .A1(\w[51][10] ),
    .A2(\w[53][10] ),
    .A3(\w[55][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02493_));
 sky130_fd_sc_hd__mux4_2 _14022_ (.A0(\w[57][10] ),
    .A1(\w[59][10] ),
    .A2(\w[61][10] ),
    .A3(\w[63][10] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02495_));
 sky130_fd_sc_hd__mux4_2 _14023_ (.A0(_02491_),
    .A1(_02492_),
    .A2(_02493_),
    .A3(_02495_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02496_));
 sky130_fd_sc_hd__mux2i_1 _14025_ (.A0(_02490_),
    .A1(_02496_),
    .S(\count16_2[5] ),
    .Y(_09161_));
 sky130_fd_sc_hd__mux4_2 _14026_ (.A0(\w[1][11] ),
    .A1(\w[3][11] ),
    .A2(\w[5][11] ),
    .A3(\w[7][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02498_));
 sky130_fd_sc_hd__mux4_2 _14027_ (.A0(\w[9][11] ),
    .A1(\w[11][11] ),
    .A2(\w[13][11] ),
    .A3(\w[15][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02499_));
 sky130_fd_sc_hd__mux4_2 _14029_ (.A0(\w[17][11] ),
    .A1(\w[19][11] ),
    .A2(\w[21][11] ),
    .A3(\w[23][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02501_));
 sky130_fd_sc_hd__mux4_2 _14030_ (.A0(\w[25][11] ),
    .A1(\w[27][11] ),
    .A2(\w[29][11] ),
    .A3(\w[31][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02502_));
 sky130_fd_sc_hd__mux4_2 _14031_ (.A0(_02498_),
    .A1(_02499_),
    .A2(_02501_),
    .A3(_02502_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02503_));
 sky130_fd_sc_hd__mux4_2 _14032_ (.A0(\w[33][11] ),
    .A1(\w[35][11] ),
    .A2(\w[37][11] ),
    .A3(\w[39][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02504_));
 sky130_fd_sc_hd__mux4_2 _14033_ (.A0(\w[41][11] ),
    .A1(\w[43][11] ),
    .A2(\w[45][11] ),
    .A3(\w[47][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02505_));
 sky130_fd_sc_hd__mux4_2 _14034_ (.A0(\w[49][11] ),
    .A1(\w[51][11] ),
    .A2(\w[53][11] ),
    .A3(\w[55][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02506_));
 sky130_fd_sc_hd__mux4_2 _14036_ (.A0(\w[57][11] ),
    .A1(\w[59][11] ),
    .A2(\w[61][11] ),
    .A3(\w[63][11] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02508_));
 sky130_fd_sc_hd__mux4_2 _14037_ (.A0(_02504_),
    .A1(_02505_),
    .A2(_02506_),
    .A3(_02508_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02509_));
 sky130_fd_sc_hd__mux2i_1 _14038_ (.A0(_02503_),
    .A1(_02509_),
    .S(\count16_2[5] ),
    .Y(_09170_));
 sky130_fd_sc_hd__mux4_2 _14039_ (.A0(\w[1][12] ),
    .A1(\w[3][12] ),
    .A2(\w[5][12] ),
    .A3(\w[7][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02510_));
 sky130_fd_sc_hd__mux4_2 _14040_ (.A0(\w[9][12] ),
    .A1(\w[11][12] ),
    .A2(\w[13][12] ),
    .A3(\w[15][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02511_));
 sky130_fd_sc_hd__mux4_2 _14042_ (.A0(\w[17][12] ),
    .A1(\w[19][12] ),
    .A2(\w[21][12] ),
    .A3(\w[23][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02513_));
 sky130_fd_sc_hd__mux4_2 _14043_ (.A0(\w[25][12] ),
    .A1(\w[27][12] ),
    .A2(\w[29][12] ),
    .A3(\w[31][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02514_));
 sky130_fd_sc_hd__mux4_2 _14044_ (.A0(_02510_),
    .A1(_02511_),
    .A2(_02513_),
    .A3(_02514_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02515_));
 sky130_fd_sc_hd__mux4_2 _14046_ (.A0(\w[33][12] ),
    .A1(\w[35][12] ),
    .A2(\w[37][12] ),
    .A3(\w[39][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02517_));
 sky130_fd_sc_hd__mux4_2 _14047_ (.A0(\w[41][12] ),
    .A1(\w[43][12] ),
    .A2(\w[45][12] ),
    .A3(\w[47][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02518_));
 sky130_fd_sc_hd__mux4_2 _14048_ (.A0(\w[49][12] ),
    .A1(\w[51][12] ),
    .A2(\w[53][12] ),
    .A3(\w[55][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02519_));
 sky130_fd_sc_hd__mux4_2 _14049_ (.A0(\w[57][12] ),
    .A1(\w[59][12] ),
    .A2(\w[61][12] ),
    .A3(\w[63][12] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02520_));
 sky130_fd_sc_hd__mux4_2 _14050_ (.A0(_02517_),
    .A1(_02518_),
    .A2(_02519_),
    .A3(_02520_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02521_));
 sky130_fd_sc_hd__mux2i_1 _14051_ (.A0(_02515_),
    .A1(_02521_),
    .S(\count16_2[5] ),
    .Y(_09179_));
 sky130_fd_sc_hd__mux4_2 _14052_ (.A0(\w[1][13] ),
    .A1(\w[3][13] ),
    .A2(\w[5][13] ),
    .A3(\w[7][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02522_));
 sky130_fd_sc_hd__mux4_2 _14053_ (.A0(\w[9][13] ),
    .A1(\w[11][13] ),
    .A2(\w[13][13] ),
    .A3(\w[15][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02523_));
 sky130_fd_sc_hd__mux4_2 _14054_ (.A0(\w[17][13] ),
    .A1(\w[19][13] ),
    .A2(\w[21][13] ),
    .A3(\w[23][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02524_));
 sky130_fd_sc_hd__mux4_2 _14055_ (.A0(\w[25][13] ),
    .A1(\w[27][13] ),
    .A2(\w[29][13] ),
    .A3(\w[31][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02525_));
 sky130_fd_sc_hd__mux4_2 _14056_ (.A0(_02522_),
    .A1(_02523_),
    .A2(_02524_),
    .A3(_02525_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02526_));
 sky130_fd_sc_hd__mux4_2 _14058_ (.A0(\w[33][13] ),
    .A1(\w[35][13] ),
    .A2(\w[37][13] ),
    .A3(\w[39][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02528_));
 sky130_fd_sc_hd__mux4_2 _14059_ (.A0(\w[41][13] ),
    .A1(\w[43][13] ),
    .A2(\w[45][13] ),
    .A3(\w[47][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02529_));
 sky130_fd_sc_hd__mux4_2 _14061_ (.A0(\w[49][13] ),
    .A1(\w[51][13] ),
    .A2(\w[53][13] ),
    .A3(\w[55][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02531_));
 sky130_fd_sc_hd__mux4_2 _14062_ (.A0(\w[57][13] ),
    .A1(\w[59][13] ),
    .A2(\w[61][13] ),
    .A3(\w[63][13] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02532_));
 sky130_fd_sc_hd__mux4_2 _14063_ (.A0(_02528_),
    .A1(_02529_),
    .A2(_02531_),
    .A3(_02532_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02533_));
 sky130_fd_sc_hd__mux2i_1 _14064_ (.A0(_02526_),
    .A1(_02533_),
    .S(\count16_2[5] ),
    .Y(_09188_));
 sky130_fd_sc_hd__mux4_2 _14065_ (.A0(\w[1][14] ),
    .A1(\w[3][14] ),
    .A2(\w[5][14] ),
    .A3(\w[7][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02534_));
 sky130_fd_sc_hd__mux4_2 _14067_ (.A0(\w[9][14] ),
    .A1(\w[11][14] ),
    .A2(\w[13][14] ),
    .A3(\w[15][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02536_));
 sky130_fd_sc_hd__mux4_2 _14068_ (.A0(\w[17][14] ),
    .A1(\w[19][14] ),
    .A2(\w[21][14] ),
    .A3(\w[23][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02537_));
 sky130_fd_sc_hd__mux4_2 _14069_ (.A0(\w[25][14] ),
    .A1(\w[27][14] ),
    .A2(\w[29][14] ),
    .A3(\w[31][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02538_));
 sky130_fd_sc_hd__mux4_2 _14070_ (.A0(_02534_),
    .A1(_02536_),
    .A2(_02537_),
    .A3(_02538_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02539_));
 sky130_fd_sc_hd__mux4_2 _14071_ (.A0(\w[33][14] ),
    .A1(\w[35][14] ),
    .A2(\w[37][14] ),
    .A3(\w[39][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02540_));
 sky130_fd_sc_hd__mux4_2 _14072_ (.A0(\w[41][14] ),
    .A1(\w[43][14] ),
    .A2(\w[45][14] ),
    .A3(\w[47][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02541_));
 sky130_fd_sc_hd__mux4_2 _14074_ (.A0(\w[49][14] ),
    .A1(\w[51][14] ),
    .A2(\w[53][14] ),
    .A3(\w[55][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02543_));
 sky130_fd_sc_hd__mux4_2 _14075_ (.A0(\w[57][14] ),
    .A1(\w[59][14] ),
    .A2(\w[61][14] ),
    .A3(\w[63][14] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02544_));
 sky130_fd_sc_hd__mux4_2 _14076_ (.A0(_02540_),
    .A1(_02541_),
    .A2(_02543_),
    .A3(_02544_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02545_));
 sky130_fd_sc_hd__mux2i_1 _14077_ (.A0(_02539_),
    .A1(_02545_),
    .S(\count16_2[5] ),
    .Y(_09197_));
 sky130_fd_sc_hd__mux4_2 _14078_ (.A0(\w[1][15] ),
    .A1(\w[3][15] ),
    .A2(\w[5][15] ),
    .A3(\w[7][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02546_));
 sky130_fd_sc_hd__mux4_2 _14080_ (.A0(\w[9][15] ),
    .A1(\w[11][15] ),
    .A2(\w[13][15] ),
    .A3(\w[15][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02548_));
 sky130_fd_sc_hd__mux4_2 _14081_ (.A0(\w[17][15] ),
    .A1(\w[19][15] ),
    .A2(\w[21][15] ),
    .A3(\w[23][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02549_));
 sky130_fd_sc_hd__mux4_2 _14082_ (.A0(\w[25][15] ),
    .A1(\w[27][15] ),
    .A2(\w[29][15] ),
    .A3(\w[31][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02550_));
 sky130_fd_sc_hd__mux4_2 _14083_ (.A0(_02546_),
    .A1(_02548_),
    .A2(_02549_),
    .A3(_02550_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02551_));
 sky130_fd_sc_hd__mux4_2 _14084_ (.A0(\w[33][15] ),
    .A1(\w[35][15] ),
    .A2(\w[37][15] ),
    .A3(\w[39][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02552_));
 sky130_fd_sc_hd__mux4_2 _14086_ (.A0(\w[41][15] ),
    .A1(\w[43][15] ),
    .A2(\w[45][15] ),
    .A3(\w[47][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02554_));
 sky130_fd_sc_hd__mux4_2 _14087_ (.A0(\w[49][15] ),
    .A1(\w[51][15] ),
    .A2(\w[53][15] ),
    .A3(\w[55][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02555_));
 sky130_fd_sc_hd__mux4_2 _14088_ (.A0(\w[57][15] ),
    .A1(\w[59][15] ),
    .A2(\w[61][15] ),
    .A3(\w[63][15] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02556_));
 sky130_fd_sc_hd__mux4_2 _14089_ (.A0(_02552_),
    .A1(_02554_),
    .A2(_02555_),
    .A3(_02556_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02557_));
 sky130_fd_sc_hd__mux2i_1 _14090_ (.A0(_02551_),
    .A1(_02557_),
    .S(\count16_2[5] ),
    .Y(_09206_));
 sky130_fd_sc_hd__mux4_2 _14091_ (.A0(\w[1][16] ),
    .A1(\w[3][16] ),
    .A2(\w[5][16] ),
    .A3(\w[7][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02558_));
 sky130_fd_sc_hd__mux4_2 _14092_ (.A0(\w[9][16] ),
    .A1(\w[11][16] ),
    .A2(\w[13][16] ),
    .A3(\w[15][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02559_));
 sky130_fd_sc_hd__mux4_2 _14093_ (.A0(\w[17][16] ),
    .A1(\w[19][16] ),
    .A2(\w[21][16] ),
    .A3(\w[23][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02560_));
 sky130_fd_sc_hd__mux4_2 _14094_ (.A0(\w[25][16] ),
    .A1(\w[27][16] ),
    .A2(\w[29][16] ),
    .A3(\w[31][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02561_));
 sky130_fd_sc_hd__mux4_2 _14095_ (.A0(_02558_),
    .A1(_02559_),
    .A2(_02560_),
    .A3(_02561_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02562_));
 sky130_fd_sc_hd__mux4_2 _14096_ (.A0(\w[33][16] ),
    .A1(\w[35][16] ),
    .A2(\w[37][16] ),
    .A3(\w[39][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02563_));
 sky130_fd_sc_hd__mux4_2 _14098_ (.A0(\w[41][16] ),
    .A1(\w[43][16] ),
    .A2(\w[45][16] ),
    .A3(\w[47][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02565_));
 sky130_fd_sc_hd__mux4_2 _14099_ (.A0(\w[49][16] ),
    .A1(\w[51][16] ),
    .A2(\w[53][16] ),
    .A3(\w[55][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02566_));
 sky130_fd_sc_hd__mux4_2 _14100_ (.A0(\w[57][16] ),
    .A1(\w[59][16] ),
    .A2(\w[61][16] ),
    .A3(\w[63][16] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02567_));
 sky130_fd_sc_hd__mux4_2 _14101_ (.A0(_02563_),
    .A1(_02565_),
    .A2(_02566_),
    .A3(_02567_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02568_));
 sky130_fd_sc_hd__mux2i_1 _14102_ (.A0(_02562_),
    .A1(_02568_),
    .S(\count16_2[5] ),
    .Y(_09215_));
 sky130_fd_sc_hd__mux4_2 _14103_ (.A0(\w[1][17] ),
    .A1(\w[3][17] ),
    .A2(\w[5][17] ),
    .A3(\w[7][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02569_));
 sky130_fd_sc_hd__mux4_2 _14104_ (.A0(\w[9][17] ),
    .A1(\w[11][17] ),
    .A2(\w[13][17] ),
    .A3(\w[15][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02570_));
 sky130_fd_sc_hd__mux4_2 _14105_ (.A0(\w[17][17] ),
    .A1(\w[19][17] ),
    .A2(\w[21][17] ),
    .A3(\w[23][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02571_));
 sky130_fd_sc_hd__mux4_2 _14106_ (.A0(\w[25][17] ),
    .A1(\w[27][17] ),
    .A2(\w[29][17] ),
    .A3(\w[31][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02572_));
 sky130_fd_sc_hd__mux4_2 _14108_ (.A0(_02569_),
    .A1(_02570_),
    .A2(_02571_),
    .A3(_02572_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02574_));
 sky130_fd_sc_hd__mux4_2 _14109_ (.A0(\w[33][17] ),
    .A1(\w[35][17] ),
    .A2(\w[37][17] ),
    .A3(\w[39][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02575_));
 sky130_fd_sc_hd__mux4_2 _14110_ (.A0(\w[41][17] ),
    .A1(\w[43][17] ),
    .A2(\w[45][17] ),
    .A3(\w[47][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02576_));
 sky130_fd_sc_hd__mux4_2 _14111_ (.A0(\w[49][17] ),
    .A1(\w[51][17] ),
    .A2(\w[53][17] ),
    .A3(\w[55][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02577_));
 sky130_fd_sc_hd__mux4_2 _14112_ (.A0(\w[57][17] ),
    .A1(\w[59][17] ),
    .A2(\w[61][17] ),
    .A3(\w[63][17] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02578_));
 sky130_fd_sc_hd__mux4_2 _14113_ (.A0(_02575_),
    .A1(_02576_),
    .A2(_02577_),
    .A3(_02578_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02579_));
 sky130_fd_sc_hd__mux2i_1 _14114_ (.A0(_02574_),
    .A1(_02579_),
    .S(\count16_2[5] ),
    .Y(_09224_));
 sky130_fd_sc_hd__mux4_2 _14115_ (.A0(\w[1][18] ),
    .A1(\w[3][18] ),
    .A2(\w[5][18] ),
    .A3(\w[7][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02580_));
 sky130_fd_sc_hd__mux4_2 _14116_ (.A0(\w[9][18] ),
    .A1(\w[11][18] ),
    .A2(\w[13][18] ),
    .A3(\w[15][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02581_));
 sky130_fd_sc_hd__mux4_2 _14117_ (.A0(\w[17][18] ),
    .A1(\w[19][18] ),
    .A2(\w[21][18] ),
    .A3(\w[23][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02582_));
 sky130_fd_sc_hd__mux4_2 _14119_ (.A0(\w[25][18] ),
    .A1(\w[27][18] ),
    .A2(\w[29][18] ),
    .A3(\w[31][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02584_));
 sky130_fd_sc_hd__mux4_2 _14121_ (.A0(_02580_),
    .A1(_02581_),
    .A2(_02582_),
    .A3(_02584_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02586_));
 sky130_fd_sc_hd__mux4_2 _14122_ (.A0(\w[33][18] ),
    .A1(\w[35][18] ),
    .A2(\w[37][18] ),
    .A3(\w[39][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02587_));
 sky130_fd_sc_hd__mux4_2 _14123_ (.A0(\w[41][18] ),
    .A1(\w[43][18] ),
    .A2(\w[45][18] ),
    .A3(\w[47][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02588_));
 sky130_fd_sc_hd__mux4_2 _14124_ (.A0(\w[49][18] ),
    .A1(\w[51][18] ),
    .A2(\w[53][18] ),
    .A3(\w[55][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02589_));
 sky130_fd_sc_hd__mux4_2 _14125_ (.A0(\w[57][18] ),
    .A1(\w[59][18] ),
    .A2(\w[61][18] ),
    .A3(\w[63][18] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02590_));
 sky130_fd_sc_hd__mux4_2 _14127_ (.A0(_02587_),
    .A1(_02588_),
    .A2(_02589_),
    .A3(_02590_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02592_));
 sky130_fd_sc_hd__mux2i_1 _14128_ (.A0(_02586_),
    .A1(_02592_),
    .S(\count16_2[5] ),
    .Y(_09233_));
 sky130_fd_sc_hd__mux4_2 _14130_ (.A0(\w[1][19] ),
    .A1(\w[3][19] ),
    .A2(\w[5][19] ),
    .A3(\w[7][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02594_));
 sky130_fd_sc_hd__mux4_2 _14131_ (.A0(\w[9][19] ),
    .A1(\w[11][19] ),
    .A2(\w[13][19] ),
    .A3(\w[15][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02595_));
 sky130_fd_sc_hd__mux4_2 _14132_ (.A0(\w[17][19] ),
    .A1(\w[19][19] ),
    .A2(\w[21][19] ),
    .A3(\w[23][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02596_));
 sky130_fd_sc_hd__mux4_2 _14134_ (.A0(\w[25][19] ),
    .A1(\w[27][19] ),
    .A2(\w[29][19] ),
    .A3(\w[31][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02598_));
 sky130_fd_sc_hd__mux4_2 _14135_ (.A0(_02594_),
    .A1(_02595_),
    .A2(_02596_),
    .A3(_02598_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02599_));
 sky130_fd_sc_hd__mux4_2 _14136_ (.A0(\w[33][19] ),
    .A1(\w[35][19] ),
    .A2(\w[37][19] ),
    .A3(\w[39][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02600_));
 sky130_fd_sc_hd__mux4_2 _14137_ (.A0(\w[41][19] ),
    .A1(\w[43][19] ),
    .A2(\w[45][19] ),
    .A3(\w[47][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02601_));
 sky130_fd_sc_hd__mux4_2 _14138_ (.A0(\w[49][19] ),
    .A1(\w[51][19] ),
    .A2(\w[53][19] ),
    .A3(\w[55][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02602_));
 sky130_fd_sc_hd__mux4_2 _14139_ (.A0(\w[57][19] ),
    .A1(\w[59][19] ),
    .A2(\w[61][19] ),
    .A3(\w[63][19] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02603_));
 sky130_fd_sc_hd__mux4_2 _14141_ (.A0(_02600_),
    .A1(_02601_),
    .A2(_02602_),
    .A3(_02603_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02605_));
 sky130_fd_sc_hd__mux2i_1 _14142_ (.A0(_02599_),
    .A1(_02605_),
    .S(\count16_2[5] ),
    .Y(_09242_));
 sky130_fd_sc_hd__mux4_2 _14143_ (.A0(\w[1][20] ),
    .A1(\w[3][20] ),
    .A2(\w[5][20] ),
    .A3(\w[7][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02606_));
 sky130_fd_sc_hd__mux4_2 _14144_ (.A0(\w[9][20] ),
    .A1(\w[11][20] ),
    .A2(\w[13][20] ),
    .A3(\w[15][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02607_));
 sky130_fd_sc_hd__mux4_2 _14145_ (.A0(\w[17][20] ),
    .A1(\w[19][20] ),
    .A2(\w[21][20] ),
    .A3(\w[23][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02608_));
 sky130_fd_sc_hd__mux4_2 _14146_ (.A0(\w[25][20] ),
    .A1(\w[27][20] ),
    .A2(\w[29][20] ),
    .A3(\w[31][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02609_));
 sky130_fd_sc_hd__mux4_2 _14147_ (.A0(_02606_),
    .A1(_02607_),
    .A2(_02608_),
    .A3(_02609_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02610_));
 sky130_fd_sc_hd__mux4_2 _14148_ (.A0(\w[33][20] ),
    .A1(\w[35][20] ),
    .A2(\w[37][20] ),
    .A3(\w[39][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02611_));
 sky130_fd_sc_hd__mux4_2 _14149_ (.A0(\w[41][20] ),
    .A1(\w[43][20] ),
    .A2(\w[45][20] ),
    .A3(\w[47][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02612_));
 sky130_fd_sc_hd__mux4_2 _14150_ (.A0(\w[49][20] ),
    .A1(\w[51][20] ),
    .A2(\w[53][20] ),
    .A3(\w[55][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02613_));
 sky130_fd_sc_hd__mux4_2 _14151_ (.A0(\w[57][20] ),
    .A1(\w[59][20] ),
    .A2(\w[61][20] ),
    .A3(\w[63][20] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02614_));
 sky130_fd_sc_hd__mux4_2 _14152_ (.A0(_02611_),
    .A1(_02612_),
    .A2(_02613_),
    .A3(_02614_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02615_));
 sky130_fd_sc_hd__mux2i_1 _14154_ (.A0(_02610_),
    .A1(_02615_),
    .S(\count16_2[5] ),
    .Y(_09251_));
 sky130_fd_sc_hd__mux4_2 _14155_ (.A0(\w[1][21] ),
    .A1(\w[3][21] ),
    .A2(\w[5][21] ),
    .A3(\w[7][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02617_));
 sky130_fd_sc_hd__mux4_2 _14156_ (.A0(\w[9][21] ),
    .A1(\w[11][21] ),
    .A2(\w[13][21] ),
    .A3(\w[15][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02618_));
 sky130_fd_sc_hd__mux4_2 _14157_ (.A0(\w[17][21] ),
    .A1(\w[19][21] ),
    .A2(\w[21][21] ),
    .A3(\w[23][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02619_));
 sky130_fd_sc_hd__mux4_2 _14158_ (.A0(\w[25][21] ),
    .A1(\w[27][21] ),
    .A2(\w[29][21] ),
    .A3(\w[31][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02620_));
 sky130_fd_sc_hd__mux4_2 _14159_ (.A0(_02617_),
    .A1(_02618_),
    .A2(_02619_),
    .A3(_02620_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02621_));
 sky130_fd_sc_hd__mux4_2 _14160_ (.A0(\w[33][21] ),
    .A1(\w[35][21] ),
    .A2(\w[37][21] ),
    .A3(\w[39][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02622_));
 sky130_fd_sc_hd__mux4_2 _14161_ (.A0(\w[41][21] ),
    .A1(\w[43][21] ),
    .A2(\w[45][21] ),
    .A3(\w[47][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02623_));
 sky130_fd_sc_hd__mux4_2 _14162_ (.A0(\w[49][21] ),
    .A1(\w[51][21] ),
    .A2(\w[53][21] ),
    .A3(\w[55][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02624_));
 sky130_fd_sc_hd__mux4_2 _14163_ (.A0(\w[57][21] ),
    .A1(\w[59][21] ),
    .A2(\w[61][21] ),
    .A3(\w[63][21] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02625_));
 sky130_fd_sc_hd__mux4_2 _14164_ (.A0(_02622_),
    .A1(_02623_),
    .A2(_02624_),
    .A3(_02625_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02626_));
 sky130_fd_sc_hd__mux2i_1 _14165_ (.A0(_02621_),
    .A1(_02626_),
    .S(\count16_2[5] ),
    .Y(_09260_));
 sky130_fd_sc_hd__mux4_2 _14166_ (.A0(\w[1][22] ),
    .A1(\w[3][22] ),
    .A2(\w[5][22] ),
    .A3(\w[7][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02627_));
 sky130_fd_sc_hd__mux4_2 _14167_ (.A0(\w[9][22] ),
    .A1(\w[11][22] ),
    .A2(\w[13][22] ),
    .A3(\w[15][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02628_));
 sky130_fd_sc_hd__mux4_2 _14168_ (.A0(\w[17][22] ),
    .A1(\w[19][22] ),
    .A2(\w[21][22] ),
    .A3(\w[23][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02629_));
 sky130_fd_sc_hd__mux4_2 _14169_ (.A0(\w[25][22] ),
    .A1(\w[27][22] ),
    .A2(\w[29][22] ),
    .A3(\w[31][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02630_));
 sky130_fd_sc_hd__mux4_2 _14170_ (.A0(_02627_),
    .A1(_02628_),
    .A2(_02629_),
    .A3(_02630_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02631_));
 sky130_fd_sc_hd__mux4_2 _14171_ (.A0(\w[33][22] ),
    .A1(\w[35][22] ),
    .A2(\w[37][22] ),
    .A3(\w[39][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02632_));
 sky130_fd_sc_hd__mux4_2 _14172_ (.A0(\w[41][22] ),
    .A1(\w[43][22] ),
    .A2(\w[45][22] ),
    .A3(\w[47][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02633_));
 sky130_fd_sc_hd__mux4_2 _14173_ (.A0(\w[49][22] ),
    .A1(\w[51][22] ),
    .A2(\w[53][22] ),
    .A3(\w[55][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02634_));
 sky130_fd_sc_hd__mux4_2 _14174_ (.A0(\w[57][22] ),
    .A1(\w[59][22] ),
    .A2(\w[61][22] ),
    .A3(\w[63][22] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02635_));
 sky130_fd_sc_hd__mux4_2 _14175_ (.A0(_02632_),
    .A1(_02633_),
    .A2(_02634_),
    .A3(_02635_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02636_));
 sky130_fd_sc_hd__mux2i_1 _14176_ (.A0(_02631_),
    .A1(_02636_),
    .S(\count16_2[5] ),
    .Y(_09269_));
 sky130_fd_sc_hd__mux4_2 _14177_ (.A0(\w[1][23] ),
    .A1(\w[3][23] ),
    .A2(\w[5][23] ),
    .A3(\w[7][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02637_));
 sky130_fd_sc_hd__mux4_2 _14178_ (.A0(\w[9][23] ),
    .A1(\w[11][23] ),
    .A2(\w[13][23] ),
    .A3(\w[15][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02638_));
 sky130_fd_sc_hd__mux4_2 _14179_ (.A0(\w[17][23] ),
    .A1(\w[19][23] ),
    .A2(\w[21][23] ),
    .A3(\w[23][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02639_));
 sky130_fd_sc_hd__mux4_2 _14180_ (.A0(\w[25][23] ),
    .A1(\w[27][23] ),
    .A2(\w[29][23] ),
    .A3(\w[31][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02640_));
 sky130_fd_sc_hd__mux4_2 _14181_ (.A0(_02637_),
    .A1(_02638_),
    .A2(_02639_),
    .A3(_02640_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02641_));
 sky130_fd_sc_hd__mux4_2 _14182_ (.A0(\w[33][23] ),
    .A1(\w[35][23] ),
    .A2(\w[37][23] ),
    .A3(\w[39][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02642_));
 sky130_fd_sc_hd__mux4_2 _14183_ (.A0(\w[41][23] ),
    .A1(\w[43][23] ),
    .A2(\w[45][23] ),
    .A3(\w[47][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02643_));
 sky130_fd_sc_hd__mux4_2 _14184_ (.A0(\w[49][23] ),
    .A1(\w[51][23] ),
    .A2(\w[53][23] ),
    .A3(\w[55][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02644_));
 sky130_fd_sc_hd__mux4_2 _14185_ (.A0(\w[57][23] ),
    .A1(\w[59][23] ),
    .A2(\w[61][23] ),
    .A3(\w[63][23] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02645_));
 sky130_fd_sc_hd__mux4_2 _14186_ (.A0(_02642_),
    .A1(_02643_),
    .A2(_02644_),
    .A3(_02645_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02646_));
 sky130_fd_sc_hd__mux2i_1 _14187_ (.A0(_02641_),
    .A1(_02646_),
    .S(\count16_2[5] ),
    .Y(_09278_));
 sky130_fd_sc_hd__mux4_2 _14188_ (.A0(\w[1][24] ),
    .A1(\w[3][24] ),
    .A2(\w[5][24] ),
    .A3(\w[7][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02647_));
 sky130_fd_sc_hd__mux4_2 _14189_ (.A0(\w[9][24] ),
    .A1(\w[11][24] ),
    .A2(\w[13][24] ),
    .A3(\w[15][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02648_));
 sky130_fd_sc_hd__mux4_2 _14190_ (.A0(\w[17][24] ),
    .A1(\w[19][24] ),
    .A2(\w[21][24] ),
    .A3(\w[23][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02649_));
 sky130_fd_sc_hd__mux4_2 _14191_ (.A0(\w[25][24] ),
    .A1(\w[27][24] ),
    .A2(\w[29][24] ),
    .A3(\w[31][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02650_));
 sky130_fd_sc_hd__mux4_2 _14192_ (.A0(_02647_),
    .A1(_02648_),
    .A2(_02649_),
    .A3(_02650_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02651_));
 sky130_fd_sc_hd__mux4_2 _14193_ (.A0(\w[33][24] ),
    .A1(\w[35][24] ),
    .A2(\w[37][24] ),
    .A3(\w[39][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02652_));
 sky130_fd_sc_hd__mux4_2 _14194_ (.A0(\w[41][24] ),
    .A1(\w[43][24] ),
    .A2(\w[45][24] ),
    .A3(\w[47][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02653_));
 sky130_fd_sc_hd__mux4_2 _14195_ (.A0(\w[49][24] ),
    .A1(\w[51][24] ),
    .A2(\w[53][24] ),
    .A3(\w[55][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02654_));
 sky130_fd_sc_hd__mux4_2 _14196_ (.A0(\w[57][24] ),
    .A1(\w[59][24] ),
    .A2(\w[61][24] ),
    .A3(\w[63][24] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02655_));
 sky130_fd_sc_hd__mux4_2 _14197_ (.A0(_02652_),
    .A1(_02653_),
    .A2(_02654_),
    .A3(_02655_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02656_));
 sky130_fd_sc_hd__mux2i_1 _14198_ (.A0(_02651_),
    .A1(_02656_),
    .S(\count16_2[5] ),
    .Y(_09287_));
 sky130_fd_sc_hd__mux4_2 _14199_ (.A0(\w[1][25] ),
    .A1(\w[3][25] ),
    .A2(\w[5][25] ),
    .A3(\w[7][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02657_));
 sky130_fd_sc_hd__mux4_2 _14200_ (.A0(\w[9][25] ),
    .A1(\w[11][25] ),
    .A2(\w[13][25] ),
    .A3(\w[15][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02658_));
 sky130_fd_sc_hd__mux4_2 _14201_ (.A0(\w[17][25] ),
    .A1(\w[19][25] ),
    .A2(\w[21][25] ),
    .A3(\w[23][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02659_));
 sky130_fd_sc_hd__mux4_2 _14202_ (.A0(\w[25][25] ),
    .A1(\w[27][25] ),
    .A2(\w[29][25] ),
    .A3(\w[31][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02660_));
 sky130_fd_sc_hd__mux4_2 _14203_ (.A0(_02657_),
    .A1(_02658_),
    .A2(_02659_),
    .A3(_02660_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02661_));
 sky130_fd_sc_hd__mux4_2 _14204_ (.A0(\w[33][25] ),
    .A1(\w[35][25] ),
    .A2(\w[37][25] ),
    .A3(\w[39][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02662_));
 sky130_fd_sc_hd__mux4_2 _14205_ (.A0(\w[41][25] ),
    .A1(\w[43][25] ),
    .A2(\w[45][25] ),
    .A3(\w[47][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02663_));
 sky130_fd_sc_hd__mux4_2 _14206_ (.A0(\w[49][25] ),
    .A1(\w[51][25] ),
    .A2(\w[53][25] ),
    .A3(\w[55][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02664_));
 sky130_fd_sc_hd__mux4_2 _14207_ (.A0(\w[57][25] ),
    .A1(\w[59][25] ),
    .A2(\w[61][25] ),
    .A3(\w[63][25] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02665_));
 sky130_fd_sc_hd__mux4_2 _14208_ (.A0(_02662_),
    .A1(_02663_),
    .A2(_02664_),
    .A3(_02665_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02666_));
 sky130_fd_sc_hd__mux2i_1 _14209_ (.A0(_02661_),
    .A1(_02666_),
    .S(\count16_2[5] ),
    .Y(_09296_));
 sky130_fd_sc_hd__mux4_2 _14210_ (.A0(\w[1][26] ),
    .A1(\w[3][26] ),
    .A2(\w[5][26] ),
    .A3(\w[7][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02667_));
 sky130_fd_sc_hd__mux4_2 _14211_ (.A0(\w[9][26] ),
    .A1(\w[11][26] ),
    .A2(\w[13][26] ),
    .A3(\w[15][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02668_));
 sky130_fd_sc_hd__mux4_2 _14212_ (.A0(\w[17][26] ),
    .A1(\w[19][26] ),
    .A2(\w[21][26] ),
    .A3(\w[23][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02669_));
 sky130_fd_sc_hd__mux4_2 _14213_ (.A0(\w[25][26] ),
    .A1(\w[27][26] ),
    .A2(\w[29][26] ),
    .A3(\w[31][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02670_));
 sky130_fd_sc_hd__mux4_2 _14214_ (.A0(_02667_),
    .A1(_02668_),
    .A2(_02669_),
    .A3(_02670_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02671_));
 sky130_fd_sc_hd__mux4_2 _14215_ (.A0(\w[33][26] ),
    .A1(\w[35][26] ),
    .A2(\w[37][26] ),
    .A3(\w[39][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02672_));
 sky130_fd_sc_hd__mux4_2 _14216_ (.A0(\w[41][26] ),
    .A1(\w[43][26] ),
    .A2(\w[45][26] ),
    .A3(\w[47][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02673_));
 sky130_fd_sc_hd__mux4_2 _14217_ (.A0(\w[49][26] ),
    .A1(\w[51][26] ),
    .A2(\w[53][26] ),
    .A3(\w[55][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02674_));
 sky130_fd_sc_hd__mux4_2 _14218_ (.A0(\w[57][26] ),
    .A1(\w[59][26] ),
    .A2(\w[61][26] ),
    .A3(\w[63][26] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02675_));
 sky130_fd_sc_hd__mux4_2 _14219_ (.A0(_02672_),
    .A1(_02673_),
    .A2(_02674_),
    .A3(_02675_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02676_));
 sky130_fd_sc_hd__mux2i_1 _14220_ (.A0(_02671_),
    .A1(_02676_),
    .S(\count16_2[5] ),
    .Y(_09305_));
 sky130_fd_sc_hd__mux4_2 _14221_ (.A0(\w[1][27] ),
    .A1(\w[3][27] ),
    .A2(\w[5][27] ),
    .A3(\w[7][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02677_));
 sky130_fd_sc_hd__mux4_2 _14222_ (.A0(\w[9][27] ),
    .A1(\w[11][27] ),
    .A2(\w[13][27] ),
    .A3(\w[15][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02678_));
 sky130_fd_sc_hd__mux4_2 _14223_ (.A0(\w[17][27] ),
    .A1(\w[19][27] ),
    .A2(\w[21][27] ),
    .A3(\w[23][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02679_));
 sky130_fd_sc_hd__mux4_2 _14224_ (.A0(\w[25][27] ),
    .A1(\w[27][27] ),
    .A2(\w[29][27] ),
    .A3(\w[31][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02680_));
 sky130_fd_sc_hd__mux4_2 _14225_ (.A0(_02677_),
    .A1(_02678_),
    .A2(_02679_),
    .A3(_02680_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02681_));
 sky130_fd_sc_hd__mux4_2 _14226_ (.A0(\w[33][27] ),
    .A1(\w[35][27] ),
    .A2(\w[37][27] ),
    .A3(\w[39][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02682_));
 sky130_fd_sc_hd__mux4_2 _14227_ (.A0(\w[41][27] ),
    .A1(\w[43][27] ),
    .A2(\w[45][27] ),
    .A3(\w[47][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02683_));
 sky130_fd_sc_hd__mux4_2 _14228_ (.A0(\w[49][27] ),
    .A1(\w[51][27] ),
    .A2(\w[53][27] ),
    .A3(\w[55][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02684_));
 sky130_fd_sc_hd__mux4_2 _14229_ (.A0(\w[57][27] ),
    .A1(\w[59][27] ),
    .A2(\w[61][27] ),
    .A3(\w[63][27] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02685_));
 sky130_fd_sc_hd__mux4_2 _14230_ (.A0(_02682_),
    .A1(_02683_),
    .A2(_02684_),
    .A3(_02685_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02686_));
 sky130_fd_sc_hd__mux2i_1 _14231_ (.A0(_02681_),
    .A1(_02686_),
    .S(\count16_2[5] ),
    .Y(_09314_));
 sky130_fd_sc_hd__inv_1 _14232_ (.A(_09324_),
    .Y(_09326_));
 sky130_fd_sc_hd__inv_1 _14233_ (.A(_09332_),
    .Y(_09335_));
 sky130_fd_sc_hd__mux4_2 _14234_ (.A0(\w[1][30] ),
    .A1(\w[3][30] ),
    .A2(\w[5][30] ),
    .A3(\w[7][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02687_));
 sky130_fd_sc_hd__mux4_2 _14235_ (.A0(\w[9][30] ),
    .A1(\w[11][30] ),
    .A2(\w[13][30] ),
    .A3(\w[15][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02688_));
 sky130_fd_sc_hd__mux4_2 _14236_ (.A0(\w[17][30] ),
    .A1(\w[19][30] ),
    .A2(\w[21][30] ),
    .A3(\w[23][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02689_));
 sky130_fd_sc_hd__mux4_2 _14237_ (.A0(\w[25][30] ),
    .A1(\w[27][30] ),
    .A2(\w[29][30] ),
    .A3(\w[31][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02690_));
 sky130_fd_sc_hd__mux4_2 _14238_ (.A0(_02687_),
    .A1(_02688_),
    .A2(_02689_),
    .A3(_02690_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02691_));
 sky130_fd_sc_hd__mux4_2 _14239_ (.A0(\w[33][30] ),
    .A1(\w[35][30] ),
    .A2(\w[37][30] ),
    .A3(\w[39][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02692_));
 sky130_fd_sc_hd__mux4_2 _14240_ (.A0(\w[41][30] ),
    .A1(\w[43][30] ),
    .A2(\w[45][30] ),
    .A3(\w[47][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02693_));
 sky130_fd_sc_hd__mux4_2 _14241_ (.A0(\w[49][30] ),
    .A1(\w[51][30] ),
    .A2(\w[53][30] ),
    .A3(\w[55][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02694_));
 sky130_fd_sc_hd__mux4_2 _14242_ (.A0(\w[57][30] ),
    .A1(\w[59][30] ),
    .A2(\w[61][30] ),
    .A3(\w[63][30] ),
    .S0(\count16_2[1] ),
    .S1(\count16_2[2] ),
    .X(_02695_));
 sky130_fd_sc_hd__mux4_2 _14243_ (.A0(_02692_),
    .A1(_02693_),
    .A2(_02694_),
    .A3(_02695_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_02696_));
 sky130_fd_sc_hd__mux2i_1 _14244_ (.A0(_02691_),
    .A1(_02696_),
    .S(\count16_2[5] ),
    .Y(_09340_));
 sky130_fd_sc_hd__inv_1 _14245_ (.A(_08827_),
    .Y(_08830_));
 sky130_fd_sc_hd__inv_1 _14246_ (.A(_08835_),
    .Y(_08838_));
 sky130_fd_sc_hd__inv_1 _14247_ (.A(_08848_),
    .Y(_08851_));
 sky130_fd_sc_hd__inv_1 _14248_ (.A(_08856_),
    .Y(_08859_));
 sky130_fd_sc_hd__inv_1 _14249_ (.A(_08864_),
    .Y(_08867_));
 sky130_fd_sc_hd__inv_1 _14250_ (.A(_08872_),
    .Y(_08875_));
 sky130_fd_sc_hd__inv_1 _14251_ (.A(_08880_),
    .Y(_08883_));
 sky130_fd_sc_hd__inv_1 _14252_ (.A(_08888_),
    .Y(_08891_));
 sky130_fd_sc_hd__inv_1 _14253_ (.A(_08896_),
    .Y(_08899_));
 sky130_fd_sc_hd__inv_1 _14254_ (.A(_08904_),
    .Y(_08907_));
 sky130_fd_sc_hd__inv_1 _14255_ (.A(_08912_),
    .Y(_08915_));
 sky130_fd_sc_hd__inv_1 _14256_ (.A(_08920_),
    .Y(_08923_));
 sky130_fd_sc_hd__inv_1 _14257_ (.A(_08928_),
    .Y(_08931_));
 sky130_fd_sc_hd__inv_1 _14258_ (.A(_08936_),
    .Y(_08939_));
 sky130_fd_sc_hd__inv_1 _14259_ (.A(_08944_),
    .Y(_08947_));
 sky130_fd_sc_hd__inv_1 _14260_ (.A(_08952_),
    .Y(_08955_));
 sky130_fd_sc_hd__inv_1 _14261_ (.A(_08960_),
    .Y(_08963_));
 sky130_fd_sc_hd__inv_1 _14262_ (.A(_08968_),
    .Y(_08971_));
 sky130_fd_sc_hd__inv_1 _14263_ (.A(_08976_),
    .Y(_08979_));
 sky130_fd_sc_hd__inv_1 _14264_ (.A(_08984_),
    .Y(_08987_));
 sky130_fd_sc_hd__inv_1 _14265_ (.A(_08992_),
    .Y(_08995_));
 sky130_fd_sc_hd__inv_1 _14266_ (.A(_09000_),
    .Y(_09003_));
 sky130_fd_sc_hd__inv_1 _14267_ (.A(_09008_),
    .Y(_09011_));
 sky130_fd_sc_hd__inv_1 _14268_ (.A(_09016_),
    .Y(_09019_));
 sky130_fd_sc_hd__inv_1 _14269_ (.A(_09024_),
    .Y(_09027_));
 sky130_fd_sc_hd__inv_1 _14270_ (.A(_09032_),
    .Y(_09035_));
 sky130_fd_sc_hd__inv_1 _14271_ (.A(_09040_),
    .Y(_09043_));
 sky130_fd_sc_hd__inv_1 _14272_ (.A(_09048_),
    .Y(_09051_));
 sky130_fd_sc_hd__inv_1 _14273_ (.A(_09056_),
    .Y(_09059_));
 sky130_fd_sc_hd__inv_1 _14274_ (.A(_09064_),
    .Y(_09067_));
 sky130_fd_sc_hd__inv_1 _14275_ (.A(_08823_),
    .Y(_08829_));
 sky130_fd_sc_hd__inv_1 _14276_ (.A(_08826_),
    .Y(_08837_));
 sky130_fd_sc_hd__inv_1 _14277_ (.A(_08834_),
    .Y(_08850_));
 sky130_fd_sc_hd__inv_1 _14278_ (.A(_08847_),
    .Y(_08858_));
 sky130_fd_sc_hd__inv_1 _14279_ (.A(_08855_),
    .Y(_08866_));
 sky130_fd_sc_hd__inv_1 _14280_ (.A(_08863_),
    .Y(_08874_));
 sky130_fd_sc_hd__inv_1 _14281_ (.A(_08871_),
    .Y(_08882_));
 sky130_fd_sc_hd__inv_1 _14282_ (.A(_08879_),
    .Y(_08890_));
 sky130_fd_sc_hd__inv_1 _14283_ (.A(_08887_),
    .Y(_08898_));
 sky130_fd_sc_hd__inv_1 _14284_ (.A(_08895_),
    .Y(_08906_));
 sky130_fd_sc_hd__inv_1 _14285_ (.A(_08903_),
    .Y(_08914_));
 sky130_fd_sc_hd__inv_1 _14286_ (.A(_08911_),
    .Y(_08922_));
 sky130_fd_sc_hd__inv_1 _14287_ (.A(_08919_),
    .Y(_08930_));
 sky130_fd_sc_hd__inv_1 _14288_ (.A(_08927_),
    .Y(_08938_));
 sky130_fd_sc_hd__inv_1 _14289_ (.A(_08935_),
    .Y(_08946_));
 sky130_fd_sc_hd__inv_1 _14290_ (.A(_08943_),
    .Y(_08954_));
 sky130_fd_sc_hd__inv_1 _14291_ (.A(_08951_),
    .Y(_08962_));
 sky130_fd_sc_hd__inv_1 _14292_ (.A(_08959_),
    .Y(_08970_));
 sky130_fd_sc_hd__inv_1 _14293_ (.A(_08967_),
    .Y(_08978_));
 sky130_fd_sc_hd__inv_1 _14294_ (.A(_08975_),
    .Y(_08986_));
 sky130_fd_sc_hd__inv_1 _14295_ (.A(_08983_),
    .Y(_08994_));
 sky130_fd_sc_hd__inv_1 _14296_ (.A(_08991_),
    .Y(_09002_));
 sky130_fd_sc_hd__inv_1 _14297_ (.A(_08999_),
    .Y(_09010_));
 sky130_fd_sc_hd__inv_1 _14298_ (.A(_09007_),
    .Y(_09018_));
 sky130_fd_sc_hd__inv_1 _14299_ (.A(_09015_),
    .Y(_09026_));
 sky130_fd_sc_hd__inv_1 _14300_ (.A(_09023_),
    .Y(_09034_));
 sky130_fd_sc_hd__inv_1 _14301_ (.A(_09031_),
    .Y(_09042_));
 sky130_fd_sc_hd__inv_1 _14302_ (.A(_09039_),
    .Y(_09050_));
 sky130_fd_sc_hd__inv_1 _14303_ (.A(_09047_),
    .Y(_09058_));
 sky130_fd_sc_hd__inv_1 _14304_ (.A(_09055_),
    .Y(_09066_));
 sky130_fd_sc_hd__inv_1 _14305_ (.A(_09323_),
    .Y(_09334_));
 sky130_fd_sc_hd__inv_1 _14306_ (.A(\count_hash2[1] ),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_4 _14307_ (.A(\count_hash1[1] ),
    .Y(_00654_));
 sky130_fd_sc_hd__mux4_2 _14308_ (.A0(\w[1][0] ),
    .A1(\w[3][0] ),
    .A2(\w[5][0] ),
    .A3(\w[7][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02697_));
 sky130_fd_sc_hd__mux4_2 _14309_ (.A0(\w[9][0] ),
    .A1(\w[11][0] ),
    .A2(\w[13][0] ),
    .A3(\w[15][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02698_));
 sky130_fd_sc_hd__mux4_2 _14310_ (.A0(\w[17][0] ),
    .A1(\w[19][0] ),
    .A2(\w[21][0] ),
    .A3(\w[23][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02699_));
 sky130_fd_sc_hd__mux4_2 _14311_ (.A0(\w[25][0] ),
    .A1(\w[27][0] ),
    .A2(\w[29][0] ),
    .A3(\w[31][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02700_));
 sky130_fd_sc_hd__mux4_2 _14312_ (.A0(_02697_),
    .A1(_02698_),
    .A2(_02699_),
    .A3(_02700_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_02701_));
 sky130_fd_sc_hd__mux4_2 _14313_ (.A0(\w[33][0] ),
    .A1(\w[35][0] ),
    .A2(\w[37][0] ),
    .A3(\w[39][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02702_));
 sky130_fd_sc_hd__mux4_2 _14314_ (.A0(\w[41][0] ),
    .A1(\w[43][0] ),
    .A2(\w[45][0] ),
    .A3(\w[47][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02703_));
 sky130_fd_sc_hd__mux4_2 _14315_ (.A0(\w[49][0] ),
    .A1(\w[51][0] ),
    .A2(\w[53][0] ),
    .A3(\w[55][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02704_));
 sky130_fd_sc_hd__mux4_2 _14316_ (.A0(\w[57][0] ),
    .A1(\w[59][0] ),
    .A2(\w[61][0] ),
    .A3(\w[63][0] ),
    .S0(\count7_1[1] ),
    .S1(\count7_1[2] ),
    .X(_02705_));
 sky130_fd_sc_hd__mux4_2 _14317_ (.A0(_02702_),
    .A1(_02703_),
    .A2(_02704_),
    .A3(_02705_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_2 _14318_ (.A0(_02701_),
    .A1(_02706_),
    .S(\count7_1[5] ),
    .X(_09368_));
 sky130_fd_sc_hd__inv_1 _14319_ (.A(_08831_),
    .Y(_08842_));
 sky130_fd_sc_hd__inv_1 _14320_ (.A(_08839_),
    .Y(_09375_));
 sky130_fd_sc_hd__inv_1 _14321_ (.A(_08852_),
    .Y(_09379_));
 sky130_fd_sc_hd__inv_1 _14322_ (.A(_08868_),
    .Y(_09383_));
 sky130_fd_sc_hd__inv_1 _14323_ (.A(_08860_),
    .Y(_09387_));
 sky130_fd_sc_hd__inv_1 _14324_ (.A(_08876_),
    .Y(_09391_));
 sky130_fd_sc_hd__inv_1 _14325_ (.A(_08884_),
    .Y(_09395_));
 sky130_fd_sc_hd__inv_1 _14326_ (.A(_08892_),
    .Y(_09399_));
 sky130_fd_sc_hd__inv_1 _14327_ (.A(_08900_),
    .Y(_09403_));
 sky130_fd_sc_hd__inv_1 _14328_ (.A(_08908_),
    .Y(_09407_));
 sky130_fd_sc_hd__inv_1 _14329_ (.A(_08916_),
    .Y(_09411_));
 sky130_fd_sc_hd__inv_1 _14330_ (.A(_08924_),
    .Y(_09415_));
 sky130_fd_sc_hd__inv_1 _14331_ (.A(_08932_),
    .Y(_09419_));
 sky130_fd_sc_hd__inv_1 _14332_ (.A(_08948_),
    .Y(_09423_));
 sky130_fd_sc_hd__inv_1 _14333_ (.A(_08940_),
    .Y(_09427_));
 sky130_fd_sc_hd__inv_1 _14334_ (.A(_08956_),
    .Y(_09431_));
 sky130_fd_sc_hd__inv_1 _14335_ (.A(_08964_),
    .Y(_09435_));
 sky130_fd_sc_hd__inv_1 _14336_ (.A(_08972_),
    .Y(_09439_));
 sky130_fd_sc_hd__inv_1 _14337_ (.A(_08980_),
    .Y(_09443_));
 sky130_fd_sc_hd__inv_1 _14338_ (.A(_08988_),
    .Y(_09447_));
 sky130_fd_sc_hd__inv_1 _14339_ (.A(_08996_),
    .Y(_09451_));
 sky130_fd_sc_hd__inv_1 _14340_ (.A(_09004_),
    .Y(_09455_));
 sky130_fd_sc_hd__inv_1 _14341_ (.A(_09012_),
    .Y(_09459_));
 sky130_fd_sc_hd__inv_1 _14342_ (.A(_09020_),
    .Y(_09463_));
 sky130_fd_sc_hd__inv_1 _14343_ (.A(_09028_),
    .Y(_09467_));
 sky130_fd_sc_hd__inv_1 _14344_ (.A(_09036_),
    .Y(_09471_));
 sky130_fd_sc_hd__inv_1 _14345_ (.A(_09044_),
    .Y(_09475_));
 sky130_fd_sc_hd__inv_1 _14346_ (.A(_09052_),
    .Y(_09479_));
 sky130_fd_sc_hd__inv_1 _14347_ (.A(_09060_),
    .Y(_09483_));
 sky130_fd_sc_hd__inv_1 _14348_ (.A(_09074_),
    .Y(_09487_));
 sky130_fd_sc_hd__inv_1 _14349_ (.A(_09073_),
    .Y(_09080_));
 sky130_fd_sc_hd__inv_1 _14350_ (.A(_09078_),
    .Y(_09089_));
 sky130_fd_sc_hd__inv_1 _14351_ (.A(_09087_),
    .Y(_09101_));
 sky130_fd_sc_hd__inv_1 _14352_ (.A(_09099_),
    .Y(_09110_));
 sky130_fd_sc_hd__inv_1 _14353_ (.A(_09108_),
    .Y(_09119_));
 sky130_fd_sc_hd__inv_1 _14354_ (.A(_09117_),
    .Y(_09128_));
 sky130_fd_sc_hd__inv_1 _14355_ (.A(_09126_),
    .Y(_09137_));
 sky130_fd_sc_hd__inv_1 _14356_ (.A(_09135_),
    .Y(_09146_));
 sky130_fd_sc_hd__inv_1 _14357_ (.A(_09144_),
    .Y(_09155_));
 sky130_fd_sc_hd__inv_1 _14358_ (.A(_09153_),
    .Y(_09164_));
 sky130_fd_sc_hd__inv_1 _14359_ (.A(_09162_),
    .Y(_09173_));
 sky130_fd_sc_hd__inv_1 _14360_ (.A(_09171_),
    .Y(_09182_));
 sky130_fd_sc_hd__inv_1 _14361_ (.A(_09180_),
    .Y(_09191_));
 sky130_fd_sc_hd__inv_1 _14362_ (.A(_09189_),
    .Y(_09200_));
 sky130_fd_sc_hd__inv_1 _14363_ (.A(_09198_),
    .Y(_09209_));
 sky130_fd_sc_hd__inv_1 _14364_ (.A(_09207_),
    .Y(_09218_));
 sky130_fd_sc_hd__inv_1 _14365_ (.A(_09216_),
    .Y(_09227_));
 sky130_fd_sc_hd__inv_1 _14366_ (.A(_09225_),
    .Y(_09236_));
 sky130_fd_sc_hd__inv_1 _14367_ (.A(_09234_),
    .Y(_09245_));
 sky130_fd_sc_hd__inv_1 _14368_ (.A(_09243_),
    .Y(_09254_));
 sky130_fd_sc_hd__inv_1 _14369_ (.A(_09252_),
    .Y(_09263_));
 sky130_fd_sc_hd__inv_1 _14370_ (.A(_09261_),
    .Y(_09272_));
 sky130_fd_sc_hd__inv_1 _14371_ (.A(_09270_),
    .Y(_09281_));
 sky130_fd_sc_hd__inv_1 _14372_ (.A(_09279_),
    .Y(_09290_));
 sky130_fd_sc_hd__inv_1 _14373_ (.A(_09288_),
    .Y(_09299_));
 sky130_fd_sc_hd__inv_1 _14374_ (.A(_09297_),
    .Y(_09308_));
 sky130_fd_sc_hd__inv_1 _14375_ (.A(_09306_),
    .Y(_09317_));
 sky130_fd_sc_hd__mux4_2 _14377_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02708_));
 sky130_fd_sc_hd__mux4_2 _14378_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02709_));
 sky130_fd_sc_hd__mux4_2 _14379_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02710_));
 sky130_fd_sc_hd__mux4_2 _14380_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02711_));
 sky130_fd_sc_hd__mux4_2 _14381_ (.A0(_02708_),
    .A1(_02709_),
    .A2(_02710_),
    .A3(_02711_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_02712_));
 sky130_fd_sc_hd__mux4_2 _14382_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02713_));
 sky130_fd_sc_hd__mux4_2 _14383_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02714_));
 sky130_fd_sc_hd__mux4_2 _14384_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02715_));
 sky130_fd_sc_hd__mux4_2 _14385_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02716_));
 sky130_fd_sc_hd__mux4_2 _14386_ (.A0(_02713_),
    .A1(_02714_),
    .A2(_02715_),
    .A3(_02716_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_02717_));
 sky130_fd_sc_hd__mux2_2 _14387_ (.A0(_02712_),
    .A1(_02717_),
    .S(\count7_2[5] ),
    .X(_09321_));
 sky130_fd_sc_hd__mux4_2 _14388_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02718_));
 sky130_fd_sc_hd__mux4_2 _14389_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02719_));
 sky130_fd_sc_hd__mux4_2 _14390_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02720_));
 sky130_fd_sc_hd__mux4_2 _14391_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02721_));
 sky130_fd_sc_hd__mux4_2 _14392_ (.A0(_02718_),
    .A1(_02719_),
    .A2(_02720_),
    .A3(_02721_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_02722_));
 sky130_fd_sc_hd__mux4_2 _14393_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02723_));
 sky130_fd_sc_hd__mux4_2 _14394_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02724_));
 sky130_fd_sc_hd__mux4_2 _14395_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02725_));
 sky130_fd_sc_hd__mux4_2 _14396_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_02726_));
 sky130_fd_sc_hd__mux4_2 _14397_ (.A0(_02723_),
    .A1(_02724_),
    .A2(_02725_),
    .A3(_02726_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_02727_));
 sky130_fd_sc_hd__mux2_2 _14398_ (.A0(_02722_),
    .A1(_02727_),
    .S(\count7_2[5] ),
    .X(_09329_));
 sky130_fd_sc_hd__inv_1 _14399_ (.A(_09327_),
    .Y(_09546_));
 sky130_fd_sc_hd__inv_1 _14400_ (.A(_09336_),
    .Y(_09550_));
 sky130_fd_sc_hd__inv_1 _14401_ (.A(\count_1[1] ),
    .Y(_00650_));
 sky130_fd_sc_hd__inv_1 _14402_ (.A(\count_2[1] ),
    .Y(_00652_));
 sky130_fd_sc_hd__inv_1 _14403_ (.A(\count_hash2[2] ),
    .Y(_09346_));
 sky130_fd_sc_hd__inv_1 _14404_ (.A(_08832_),
    .Y(_09371_));
 sky130_fd_sc_hd__inv_1 _14405_ (.A(_08840_),
    .Y(_08843_));
 sky130_fd_sc_hd__inv_1 _14406_ (.A(_08853_),
    .Y(_09376_));
 sky130_fd_sc_hd__inv_1 _14407_ (.A(_08861_),
    .Y(_09380_));
 sky130_fd_sc_hd__inv_1 _14408_ (.A(_08877_),
    .Y(_09384_));
 sky130_fd_sc_hd__inv_1 _14409_ (.A(_08869_),
    .Y(_09388_));
 sky130_fd_sc_hd__inv_1 _14410_ (.A(_08885_),
    .Y(_09392_));
 sky130_fd_sc_hd__inv_1 _14411_ (.A(_08893_),
    .Y(_09396_));
 sky130_fd_sc_hd__inv_1 _14412_ (.A(_08901_),
    .Y(_09400_));
 sky130_fd_sc_hd__inv_1 _14413_ (.A(_08909_),
    .Y(_09404_));
 sky130_fd_sc_hd__inv_1 _14414_ (.A(_08917_),
    .Y(_09408_));
 sky130_fd_sc_hd__inv_1 _14415_ (.A(_08925_),
    .Y(_09412_));
 sky130_fd_sc_hd__inv_1 _14416_ (.A(_08933_),
    .Y(_09416_));
 sky130_fd_sc_hd__inv_1 _14417_ (.A(_08941_),
    .Y(_09420_));
 sky130_fd_sc_hd__inv_1 _14418_ (.A(_08957_),
    .Y(_09424_));
 sky130_fd_sc_hd__inv_1 _14419_ (.A(_08949_),
    .Y(_09428_));
 sky130_fd_sc_hd__inv_1 _14420_ (.A(_08965_),
    .Y(_09432_));
 sky130_fd_sc_hd__inv_1 _14421_ (.A(_08973_),
    .Y(_09436_));
 sky130_fd_sc_hd__inv_1 _14422_ (.A(_08981_),
    .Y(_09440_));
 sky130_fd_sc_hd__inv_1 _14423_ (.A(_08989_),
    .Y(_09444_));
 sky130_fd_sc_hd__inv_1 _14424_ (.A(_08997_),
    .Y(_09448_));
 sky130_fd_sc_hd__inv_1 _14425_ (.A(_09005_),
    .Y(_09452_));
 sky130_fd_sc_hd__inv_1 _14426_ (.A(_09013_),
    .Y(_09456_));
 sky130_fd_sc_hd__inv_1 _14427_ (.A(_09021_),
    .Y(_09460_));
 sky130_fd_sc_hd__inv_1 _14428_ (.A(_09029_),
    .Y(_09464_));
 sky130_fd_sc_hd__inv_1 _14429_ (.A(_09037_),
    .Y(_09468_));
 sky130_fd_sc_hd__inv_1 _14430_ (.A(_09045_),
    .Y(_09472_));
 sky130_fd_sc_hd__inv_1 _14431_ (.A(_09053_),
    .Y(_09476_));
 sky130_fd_sc_hd__inv_1 _14432_ (.A(_09061_),
    .Y(_09480_));
 sky130_fd_sc_hd__inv_1 _14433_ (.A(_09069_),
    .Y(_09484_));
 sky130_fd_sc_hd__inv_1 _14434_ (.A(_09079_),
    .Y(_09081_));
 sky130_fd_sc_hd__inv_1 _14435_ (.A(_09088_),
    .Y(_09090_));
 sky130_fd_sc_hd__inv_1 _14436_ (.A(_09100_),
    .Y(_09102_));
 sky130_fd_sc_hd__inv_1 _14437_ (.A(_09109_),
    .Y(_09111_));
 sky130_fd_sc_hd__inv_1 _14438_ (.A(_09118_),
    .Y(_09120_));
 sky130_fd_sc_hd__inv_1 _14439_ (.A(_09127_),
    .Y(_09129_));
 sky130_fd_sc_hd__inv_1 _14440_ (.A(_09136_),
    .Y(_09138_));
 sky130_fd_sc_hd__inv_1 _14441_ (.A(_09145_),
    .Y(_09147_));
 sky130_fd_sc_hd__inv_1 _14442_ (.A(_09154_),
    .Y(_09156_));
 sky130_fd_sc_hd__inv_1 _14443_ (.A(_09163_),
    .Y(_09165_));
 sky130_fd_sc_hd__inv_1 _14444_ (.A(_09172_),
    .Y(_09174_));
 sky130_fd_sc_hd__inv_1 _14445_ (.A(_09181_),
    .Y(_09183_));
 sky130_fd_sc_hd__inv_1 _14446_ (.A(_09190_),
    .Y(_09192_));
 sky130_fd_sc_hd__inv_1 _14447_ (.A(_09199_),
    .Y(_09201_));
 sky130_fd_sc_hd__inv_1 _14448_ (.A(_09208_),
    .Y(_09210_));
 sky130_fd_sc_hd__inv_1 _14449_ (.A(_09217_),
    .Y(_09219_));
 sky130_fd_sc_hd__inv_1 _14450_ (.A(_09226_),
    .Y(_09228_));
 sky130_fd_sc_hd__inv_1 _14451_ (.A(_09235_),
    .Y(_09237_));
 sky130_fd_sc_hd__inv_1 _14452_ (.A(_09244_),
    .Y(_09246_));
 sky130_fd_sc_hd__inv_1 _14453_ (.A(_09253_),
    .Y(_09255_));
 sky130_fd_sc_hd__inv_1 _14454_ (.A(_09262_),
    .Y(_09264_));
 sky130_fd_sc_hd__inv_1 _14455_ (.A(_09271_),
    .Y(_09273_));
 sky130_fd_sc_hd__inv_1 _14456_ (.A(_09280_),
    .Y(_09282_));
 sky130_fd_sc_hd__inv_1 _14457_ (.A(_09289_),
    .Y(_09291_));
 sky130_fd_sc_hd__inv_1 _14458_ (.A(_09298_),
    .Y(_09300_));
 sky130_fd_sc_hd__inv_1 _14459_ (.A(_09307_),
    .Y(_09309_));
 sky130_fd_sc_hd__inv_1 _14460_ (.A(_09316_),
    .Y(_09318_));
 sky130_fd_sc_hd__inv_1 _14461_ (.A(_09328_),
    .Y(_09543_));
 sky130_fd_sc_hd__inv_1 _14462_ (.A(_09337_),
    .Y(_09547_));
 sky130_fd_sc_hd__inv_1 _14463_ (.A(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__inv_1 _14464_ (.A(\count_1[2] ),
    .Y(_09553_));
 sky130_fd_sc_hd__inv_1 _14465_ (.A(\count_2[2] ),
    .Y(_09561_));
 sky130_fd_sc_hd__nor2_1 _14470_ (.A(\count15_1[1] ),
    .B(reset),
    .Y(_00658_));
 sky130_fd_sc_hd__nor2b_1 _14472_ (.A(reset),
    .B_N(_00644_),
    .Y(_00659_));
 sky130_fd_sc_hd__xnor2_1 _14476_ (.A(\count15_1[3] ),
    .B(_09575_),
    .Y(_02736_));
 sky130_fd_sc_hd__nor2_1 _14477_ (.A(reset),
    .B(_02736_),
    .Y(_00660_));
 sky130_fd_sc_hd__nand3_2 _14483_ (.A(\count15_1[1] ),
    .B(\count15_1[2] ),
    .C(\count15_1[3] ),
    .Y(_02742_));
 sky130_fd_sc_hd__xor2_1 _14484_ (.A(\count15_1[4] ),
    .B(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__nor2_1 _14485_ (.A(reset),
    .B(_02743_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand3_1 _14487_ (.A(\count15_1[3] ),
    .B(\count15_1[4] ),
    .C(_09575_),
    .Y(_02745_));
 sky130_fd_sc_hd__xor2_1 _14488_ (.A(\count15_1[5] ),
    .B(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__nor2_1 _14489_ (.A(reset),
    .B(_02746_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _14493_ (.A(_05334_),
    .B(\count15_2[1] ),
    .Y(_00663_));
 sky130_fd_sc_hd__nor2b_1 _14494_ (.A(reset),
    .B_N(_00648_),
    .Y(_00664_));
 sky130_fd_sc_hd__xnor2_1 _14498_ (.A(\count15_2[3] ),
    .B(_09570_),
    .Y(_02753_));
 sky130_fd_sc_hd__nor2_1 _14499_ (.A(reset),
    .B(_02753_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand3_2 _14505_ (.A(\count15_2[1] ),
    .B(\count15_2[2] ),
    .C(\count15_2[3] ),
    .Y(_02759_));
 sky130_fd_sc_hd__xor2_1 _14506_ (.A(\count15_2[4] ),
    .B(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__nor2_1 _14507_ (.A(reset),
    .B(_02760_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand3_1 _14509_ (.A(\count15_2[3] ),
    .B(\count15_2[4] ),
    .C(_09570_),
    .Y(_02762_));
 sky130_fd_sc_hd__xor2_1 _14510_ (.A(\count15_2[5] ),
    .B(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__nor2_1 _14511_ (.A(reset),
    .B(_02763_),
    .Y(_00667_));
 sky130_fd_sc_hd__nor2_1 _14512_ (.A(\count16_1[1] ),
    .B(reset),
    .Y(_00668_));
 sky130_fd_sc_hd__nor2b_1 _14513_ (.A(reset),
    .B_N(_00645_),
    .Y(_00669_));
 sky130_fd_sc_hd__xnor2_1 _14514_ (.A(\count16_1[3] ),
    .B(_09574_),
    .Y(_02764_));
 sky130_fd_sc_hd__nor2_1 _14515_ (.A(reset),
    .B(_02764_),
    .Y(_00670_));
 sky130_fd_sc_hd__nand3_2 _14517_ (.A(\count16_1[1] ),
    .B(\count16_1[2] ),
    .C(\count16_1[3] ),
    .Y(_02766_));
 sky130_fd_sc_hd__xor2_1 _14518_ (.A(\count16_1[4] ),
    .B(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_1 _14519_ (.A(reset),
    .B(_02767_),
    .Y(_00671_));
 sky130_fd_sc_hd__nand3_1 _14520_ (.A(\count16_1[3] ),
    .B(\count16_1[4] ),
    .C(_09574_),
    .Y(_02768_));
 sky130_fd_sc_hd__xor2_1 _14521_ (.A(\count16_1[5] ),
    .B(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__nor2_1 _14522_ (.A(reset),
    .B(_02769_),
    .Y(_00672_));
 sky130_fd_sc_hd__nor2_1 _14523_ (.A(reset),
    .B(\count16_2[1] ),
    .Y(_00673_));
 sky130_fd_sc_hd__nor2b_1 _14524_ (.A(reset),
    .B_N(_00649_),
    .Y(_00674_));
 sky130_fd_sc_hd__xnor2_1 _14525_ (.A(\count16_2[3] ),
    .B(_09571_),
    .Y(_02770_));
 sky130_fd_sc_hd__nor2_1 _14526_ (.A(reset),
    .B(_02770_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand3_2 _14527_ (.A(\count16_2[1] ),
    .B(\count16_2[2] ),
    .C(\count16_2[3] ),
    .Y(_02771_));
 sky130_fd_sc_hd__xor2_1 _14528_ (.A(\count16_2[4] ),
    .B(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__nor2_1 _14529_ (.A(reset),
    .B(_02772_),
    .Y(_00676_));
 sky130_fd_sc_hd__nand3_1 _14530_ (.A(\count16_2[3] ),
    .B(\count16_2[4] ),
    .C(_09571_),
    .Y(_02773_));
 sky130_fd_sc_hd__xor2_1 _14531_ (.A(\count16_2[5] ),
    .B(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__nor2_1 _14532_ (.A(reset),
    .B(_02774_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _14536_ (.A(_05334_),
    .B(\count2_1[1] ),
    .Y(_00678_));
 sky130_fd_sc_hd__or2_2 _14537_ (.A(reset),
    .B(_00642_),
    .X(_00679_));
 sky130_fd_sc_hd__xnor2_1 _14541_ (.A(\count2_1[3] ),
    .B(_09569_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand2_1 _14542_ (.A(_05334_),
    .B(_02781_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand3_2 _14548_ (.A(\count2_1[1] ),
    .B(\count2_1[2] ),
    .C(\count2_1[3] ),
    .Y(_02787_));
 sky130_fd_sc_hd__xor2_1 _14549_ (.A(\count2_1[4] ),
    .B(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__nor2_1 _14550_ (.A(reset),
    .B(_02788_),
    .Y(_00681_));
 sky130_fd_sc_hd__nand3_1 _14552_ (.A(\count2_1[3] ),
    .B(\count2_1[4] ),
    .C(_09569_),
    .Y(_02790_));
 sky130_fd_sc_hd__xor2_1 _14553_ (.A(\count2_1[5] ),
    .B(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__nor2_1 _14554_ (.A(reset),
    .B(_02791_),
    .Y(_00682_));
 sky130_fd_sc_hd__nand2_1 _14558_ (.A(\count2_2[1] ),
    .B(_05334_),
    .Y(_00683_));
 sky130_fd_sc_hd__or2_2 _14559_ (.A(reset),
    .B(_00646_),
    .X(_00684_));
 sky130_fd_sc_hd__xnor2_1 _14563_ (.A(\count2_2[3] ),
    .B(_09573_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_1 _14564_ (.A(_05334_),
    .B(_02798_),
    .Y(_00685_));
 sky130_fd_sc_hd__nand3_2 _14570_ (.A(\count2_2[1] ),
    .B(\count2_2[2] ),
    .C(\count2_2[3] ),
    .Y(_02804_));
 sky130_fd_sc_hd__xor2_1 _14571_ (.A(\count2_2[4] ),
    .B(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__nor2_1 _14572_ (.A(reset),
    .B(_02805_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand3_1 _14574_ (.A(\count2_2[3] ),
    .B(\count2_2[4] ),
    .C(_09573_),
    .Y(_02807_));
 sky130_fd_sc_hd__xor2_1 _14575_ (.A(\count2_2[5] ),
    .B(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__nor2_1 _14576_ (.A(reset),
    .B(_02808_),
    .Y(_00687_));
 sky130_fd_sc_hd__nor2_1 _14577_ (.A(\count7_1[1] ),
    .B(reset),
    .Y(_00688_));
 sky130_fd_sc_hd__nor2b_1 _14578_ (.A(reset),
    .B_N(_00643_),
    .Y(_00689_));
 sky130_fd_sc_hd__xnor2_1 _14579_ (.A(\count7_1[3] ),
    .B(_09576_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2_1 _14580_ (.A(_05334_),
    .B(_02809_),
    .Y(_00690_));
 sky130_fd_sc_hd__nand3_2 _14582_ (.A(\count7_1[1] ),
    .B(\count7_1[2] ),
    .C(\count7_1[3] ),
    .Y(_02811_));
 sky130_fd_sc_hd__xor2_1 _14583_ (.A(\count7_1[4] ),
    .B(_02811_),
    .X(_02812_));
 sky130_fd_sc_hd__nor2_1 _14584_ (.A(reset),
    .B(_02812_),
    .Y(_00691_));
 sky130_fd_sc_hd__nand3_1 _14585_ (.A(\count7_1[3] ),
    .B(\count7_1[4] ),
    .C(_09576_),
    .Y(_02813_));
 sky130_fd_sc_hd__xor2_1 _14586_ (.A(\count7_1[5] ),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__nor2_1 _14587_ (.A(reset),
    .B(_02814_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _14588_ (.A(\count7_2[1] ),
    .B(_05334_),
    .Y(_00693_));
 sky130_fd_sc_hd__nor2b_1 _14589_ (.A(reset),
    .B_N(_00647_),
    .Y(_00694_));
 sky130_fd_sc_hd__xnor2_1 _14590_ (.A(\count7_2[3] ),
    .B(_09572_),
    .Y(_02815_));
 sky130_fd_sc_hd__nand2_1 _14591_ (.A(_05334_),
    .B(_02815_),
    .Y(_00695_));
 sky130_fd_sc_hd__nand3_2 _14592_ (.A(\count7_2[1] ),
    .B(\count7_2[2] ),
    .C(\count7_2[3] ),
    .Y(_02816_));
 sky130_fd_sc_hd__xor2_1 _14593_ (.A(\count7_2[4] ),
    .B(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__nor2_1 _14594_ (.A(reset),
    .B(_02817_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand3_1 _14595_ (.A(\count7_2[3] ),
    .B(\count7_2[4] ),
    .C(_09572_),
    .Y(_02818_));
 sky130_fd_sc_hd__xor2_1 _14596_ (.A(\count7_2[5] ),
    .B(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__nor2_1 _14597_ (.A(reset),
    .B(_02819_),
    .Y(_00697_));
 sky130_fd_sc_hd__xnor2_1 _14598_ (.A(_00650_),
    .B(_00128_),
    .Y(_02820_));
 sky130_fd_sc_hd__nor2_1 _14599_ (.A(reset),
    .B(_02820_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _14600_ (.A(\count_1[2] ),
    .B(_00128_),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_1 _14601_ (.A(_00651_),
    .B(_05331_),
    .Y(_02822_));
 sky130_fd_sc_hd__a21oi_1 _14602_ (.A1(_02821_),
    .A2(_02822_),
    .B1(reset),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _14603_ (.A(_09559_),
    .B(_05331_),
    .Y(_02823_));
 sky130_fd_sc_hd__xor2_1 _14604_ (.A(\count_1[3] ),
    .B(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__nor2_1 _14605_ (.A(reset),
    .B(_02824_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand4_1 _14606_ (.A(\count_1[3] ),
    .B(\count_1[2] ),
    .C(\count_1[1] ),
    .D(_05331_),
    .Y(_02825_));
 sky130_fd_sc_hd__xor2_1 _14607_ (.A(\count_1[4] ),
    .B(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__nand2_1 _14608_ (.A(_05334_),
    .B(_02826_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand4_1 _14609_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C(_09559_),
    .D(_05331_),
    .Y(_02827_));
 sky130_fd_sc_hd__xor2_1 _14610_ (.A(\count_1[5] ),
    .B(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__nor2_1 _14611_ (.A(reset),
    .B(_02828_),
    .Y(_00702_));
 sky130_fd_sc_hd__xnor2_1 _14612_ (.A(_00652_),
    .B(_00128_),
    .Y(_02829_));
 sky130_fd_sc_hd__nor2_1 _14613_ (.A(reset),
    .B(_02829_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_1 _14614_ (.A(\count_2[2] ),
    .B(_00128_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand2_1 _14615_ (.A(_00653_),
    .B(_05331_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21oi_1 _14616_ (.A1(_02830_),
    .A2(_02831_),
    .B1(reset),
    .Y(_00704_));
 sky130_fd_sc_hd__xnor2_1 _14617_ (.A(\count_2[3] ),
    .B(_09567_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21oi_1 _14618_ (.A1(_05331_),
    .A2(_02832_),
    .B1(reset),
    .Y(_00705_));
 sky130_fd_sc_hd__nand3_1 _14619_ (.A(\count_2[3] ),
    .B(\count_2[2] ),
    .C(\count_2[1] ),
    .Y(_02833_));
 sky130_fd_sc_hd__xor2_1 _14620_ (.A(\count_2[4] ),
    .B(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__nand3_1 _14621_ (.A(_05334_),
    .B(_05331_),
    .C(_02834_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand3_1 _14622_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_09567_),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_1 _14623_ (.A(\count_2[6] ),
    .B(\count_2[5] ),
    .Y(_02836_));
 sky130_fd_sc_hd__nor2_1 _14624_ (.A(_02835_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__a211oi_1 _14625_ (.A1(_05408_),
    .A2(_02835_),
    .B1(_02837_),
    .C1(reset),
    .Y(_00707_));
 sky130_fd_sc_hd__nor2b_1 _14626_ (.A(\count_2[6] ),
    .B_N(_05330_),
    .Y(_02838_));
 sky130_fd_sc_hd__nand2_1 _14627_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .Y(_02839_));
 sky130_fd_sc_hd__nor2_1 _14628_ (.A(_02833_),
    .B(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__mux2i_1 _14629_ (.A0(\count_2[6] ),
    .A1(_02838_),
    .S(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__nor2_1 _14630_ (.A(reset),
    .B(_02841_),
    .Y(_00708_));
 sky130_fd_sc_hd__nor2_1 _14633_ (.A(\count_hash1[6] ),
    .B(_05479_),
    .Y(_02844_));
 sky130_fd_sc_hd__nand2_1 _14634_ (.A(_09366_),
    .B(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__xnor2_1 _14635_ (.A(\count_hash1[1] ),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__nor2_1 _14636_ (.A(reset_hash),
    .B(_02846_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand3_1 _14637_ (.A(_09366_),
    .B(\count_hash1[2] ),
    .C(_02844_),
    .Y(_02847_));
 sky130_fd_sc_hd__nand2_1 _14638_ (.A(_00655_),
    .B(_02845_),
    .Y(_02848_));
 sky130_fd_sc_hd__a21oi_1 _14639_ (.A1(_02847_),
    .A2(_02848_),
    .B1(reset_hash),
    .Y(_00710_));
 sky130_fd_sc_hd__nor2_1 _14642_ (.A(_05953_),
    .B(_02844_),
    .Y(_02851_));
 sky130_fd_sc_hd__nor2_1 _14643_ (.A(reset_hash),
    .B(_02851_),
    .Y(_00711_));
 sky130_fd_sc_hd__a21oi_1 _14645_ (.A1(_05958_),
    .A2(_02845_),
    .B1(reset_hash),
    .Y(_00712_));
 sky130_fd_sc_hd__xor2_2 _14646_ (.A(\count_hash1[5] ),
    .B(_05977_),
    .X(_02853_));
 sky130_fd_sc_hd__a21oi_1 _14650_ (.A1(_02853_),
    .A2(_02845_),
    .B1(reset_hash),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_2 _14651_ (.A(\count_hash1[2] ),
    .B(\count_hash1[1] ),
    .Y(_02857_));
 sky130_fd_sc_hd__o21ai_0 _14652_ (.A1(_05479_),
    .A2(_02857_),
    .B1(\count_hash1[6] ),
    .Y(_02858_));
 sky130_fd_sc_hd__nor2_1 _14653_ (.A(_09366_),
    .B(_02857_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_1 _14654_ (.A(_02844_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__a21oi_1 _14655_ (.A1(_02858_),
    .A2(_02860_),
    .B1(reset_hash),
    .Y(_00714_));
 sky130_fd_sc_hd__xnor2_1 _14656_ (.A(\count_hash2[1] ),
    .B(_02845_),
    .Y(_02861_));
 sky130_fd_sc_hd__nor2_1 _14657_ (.A(reset_hash),
    .B(_02861_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand3_1 _14658_ (.A(\count_hash2[2] ),
    .B(_09366_),
    .C(_02844_),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_1 _14659_ (.A(_00657_),
    .B(_02845_),
    .Y(_02863_));
 sky130_fd_sc_hd__a21oi_1 _14660_ (.A1(_02862_),
    .A2(_02863_),
    .B1(reset_hash),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2_1 _14661_ (.A(_09354_),
    .B(_02845_),
    .Y(_02864_));
 sky130_fd_sc_hd__xor2_1 _14662_ (.A(\count_hash2[3] ),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__nor2_1 _14663_ (.A(reset_hash),
    .B(_02865_),
    .Y(_00717_));
 sky130_fd_sc_hd__a21oi_1 _14664_ (.A1(_09366_),
    .A2(_02844_),
    .B1(_05460_),
    .Y(_02866_));
 sky130_fd_sc_hd__xnor2_1 _14665_ (.A(\count_hash2[4] ),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__nor2_1 _14666_ (.A(reset_hash),
    .B(_02867_),
    .Y(_00718_));
 sky130_fd_sc_hd__a21oi_1 _14667_ (.A1(_09366_),
    .A2(_02844_),
    .B1(_05471_),
    .Y(_02868_));
 sky130_fd_sc_hd__xnor2_1 _14668_ (.A(\count_hash2[5] ),
    .B(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__nor2_1 _14669_ (.A(reset_hash),
    .B(_02869_),
    .Y(_00719_));
 sky130_fd_sc_hd__or2_2 _14671_ (.A(_09358_),
    .B(_09362_),
    .X(_02871_));
 sky130_fd_sc_hd__and2_1 _14672_ (.A(\count_hash1[2] ),
    .B(\count_hash1[1] ),
    .X(_02872_));
 sky130_fd_sc_hd__nor2b_1 _14673_ (.A(\count_hash1[4] ),
    .B_N(\count_hash1[3] ),
    .Y(_02873_));
 sky130_fd_sc_hd__nand2_1 _14674_ (.A(\count_hash1[3] ),
    .B(_09366_),
    .Y(_02874_));
 sky130_fd_sc_hd__or2_2 _14675_ (.A(\count_hash1[3] ),
    .B(_09366_),
    .X(_02875_));
 sky130_fd_sc_hd__o21ai_0 _14676_ (.A1(_02872_),
    .A2(_02874_),
    .B1(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__a32oi_1 _14677_ (.A1(_09366_),
    .A2(_02872_),
    .A3(_02873_),
    .B1(_02876_),
    .B2(\count_hash1[4] ),
    .Y(_02877_));
 sky130_fd_sc_hd__nor2_1 _14679_ (.A(_02853_),
    .B(_02877_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_1 _14684_ (.A(_09358_),
    .B(_05978_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _14685_ (.A(_09362_),
    .B(_02853_),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_1 _14686_ (.A(_02884_),
    .B(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__nand2_1 _14687_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .Y(_02887_));
 sky130_fd_sc_hd__a21oi_1 _14688_ (.A1(_02857_),
    .A2(_05951_),
    .B1(_05952_),
    .Y(_02888_));
 sky130_fd_sc_hd__o32ai_1 _14689_ (.A1(_09366_),
    .A2(_02887_),
    .A3(_02857_),
    .B1(_02888_),
    .B2(\count_hash1[4] ),
    .Y(_02889_));
 sky130_fd_sc_hd__nor2_1 _14690_ (.A(_02853_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__a21oi_1 _14691_ (.A1(_02853_),
    .A2(_02877_),
    .B1(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__o21ai_0 _14692_ (.A1(_09364_),
    .A2(_02886_),
    .B1(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__a21boi_0 _14693_ (.A1(_02871_),
    .A2(_02879_),
    .B1_N(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__xnor2_1 _14694_ (.A(\count_hash1[4] ),
    .B(_05957_),
    .Y(_02894_));
 sky130_fd_sc_hd__nor2_1 _14695_ (.A(_02894_),
    .B(_05953_),
    .Y(_02895_));
 sky130_fd_sc_hd__nor2_1 _14701_ (.A(_09357_),
    .B(_09362_),
    .Y(_02901_));
 sky130_fd_sc_hd__nor2_1 _14702_ (.A(_05978_),
    .B(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__a21o_1 _14703_ (.A1(_09364_),
    .A2(_05978_),
    .B1(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__nand2_1 _14705_ (.A(_05958_),
    .B(_05978_),
    .Y(_02905_));
 sky130_fd_sc_hd__nand2_1 _14706_ (.A(_02894_),
    .B(_02853_),
    .Y(_02906_));
 sky130_fd_sc_hd__nand2_1 _14707_ (.A(_02905_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__nand2_1 _14708_ (.A(_09362_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand2_1 _14710_ (.A(_09358_),
    .B(_02905_),
    .Y(_02910_));
 sky130_fd_sc_hd__nor2_1 _14711_ (.A(_05951_),
    .B(_05952_),
    .Y(_02911_));
 sky130_fd_sc_hd__a21oi_1 _14714_ (.A1(_02908_),
    .A2(_02910_),
    .B1(_02911_),
    .Y(_02914_));
 sky130_fd_sc_hd__a21oi_1 _14715_ (.A1(_02895_),
    .A2(_02903_),
    .B1(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__or2_2 _14716_ (.A(\count_hash1[6] ),
    .B(_05480_),
    .X(_02916_));
 sky130_fd_sc_hd__nor2_1 _14718_ (.A(reset_hash),
    .B(_02916_),
    .Y(_02918_));
 sky130_fd_sc_hd__a2bb2oi_1 _14719_ (.A1_N(_05956_),
    .A2_N(_02888_),
    .B1(_02873_),
    .B2(_02859_),
    .Y(_02919_));
 sky130_fd_sc_hd__nor2_1 _14720_ (.A(_09358_),
    .B(_09362_),
    .Y(_02920_));
 sky130_fd_sc_hd__nor2_1 _14721_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__nor2_1 _14722_ (.A(_09357_),
    .B(_09364_),
    .Y(_02922_));
 sky130_fd_sc_hd__a21oi_1 _14723_ (.A1(_02920_),
    .A2(_02922_),
    .B1(_02877_),
    .Y(_02923_));
 sky130_fd_sc_hd__o21ai_0 _14724_ (.A1(_02921_),
    .A2(_02923_),
    .B1(_02853_),
    .Y(_02924_));
 sky130_fd_sc_hd__nor2_1 _14725_ (.A(_02853_),
    .B(_02919_),
    .Y(_02925_));
 sky130_fd_sc_hd__o21bai_1 _14726_ (.A1(_02853_),
    .A2(_02919_),
    .B1_N(_02889_),
    .Y(_02926_));
 sky130_fd_sc_hd__and2_1 _14727_ (.A(_09357_),
    .B(_02889_),
    .X(_02927_));
 sky130_fd_sc_hd__a221oi_1 _14728_ (.A1(_09358_),
    .A2(_02925_),
    .B1(_02926_),
    .B2(_09364_),
    .C1(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__nor2_1 _14729_ (.A(_09362_),
    .B(_09364_),
    .Y(_02929_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(_05958_),
    .B(_02911_),
    .Y(_02930_));
 sky130_fd_sc_hd__nor2_1 _14731_ (.A(_02929_),
    .B(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__nor2_1 _14732_ (.A(_09358_),
    .B(_09364_),
    .Y(_02932_));
 sky130_fd_sc_hd__nor2_1 _14733_ (.A(_02877_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _14734_ (.A(_09358_),
    .B(_05958_),
    .Y(_02934_));
 sky130_fd_sc_hd__a21oi_1 _14735_ (.A1(_09362_),
    .A2(_02894_),
    .B1(_09357_),
    .Y(_02935_));
 sky130_fd_sc_hd__a21oi_1 _14736_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_05953_),
    .Y(_02936_));
 sky130_fd_sc_hd__o31ai_1 _14737_ (.A1(_02931_),
    .A2(_02933_),
    .A3(_02936_),
    .B1(_05978_),
    .Y(_02937_));
 sky130_fd_sc_hd__or2_2 _14738_ (.A(_09357_),
    .B(_09362_),
    .X(_02938_));
 sky130_fd_sc_hd__nor2_1 _14739_ (.A(_09358_),
    .B(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__o22ai_1 _14740_ (.A1(_02919_),
    .A2(_02922_),
    .B1(_02930_),
    .B2(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__a222oi_1 _14741_ (.A1(_02871_),
    .A2(_02889_),
    .B1(_02925_),
    .B2(_02938_),
    .C1(_02940_),
    .C2(_02853_),
    .Y(_02941_));
 sky130_fd_sc_hd__nand4_1 _14742_ (.A(_02924_),
    .B(_02928_),
    .C(_02937_),
    .D(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2_1 _14743_ (.A(_02918_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__a21oi_1 _14745_ (.A1(_02893_),
    .A2(_02915_),
    .B1(_02943_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand2_1 _14749_ (.A(_09358_),
    .B(_02889_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_1 _14750_ (.A(_05958_),
    .B(_02853_),
    .Y(_02949_));
 sky130_fd_sc_hd__inv_1 _14751_ (.A(_09357_),
    .Y(_02950_));
 sky130_fd_sc_hd__nor2_1 _14753_ (.A(_02911_),
    .B(_02853_),
    .Y(_02952_));
 sky130_fd_sc_hd__nor2_1 _14754_ (.A(_02950_),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__o21ai_0 _14755_ (.A1(_05953_),
    .A2(_02949_),
    .B1(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__a32o_1 _14756_ (.A1(_09366_),
    .A2(_02872_),
    .A3(_02873_),
    .B1(_02876_),
    .B2(\count_hash1[4] ),
    .X(_02955_));
 sky130_fd_sc_hd__nor2_1 _14757_ (.A(_05958_),
    .B(_02853_),
    .Y(_02956_));
 sky130_fd_sc_hd__nor2_1 _14758_ (.A(_02911_),
    .B(_02949_),
    .Y(_02957_));
 sky130_fd_sc_hd__o31ai_1 _14760_ (.A1(_02955_),
    .A2(_02956_),
    .A3(_02957_),
    .B1(_09362_),
    .Y(_02959_));
 sky130_fd_sc_hd__a41o_1 _14761_ (.A1(_02942_),
    .A2(_02948_),
    .A3(_02954_),
    .A4(_02959_),
    .B1(_02916_),
    .X(_02960_));
 sky130_fd_sc_hd__nand2_1 _14762_ (.A(_05476_),
    .B(_02960_),
    .Y(_00721_));
 sky130_fd_sc_hd__o21a_1 _14763_ (.A1(_02877_),
    .A2(_02884_),
    .B1(_02942_),
    .X(_02961_));
 sky130_fd_sc_hd__nand2_1 _14765_ (.A(_02853_),
    .B(_02923_),
    .Y(_02963_));
 sky130_fd_sc_hd__o21ai_0 _14767_ (.A1(_02895_),
    .A2(_02952_),
    .B1(_09357_),
    .Y(_02965_));
 sky130_fd_sc_hd__a21oi_1 _14768_ (.A1(_05958_),
    .A2(_02932_),
    .B1(_02853_),
    .Y(_02966_));
 sky130_fd_sc_hd__nor2_1 _14770_ (.A(_09364_),
    .B(_02911_),
    .Y(_02968_));
 sky130_fd_sc_hd__nor2_1 _14771_ (.A(_02894_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__o22ai_1 _14772_ (.A1(_05953_),
    .A2(_02966_),
    .B1(_02969_),
    .B2(_09362_),
    .Y(_02970_));
 sky130_fd_sc_hd__nand4_1 _14773_ (.A(_02961_),
    .B(_02963_),
    .C(_02965_),
    .D(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__a21o_1 _14774_ (.A1(_05481_),
    .A2(_02971_),
    .B1(reset_hash),
    .X(_00722_));
 sky130_fd_sc_hd__and2_1 _14775_ (.A(_05978_),
    .B(_02889_),
    .X(_02972_));
 sky130_fd_sc_hd__nand2_1 _14776_ (.A(_09357_),
    .B(_02911_),
    .Y(_02973_));
 sky130_fd_sc_hd__nor2_1 _14777_ (.A(_05958_),
    .B(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_1 _14778_ (.A(_09362_),
    .B(_02889_),
    .Y(_02975_));
 sky130_fd_sc_hd__a21oi_1 _14779_ (.A1(_02973_),
    .A2(_02975_),
    .B1(_05978_),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2_1 _14781_ (.A(_09364_),
    .B(_02853_),
    .Y(_02978_));
 sky130_fd_sc_hd__nand2_1 _14782_ (.A(_02859_),
    .B(_02873_),
    .Y(_02979_));
 sky130_fd_sc_hd__o21ai_0 _14783_ (.A1(_05956_),
    .A2(_02888_),
    .B1(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__nor2_1 _14784_ (.A(_02955_),
    .B(_02889_),
    .Y(_02981_));
 sky130_fd_sc_hd__a22oi_1 _14785_ (.A1(_09357_),
    .A2(_02980_),
    .B1(_02981_),
    .B2(_09362_),
    .Y(_02982_));
 sky130_fd_sc_hd__o22ai_1 _14786_ (.A1(_02919_),
    .A2(_02978_),
    .B1(_02982_),
    .B2(_02853_),
    .Y(_02983_));
 sky130_fd_sc_hd__a2111oi_0 _14787_ (.A1(_09358_),
    .A2(_02972_),
    .B1(_02974_),
    .C1(_02976_),
    .D1(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__nor2_1 _14788_ (.A(_02943_),
    .B(_02984_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand2_1 _14789_ (.A(_09358_),
    .B(_02911_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand2_1 _14790_ (.A(_09357_),
    .B(_05953_),
    .Y(_02986_));
 sky130_fd_sc_hd__a21oi_1 _14791_ (.A1(_02985_),
    .A2(_02986_),
    .B1(_02906_),
    .Y(_02987_));
 sky130_fd_sc_hd__a21oi_1 _14792_ (.A1(_09362_),
    .A2(_02891_),
    .B1(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__nand2_1 _14793_ (.A(_02942_),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__nor3_1 _14794_ (.A(_02853_),
    .B(_02919_),
    .C(_02939_),
    .Y(_02990_));
 sky130_fd_sc_hd__nor2_1 _14795_ (.A(_02894_),
    .B(_02853_),
    .Y(_02991_));
 sky130_fd_sc_hd__nor2_1 _14796_ (.A(_05958_),
    .B(_05978_),
    .Y(_02992_));
 sky130_fd_sc_hd__a221oi_1 _14797_ (.A1(_09362_),
    .A2(_02991_),
    .B1(_02992_),
    .B2(_09364_),
    .C1(_05953_),
    .Y(_02993_));
 sky130_fd_sc_hd__a221oi_1 _14798_ (.A1(_09364_),
    .A2(_05958_),
    .B1(_02907_),
    .B2(_09358_),
    .C1(_02911_),
    .Y(_02994_));
 sky130_fd_sc_hd__o21ai_0 _14799_ (.A1(_02895_),
    .A2(_02879_),
    .B1(_09357_),
    .Y(_02995_));
 sky130_fd_sc_hd__o21ai_0 _14800_ (.A1(_02993_),
    .A2(_02994_),
    .B1(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__nor3_1 _14801_ (.A(_02989_),
    .B(_02990_),
    .C(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__o21ai_0 _14802_ (.A1(_02916_),
    .A2(_02997_),
    .B1(_05476_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _14803_ (.A(_05978_),
    .B(_02933_),
    .Y(_02998_));
 sky130_fd_sc_hd__o2bb2ai_1 _14804_ (.A1_N(_02950_),
    .A2_N(_02998_),
    .B1(_02879_),
    .B2(_02895_),
    .Y(_02999_));
 sky130_fd_sc_hd__nand2_1 _14805_ (.A(_09362_),
    .B(_02906_),
    .Y(_03000_));
 sky130_fd_sc_hd__nor2_1 _14806_ (.A(_02853_),
    .B(_02895_),
    .Y(_03001_));
 sky130_fd_sc_hd__o21ai_0 _14808_ (.A1(_05978_),
    .A2(_02980_),
    .B1(_09358_),
    .Y(_03003_));
 sky130_fd_sc_hd__o22ai_1 _14809_ (.A1(_02890_),
    .A2(_03000_),
    .B1(_03001_),
    .B2(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__a211oi_1 _14810_ (.A1(_09364_),
    .A2(_02891_),
    .B1(_02983_),
    .C1(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__a21oi_1 _14811_ (.A1(_02999_),
    .A2(_03005_),
    .B1(_02943_),
    .Y(_00725_));
 sky130_fd_sc_hd__o21ai_0 _14812_ (.A1(_09357_),
    .A2(_09364_),
    .B1(_02889_),
    .Y(_03006_));
 sky130_fd_sc_hd__nand2_1 _14813_ (.A(_09357_),
    .B(_02853_),
    .Y(_03007_));
 sky130_fd_sc_hd__a21oi_1 _14814_ (.A1(_09364_),
    .A2(_05978_),
    .B1(_09358_),
    .Y(_03008_));
 sky130_fd_sc_hd__a21oi_1 _14815_ (.A1(_03007_),
    .A2(_03008_),
    .B1(_02877_),
    .Y(_03009_));
 sky130_fd_sc_hd__a21oi_1 _14816_ (.A1(_09358_),
    .A2(_02925_),
    .B1(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _14817_ (.A(_05953_),
    .B(_02853_),
    .Y(_03011_));
 sky130_fd_sc_hd__or3_1 _14818_ (.A(_09358_),
    .B(_05953_),
    .C(_02853_),
    .X(_03012_));
 sky130_fd_sc_hd__o21ai_0 _14819_ (.A1(_09357_),
    .A2(_05978_),
    .B1(_02911_),
    .Y(_03013_));
 sky130_fd_sc_hd__nand2b_1 _14820_ (.A_N(_09362_),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_1 _14821_ (.A(_09358_),
    .B(_02895_),
    .Y(_03015_));
 sky130_fd_sc_hd__nor2_1 _14822_ (.A(_02919_),
    .B(_02929_),
    .Y(_03016_));
 sky130_fd_sc_hd__nand2_1 _14823_ (.A(_05978_),
    .B(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__o21ai_0 _14824_ (.A1(_05978_),
    .A2(_03015_),
    .B1(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__a41oi_1 _14825_ (.A1(_05958_),
    .A2(_03011_),
    .A3(_03012_),
    .A4(_03014_),
    .B1(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__a31oi_1 _14826_ (.A1(_03006_),
    .A2(_03010_),
    .A3(_03019_),
    .B1(_02943_),
    .Y(_00726_));
 sky130_fd_sc_hd__a21oi_1 _14827_ (.A1(_09362_),
    .A2(_02911_),
    .B1(_09357_),
    .Y(_03020_));
 sky130_fd_sc_hd__nor2_1 _14828_ (.A(_02906_),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__nand2_1 _14829_ (.A(_09364_),
    .B(_02907_),
    .Y(_03022_));
 sky130_fd_sc_hd__nand3_1 _14830_ (.A(_09358_),
    .B(_05958_),
    .C(_02853_),
    .Y(_03023_));
 sky130_fd_sc_hd__a21oi_1 _14831_ (.A1(_03022_),
    .A2(_03023_),
    .B1(_05953_),
    .Y(_03024_));
 sky130_fd_sc_hd__nor2_1 _14832_ (.A(_03021_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__a21oi_1 _14833_ (.A1(_02928_),
    .A2(_03025_),
    .B1(_02943_),
    .Y(_00727_));
 sky130_fd_sc_hd__o21ai_0 _14834_ (.A1(_09362_),
    .A2(_09364_),
    .B1(_02895_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand3_1 _14835_ (.A(_09357_),
    .B(_02853_),
    .C(_02980_),
    .Y(_03027_));
 sky130_fd_sc_hd__o211a_1 _14836_ (.A1(_02853_),
    .A2(_03026_),
    .B1(_02942_),
    .C1(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__nand2_1 _14837_ (.A(_09364_),
    .B(_02894_),
    .Y(_03029_));
 sky130_fd_sc_hd__nand2_1 _14838_ (.A(_09362_),
    .B(_02895_),
    .Y(_03030_));
 sky130_fd_sc_hd__o21ai_0 _14839_ (.A1(_02911_),
    .A2(_03029_),
    .B1(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__a21oi_1 _14840_ (.A1(_02853_),
    .A2(_03031_),
    .B1(_03018_),
    .Y(_03032_));
 sky130_fd_sc_hd__nor3_1 _14841_ (.A(_09357_),
    .B(_09362_),
    .C(_09364_),
    .Y(_03033_));
 sky130_fd_sc_hd__nor2_1 _14842_ (.A(_02911_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__o21ai_0 _14843_ (.A1(_09358_),
    .A2(_03034_),
    .B1(_02991_),
    .Y(_03035_));
 sky130_fd_sc_hd__nor2_1 _14844_ (.A(_09362_),
    .B(_02894_),
    .Y(_03036_));
 sky130_fd_sc_hd__nor2_1 _14845_ (.A(_02911_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__nor2_1 _14846_ (.A(_05978_),
    .B(_02895_),
    .Y(_03038_));
 sky130_fd_sc_hd__o221ai_1 _14847_ (.A1(_09358_),
    .A2(_02919_),
    .B1(_03037_),
    .B2(_09364_),
    .C1(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__nand4_1 _14848_ (.A(_03028_),
    .B(_03032_),
    .C(_03035_),
    .D(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__a21o_1 _14849_ (.A1(_05481_),
    .A2(_03040_),
    .B1(reset_hash),
    .X(_00728_));
 sky130_fd_sc_hd__o21ai_0 _14850_ (.A1(_02879_),
    .A2(_02957_),
    .B1(_09362_),
    .Y(_03041_));
 sky130_fd_sc_hd__nor2_1 _14851_ (.A(_02911_),
    .B(_02932_),
    .Y(_03042_));
 sky130_fd_sc_hd__nor3_1 _14852_ (.A(_05953_),
    .B(_02853_),
    .C(_02922_),
    .Y(_03043_));
 sky130_fd_sc_hd__o21ai_0 _14853_ (.A1(_03042_),
    .A2(_03043_),
    .B1(_05958_),
    .Y(_03044_));
 sky130_fd_sc_hd__a41oi_1 _14854_ (.A1(_02998_),
    .A2(_03032_),
    .A3(_03041_),
    .A4(_03044_),
    .B1(_02943_),
    .Y(_00729_));
 sky130_fd_sc_hd__o22ai_1 _14855_ (.A1(_02920_),
    .A2(_02949_),
    .B1(_03029_),
    .B2(_02853_),
    .Y(_03045_));
 sky130_fd_sc_hd__a21oi_1 _14856_ (.A1(_05953_),
    .A2(_03045_),
    .B1(_02990_),
    .Y(_03046_));
 sky130_fd_sc_hd__and3_1 _14857_ (.A(_05476_),
    .B(_02942_),
    .C(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__nor2_1 _14858_ (.A(_02894_),
    .B(_03020_),
    .Y(_03048_));
 sky130_fd_sc_hd__a22oi_1 _14859_ (.A1(_09364_),
    .A2(_05953_),
    .B1(_02877_),
    .B2(_09358_),
    .Y(_03049_));
 sky130_fd_sc_hd__o21ai_0 _14860_ (.A1(_02889_),
    .A2(_03049_),
    .B1(_02853_),
    .Y(_03050_));
 sky130_fd_sc_hd__o31ai_1 _14861_ (.A1(_02853_),
    .A2(_02974_),
    .A3(_03048_),
    .B1(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__nor2_1 _14862_ (.A(reset_hash),
    .B(_05481_),
    .Y(_03052_));
 sky130_fd_sc_hd__a31oi_1 _14863_ (.A1(_02893_),
    .A2(_03047_),
    .A3(_03051_),
    .B1(_03052_),
    .Y(_00730_));
 sky130_fd_sc_hd__nor2_1 _14864_ (.A(_02919_),
    .B(_02932_),
    .Y(_03053_));
 sky130_fd_sc_hd__a21oi_1 _14865_ (.A1(_09362_),
    .A2(_02894_),
    .B1(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__nor2_1 _14866_ (.A(_02853_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__a31oi_1 _14867_ (.A1(_09357_),
    .A2(_02853_),
    .A3(_02889_),
    .B1(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__a31oi_1 _14868_ (.A1(_09364_),
    .A2(_02894_),
    .A3(_05978_),
    .B1(_02902_),
    .Y(_03057_));
 sky130_fd_sc_hd__nor2_1 _14869_ (.A(_05953_),
    .B(_02853_),
    .Y(_03058_));
 sky130_fd_sc_hd__o21ai_0 _14870_ (.A1(_02957_),
    .A2(_03058_),
    .B1(_09358_),
    .Y(_03059_));
 sky130_fd_sc_hd__o21ai_0 _14871_ (.A1(_05953_),
    .A2(_03057_),
    .B1(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__a21oi_1 _14872_ (.A1(_02853_),
    .A2(_03016_),
    .B1(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__a21oi_1 _14873_ (.A1(_03056_),
    .A2(_03061_),
    .B1(_02943_),
    .Y(_00731_));
 sky130_fd_sc_hd__o21ai_0 _14874_ (.A1(_02927_),
    .A2(_02933_),
    .B1(_02853_),
    .Y(_03062_));
 sky130_fd_sc_hd__nor2_1 _14875_ (.A(_05978_),
    .B(_02919_),
    .Y(_03063_));
 sky130_fd_sc_hd__o21ai_0 _14876_ (.A1(_02991_),
    .A2(_03063_),
    .B1(_09364_),
    .Y(_03064_));
 sky130_fd_sc_hd__nor2_1 _14877_ (.A(_02991_),
    .B(_02992_),
    .Y(_03065_));
 sky130_fd_sc_hd__o21ai_0 _14878_ (.A1(_02853_),
    .A2(_02895_),
    .B1(_02949_),
    .Y(_03066_));
 sky130_fd_sc_hd__a22oi_1 _14879_ (.A1(_09358_),
    .A2(_03065_),
    .B1(_03066_),
    .B2(_09362_),
    .Y(_03067_));
 sky130_fd_sc_hd__a31oi_1 _14880_ (.A1(_03062_),
    .A2(_03064_),
    .A3(_03067_),
    .B1(_02943_),
    .Y(_00732_));
 sky130_fd_sc_hd__a21oi_1 _14881_ (.A1(_09362_),
    .A2(_02894_),
    .B1(_09358_),
    .Y(_03068_));
 sky130_fd_sc_hd__o221ai_1 _14882_ (.A1(_02922_),
    .A2(_02905_),
    .B1(_03068_),
    .B2(_05978_),
    .C1(_02911_),
    .Y(_03069_));
 sky130_fd_sc_hd__nand2_1 _14883_ (.A(_09362_),
    .B(_02992_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand3_1 _14884_ (.A(_05953_),
    .B(_03022_),
    .C(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__nand2_1 _14885_ (.A(_02980_),
    .B(_02871_),
    .Y(_03072_));
 sky130_fd_sc_hd__o21ai_0 _14886_ (.A1(_05953_),
    .A2(_03029_),
    .B1(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__a222oi_1 _14887_ (.A1(_02889_),
    .A2(_02902_),
    .B1(_03069_),
    .B2(_03071_),
    .C1(_03073_),
    .C2(_05978_),
    .Y(_03074_));
 sky130_fd_sc_hd__nor2_1 _14888_ (.A(_02943_),
    .B(_03074_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand2_1 _14889_ (.A(_09358_),
    .B(_02981_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2_1 _14890_ (.A(_02950_),
    .B(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__o211ai_1 _14891_ (.A1(_09358_),
    .A2(_02930_),
    .B1(_03076_),
    .C1(_05978_),
    .Y(_03077_));
 sky130_fd_sc_hd__nor2_1 _14892_ (.A(_05953_),
    .B(_02938_),
    .Y(_03078_));
 sky130_fd_sc_hd__a21oi_1 _14893_ (.A1(_05953_),
    .A2(_03068_),
    .B1(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_1 _14894_ (.A(_02853_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__a21oi_1 _14895_ (.A1(_03077_),
    .A2(_03080_),
    .B1(_02943_),
    .Y(_00734_));
 sky130_fd_sc_hd__a21oi_1 _14896_ (.A1(_09362_),
    .A2(_05953_),
    .B1(_09364_),
    .Y(_03081_));
 sky130_fd_sc_hd__nand3_1 _14897_ (.A(_09357_),
    .B(_02911_),
    .C(_02853_),
    .Y(_03082_));
 sky130_fd_sc_hd__o21ai_0 _14898_ (.A1(_02853_),
    .A2(_03081_),
    .B1(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__nand2_1 _14899_ (.A(_02911_),
    .B(_05978_),
    .Y(_03084_));
 sky130_fd_sc_hd__a21oi_1 _14900_ (.A1(_09364_),
    .A2(_02894_),
    .B1(_09358_),
    .Y(_03085_));
 sky130_fd_sc_hd__nor2_1 _14901_ (.A(_03084_),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__a21oi_1 _14902_ (.A1(_05958_),
    .A2(_03083_),
    .B1(_03086_),
    .Y(_03087_));
 sky130_fd_sc_hd__a31oi_1 _14903_ (.A1(_02924_),
    .A2(_03047_),
    .A3(_03087_),
    .B1(_03052_),
    .Y(_00735_));
 sky130_fd_sc_hd__a211oi_1 _14904_ (.A1(_05953_),
    .A2(_02934_),
    .B1(_03078_),
    .C1(_05978_),
    .Y(_03088_));
 sky130_fd_sc_hd__a21oi_1 _14905_ (.A1(_09362_),
    .A2(_02972_),
    .B1(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__a21oi_1 _14906_ (.A1(_02937_),
    .A2(_03089_),
    .B1(_02943_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand2_1 _14907_ (.A(_09364_),
    .B(_03058_),
    .Y(_03090_));
 sky130_fd_sc_hd__o21ai_0 _14908_ (.A1(_02920_),
    .A2(_03011_),
    .B1(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__o22ai_1 _14909_ (.A1(_02919_),
    .A2(_02885_),
    .B1(_03006_),
    .B2(_02853_),
    .Y(_03092_));
 sky130_fd_sc_hd__a21oi_1 _14910_ (.A1(_05958_),
    .A2(_03091_),
    .B1(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__o21ai_0 _14911_ (.A1(_05953_),
    .A2(_02949_),
    .B1(_02919_),
    .Y(_03094_));
 sky130_fd_sc_hd__a21oi_1 _14912_ (.A1(_09358_),
    .A2(_03094_),
    .B1(_02974_),
    .Y(_03095_));
 sky130_fd_sc_hd__and3_1 _14913_ (.A(_02961_),
    .B(_03093_),
    .C(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__o21ai_0 _14914_ (.A1(_02916_),
    .A2(_03096_),
    .B1(_05476_),
    .Y(_00737_));
 sky130_fd_sc_hd__nor3_1 _14915_ (.A(_09357_),
    .B(_09358_),
    .C(_09364_),
    .Y(_03097_));
 sky130_fd_sc_hd__o21ai_0 _14916_ (.A1(_02919_),
    .A2(_03097_),
    .B1(_03026_),
    .Y(_03098_));
 sky130_fd_sc_hd__a21oi_1 _14917_ (.A1(_09358_),
    .A2(_02889_),
    .B1(_02974_),
    .Y(_03099_));
 sky130_fd_sc_hd__o22ai_1 _14918_ (.A1(_02949_),
    .A2(_02973_),
    .B1(_03099_),
    .B2(_02853_),
    .Y(_03100_));
 sky130_fd_sc_hd__a21oi_1 _14919_ (.A1(_05978_),
    .A2(_03098_),
    .B1(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _14920_ (.A(_03011_),
    .B(_03084_),
    .Y(_03102_));
 sky130_fd_sc_hd__nand3_1 _14921_ (.A(_09357_),
    .B(_05958_),
    .C(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__a31oi_1 _14922_ (.A1(_02924_),
    .A2(_03101_),
    .A3(_03103_),
    .B1(_02943_),
    .Y(_00738_));
 sky130_fd_sc_hd__a21oi_1 _14923_ (.A1(_09358_),
    .A2(_05958_),
    .B1(_09364_),
    .Y(_03104_));
 sky130_fd_sc_hd__nor2_1 _14924_ (.A(_02950_),
    .B(_02905_),
    .Y(_03105_));
 sky130_fd_sc_hd__a21oi_1 _14925_ (.A1(_09362_),
    .A2(_02905_),
    .B1(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__o22a_1 _14926_ (.A1(_03011_),
    .A2(_03104_),
    .B1(_03106_),
    .B2(_05953_),
    .X(_03107_));
 sky130_fd_sc_hd__a21oi_1 _14927_ (.A1(_03010_),
    .A2(_03107_),
    .B1(_02943_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _14928_ (.A(_02853_),
    .B(_02940_),
    .Y(_03108_));
 sky130_fd_sc_hd__o21ai_0 _14929_ (.A1(_02879_),
    .A2(_02957_),
    .B1(_09364_),
    .Y(_03109_));
 sky130_fd_sc_hd__a21oi_1 _14930_ (.A1(_09362_),
    .A2(_02889_),
    .B1(_09358_),
    .Y(_03110_));
 sky130_fd_sc_hd__nor2_1 _14931_ (.A(_02981_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__nor2_1 _14932_ (.A(_03055_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__a31oi_1 _14933_ (.A1(_03108_),
    .A2(_03109_),
    .A3(_03112_),
    .B1(_02943_),
    .Y(_00740_));
 sky130_fd_sc_hd__nor2_1 _14934_ (.A(_02877_),
    .B(_02901_),
    .Y(_03113_));
 sky130_fd_sc_hd__a21oi_1 _14935_ (.A1(_09362_),
    .A2(_05958_),
    .B1(_09357_),
    .Y(_03114_));
 sky130_fd_sc_hd__o21ai_0 _14936_ (.A1(_02955_),
    .A2(_03114_),
    .B1(_02853_),
    .Y(_03115_));
 sky130_fd_sc_hd__o41ai_1 _14937_ (.A1(_02853_),
    .A2(_02931_),
    .A3(_03053_),
    .A4(_03113_),
    .B1(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__a21oi_1 _14938_ (.A1(_02892_),
    .A2(_03116_),
    .B1(_02943_),
    .Y(_00741_));
 sky130_fd_sc_hd__a22oi_1 _14939_ (.A1(_02911_),
    .A2(_02853_),
    .B1(_02885_),
    .B2(_02950_),
    .Y(_03117_));
 sky130_fd_sc_hd__nor2_1 _14940_ (.A(_09358_),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__o32ai_1 _14941_ (.A1(_02894_),
    .A2(_02952_),
    .A3(_03118_),
    .B1(_02877_),
    .B2(_02885_),
    .Y(_03119_));
 sky130_fd_sc_hd__nor2_1 _14942_ (.A(_03009_),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__a21oi_1 _14943_ (.A1(_03101_),
    .A2(_03120_),
    .B1(_02943_),
    .Y(_00742_));
 sky130_fd_sc_hd__nand3_1 _14944_ (.A(_09364_),
    .B(_02853_),
    .C(_02955_),
    .Y(_03121_));
 sky130_fd_sc_hd__o21ai_0 _14945_ (.A1(_02955_),
    .A2(_02972_),
    .B1(_09358_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_1 _14946_ (.A(_03121_),
    .B(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__nand2_1 _14947_ (.A(_09357_),
    .B(_05978_),
    .Y(_03124_));
 sky130_fd_sc_hd__nand2_1 _14948_ (.A(_09362_),
    .B(_03102_),
    .Y(_03125_));
 sky130_fd_sc_hd__a21oi_1 _14949_ (.A1(_03124_),
    .A2(_03125_),
    .B1(_02894_),
    .Y(_03126_));
 sky130_fd_sc_hd__nand2_1 _14950_ (.A(_09364_),
    .B(_03065_),
    .Y(_03127_));
 sky130_fd_sc_hd__a21oi_1 _14951_ (.A1(_02908_),
    .A2(_03127_),
    .B1(_02911_),
    .Y(_03128_));
 sky130_fd_sc_hd__nor4b_1 _14952_ (.A(_03123_),
    .B(_03126_),
    .C(_03128_),
    .D_N(_02942_),
    .Y(_03129_));
 sky130_fd_sc_hd__o21ai_0 _14953_ (.A1(_02916_),
    .A2(_03129_),
    .B1(_05476_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_1 _14954_ (.A(_09357_),
    .B(_02877_),
    .Y(_03130_));
 sky130_fd_sc_hd__o21ai_0 _14955_ (.A1(_09358_),
    .A2(_05953_),
    .B1(_05958_),
    .Y(_03131_));
 sky130_fd_sc_hd__a221o_1 _14956_ (.A1(_02889_),
    .A2(_02932_),
    .B1(_03130_),
    .B2(_03131_),
    .C1(_05978_),
    .X(_03132_));
 sky130_fd_sc_hd__nand2_1 _14957_ (.A(_02853_),
    .B(_02929_),
    .Y(_03133_));
 sky130_fd_sc_hd__nand2_1 _14958_ (.A(_05978_),
    .B(_02939_),
    .Y(_03134_));
 sky130_fd_sc_hd__nand3_1 _14959_ (.A(_02980_),
    .B(_03133_),
    .C(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__a41oi_1 _14960_ (.A1(_03035_),
    .A2(_03121_),
    .A3(_03132_),
    .A4(_03135_),
    .B1(_02943_),
    .Y(_00744_));
 sky130_fd_sc_hd__nor2_1 _14961_ (.A(_09357_),
    .B(_09358_),
    .Y(_03136_));
 sky130_fd_sc_hd__nor2_1 _14962_ (.A(_02877_),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__nor2_1 _14963_ (.A(_03016_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__nor2_1 _14964_ (.A(_09358_),
    .B(_02853_),
    .Y(_03139_));
 sky130_fd_sc_hd__nor3_1 _14965_ (.A(_09362_),
    .B(_05953_),
    .C(_05978_),
    .Y(_03140_));
 sky130_fd_sc_hd__nor2_1 _14966_ (.A(_03139_),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__o21ai_0 _14967_ (.A1(_05978_),
    .A2(_02922_),
    .B1(_05953_),
    .Y(_03142_));
 sky130_fd_sc_hd__o211ai_1 _14968_ (.A1(_09357_),
    .A2(_03141_),
    .B1(_03142_),
    .C1(_05958_),
    .Y(_03143_));
 sky130_fd_sc_hd__o2111a_1 _14969_ (.A1(_02853_),
    .A2(_03138_),
    .B1(_03143_),
    .C1(_02988_),
    .D1(_02942_),
    .X(_03144_));
 sky130_fd_sc_hd__o21ai_0 _14970_ (.A1(_02916_),
    .A2(_03144_),
    .B1(_05476_),
    .Y(_00745_));
 sky130_fd_sc_hd__o21ai_0 _14971_ (.A1(_05958_),
    .A2(_02879_),
    .B1(_09362_),
    .Y(_03145_));
 sky130_fd_sc_hd__a21oi_1 _14972_ (.A1(_03072_),
    .A2(_03006_),
    .B1(_05978_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand2_1 _14973_ (.A(_09364_),
    .B(_03102_),
    .Y(_03147_));
 sky130_fd_sc_hd__nand3_1 _14974_ (.A(_09358_),
    .B(_02911_),
    .C(_02853_),
    .Y(_03148_));
 sky130_fd_sc_hd__a21oi_1 _14975_ (.A1(_03147_),
    .A2(_03148_),
    .B1(_05958_),
    .Y(_03149_));
 sky130_fd_sc_hd__a2111oi_0 _14976_ (.A1(_09357_),
    .A2(_02991_),
    .B1(_02990_),
    .C1(_03146_),
    .D1(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__and3_1 _14977_ (.A(_02942_),
    .B(_03145_),
    .C(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__o21ai_0 _14978_ (.A1(_02916_),
    .A2(_03151_),
    .B1(_05476_),
    .Y(_00746_));
 sky130_fd_sc_hd__nor3_1 _14979_ (.A(_03055_),
    .B(_03092_),
    .C(_03119_),
    .Y(_03152_));
 sky130_fd_sc_hd__nor2_1 _14980_ (.A(_02943_),
    .B(_03152_),
    .Y(_00747_));
 sky130_fd_sc_hd__o22ai_1 _14981_ (.A1(_02919_),
    .A2(_02922_),
    .B1(_02930_),
    .B2(_02901_),
    .Y(_03153_));
 sky130_fd_sc_hd__nand2_1 _14982_ (.A(_02853_),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__nand2_1 _14983_ (.A(_09358_),
    .B(_02980_),
    .Y(_03155_));
 sky130_fd_sc_hd__a21oi_1 _14984_ (.A1(_03138_),
    .A2(_03155_),
    .B1(_02853_),
    .Y(_03156_));
 sky130_fd_sc_hd__nor2_1 _14985_ (.A(_03126_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__a31oi_1 _14986_ (.A1(_02924_),
    .A2(_03154_),
    .A3(_03157_),
    .B1(_02943_),
    .Y(_00748_));
 sky130_fd_sc_hd__o311a_1 _14987_ (.A1(_05978_),
    .A2(_02877_),
    .A3(_03097_),
    .B1(_02942_),
    .C1(_05476_),
    .X(_03158_));
 sky130_fd_sc_hd__nand2_1 _14988_ (.A(_05953_),
    .B(_02932_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_1 _14989_ (.A(_02911_),
    .B(_02922_),
    .Y(_03160_));
 sky130_fd_sc_hd__a32oi_1 _14990_ (.A1(_02991_),
    .A2(_03159_),
    .A3(_03160_),
    .B1(_03063_),
    .B2(_09362_),
    .Y(_03161_));
 sky130_fd_sc_hd__a41oi_1 _14991_ (.A1(_03056_),
    .A2(_03132_),
    .A3(_03158_),
    .A4(_03161_),
    .B1(_03052_),
    .Y(_00749_));
 sky130_fd_sc_hd__a21oi_1 _14992_ (.A1(_02920_),
    .A2(_02922_),
    .B1(_02919_),
    .Y(_03162_));
 sky130_fd_sc_hd__o221ai_1 _14993_ (.A1(_02950_),
    .A2(_02894_),
    .B1(_02920_),
    .B2(_02930_),
    .C1(_05978_),
    .Y(_03163_));
 sky130_fd_sc_hd__o21ai_0 _14994_ (.A1(_05978_),
    .A2(_03162_),
    .B1(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__a221oi_1 _14995_ (.A1(_02889_),
    .A2(_02902_),
    .B1(_03073_),
    .B2(_05978_),
    .C1(_03100_),
    .Y(_03165_));
 sky130_fd_sc_hd__a31oi_1 _14996_ (.A1(_03158_),
    .A2(_03164_),
    .A3(_03165_),
    .B1(_03052_),
    .Y(_00750_));
 sky130_fd_sc_hd__nor2_1 _14997_ (.A(_02968_),
    .B(_03078_),
    .Y(_03166_));
 sky130_fd_sc_hd__o21ai_0 _14998_ (.A1(_09358_),
    .A2(_03166_),
    .B1(_05958_),
    .Y(_03167_));
 sky130_fd_sc_hd__a21oi_1 _14999_ (.A1(_03072_),
    .A2(_03167_),
    .B1(_05978_),
    .Y(_03168_));
 sky130_fd_sc_hd__a211oi_1 _15000_ (.A1(_05978_),
    .A2(_02927_),
    .B1(_03156_),
    .C1(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_1 _15001_ (.A(_03028_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__a21o_1 _15002_ (.A1(_05481_),
    .A2(_03170_),
    .B1(reset_hash),
    .X(_00751_));
 sky130_fd_sc_hd__nor2_1 _15004_ (.A(_09347_),
    .B(_09348_),
    .Y(_03172_));
 sky130_fd_sc_hd__nor2_1 _15006_ (.A(_09350_),
    .B(_09352_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand2_1 _15007_ (.A(_03172_),
    .B(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand2_1 _15008_ (.A(_02918_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__xnor2_1 _15009_ (.A(\count_hash2[4] ),
    .B(_05460_),
    .Y(_03177_));
 sky130_fd_sc_hd__xor2_1 _15010_ (.A(\count_hash2[5] ),
    .B(_05471_),
    .X(_03178_));
 sky130_fd_sc_hd__nand2_1 _15011_ (.A(_03177_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__xnor2_2 _15013_ (.A(\count_hash2[3] ),
    .B(_09354_),
    .Y(_03181_));
 sky130_fd_sc_hd__nand2_1 _15014_ (.A(_03181_),
    .B(_03172_),
    .Y(_03182_));
 sky130_fd_sc_hd__clkinv_1 _15015_ (.A(_09347_),
    .Y(_03183_));
 sky130_fd_sc_hd__nor2_1 _15019_ (.A(_09352_),
    .B(_03181_),
    .Y(_03187_));
 sky130_fd_sc_hd__o21ai_0 _15020_ (.A1(_03183_),
    .A2(_03177_),
    .B1(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__inv_1 _15021_ (.A(_09350_),
    .Y(_03189_));
 sky130_fd_sc_hd__nor2_1 _15022_ (.A(_05461_),
    .B(_03178_),
    .Y(_03190_));
 sky130_fd_sc_hd__a22oi_1 _15023_ (.A1(_03182_),
    .A2(_03190_),
    .B1(_03188_),
    .B2(_05461_),
    .Y(_03191_));
 sky130_fd_sc_hd__nand2_1 _15025_ (.A(_05461_),
    .B(_05458_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2_1 _15026_ (.A(_03177_),
    .B(_03181_),
    .Y(_03194_));
 sky130_fd_sc_hd__and2_1 _15027_ (.A(_03193_),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__nor3_1 _15030_ (.A(_09347_),
    .B(_09348_),
    .C(_09350_),
    .Y(_03198_));
 sky130_fd_sc_hd__nand2_1 _15031_ (.A(_03177_),
    .B(_05458_),
    .Y(_03199_));
 sky130_fd_sc_hd__nor2_1 _15032_ (.A(_03198_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__a21oi_1 _15033_ (.A1(_09352_),
    .A2(_03195_),
    .B1(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__o22ai_1 _15034_ (.A1(_03189_),
    .A2(_03191_),
    .B1(_03201_),
    .B2(_05472_),
    .Y(_03202_));
 sky130_fd_sc_hd__a31oi_1 _15035_ (.A1(_03179_),
    .A2(_03182_),
    .A3(_03188_),
    .B1(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__o21ai_0 _15036_ (.A1(_03176_),
    .A2(_03203_),
    .B1(_05476_),
    .Y(_00752_));
 sky130_fd_sc_hd__o21ai_0 _15043_ (.A1(_03177_),
    .A2(_03172_),
    .B1(_03181_),
    .Y(_03210_));
 sky130_fd_sc_hd__a32oi_1 _15045_ (.A1(_09352_),
    .A2(_05461_),
    .A3(_03182_),
    .B1(_03210_),
    .B2(_09350_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _15047_ (.A(_05461_),
    .B(_05472_),
    .Y(_03214_));
 sky130_fd_sc_hd__nor2_1 _15048_ (.A(_05458_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__o21ai_0 _15049_ (.A1(_03172_),
    .A2(_03215_),
    .B1(_03174_),
    .Y(_03216_));
 sky130_fd_sc_hd__nor2_1 _15052_ (.A(_05461_),
    .B(_05472_),
    .Y(_03219_));
 sky130_fd_sc_hd__nand3_1 _15053_ (.A(_09350_),
    .B(_03181_),
    .C(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__a21oi_1 _15054_ (.A1(_03183_),
    .A2(_05461_),
    .B1(_05472_),
    .Y(_03221_));
 sky130_fd_sc_hd__o21ai_0 _15056_ (.A1(_09348_),
    .A2(_03177_),
    .B1(_03179_),
    .Y(_03223_));
 sky130_fd_sc_hd__a21oi_1 _15058_ (.A1(_09348_),
    .A2(_03181_),
    .B1(_09347_),
    .Y(_03225_));
 sky130_fd_sc_hd__a21oi_1 _15059_ (.A1(_03181_),
    .A2(_03223_),
    .B1(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__o221ai_1 _15060_ (.A1(_03181_),
    .A2(_03221_),
    .B1(_03226_),
    .B2(_09352_),
    .C1(_03214_),
    .Y(_03227_));
 sky130_fd_sc_hd__o2111ai_1 _15061_ (.A1(_03178_),
    .A2(_03212_),
    .B1(_03216_),
    .C1(_03220_),
    .D1(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_1 _15062_ (.A(_05481_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _15063_ (.A(_05476_),
    .B(_03229_),
    .Y(_00753_));
 sky130_fd_sc_hd__a21oi_1 _15064_ (.A1(_09352_),
    .A2(_05461_),
    .B1(_09347_),
    .Y(_03230_));
 sky130_fd_sc_hd__nand2_1 _15065_ (.A(_09348_),
    .B(_03177_),
    .Y(_03231_));
 sky130_fd_sc_hd__o21ai_0 _15066_ (.A1(_03181_),
    .A2(_03230_),
    .B1(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__nand2_1 _15067_ (.A(_05461_),
    .B(_03181_),
    .Y(_03233_));
 sky130_fd_sc_hd__nor3_1 _15068_ (.A(_03178_),
    .B(_03198_),
    .C(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__a21oi_1 _15069_ (.A1(_03178_),
    .A2(_03232_),
    .B1(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__nor2_1 _15071_ (.A(_03177_),
    .B(_03178_),
    .Y(_03237_));
 sky130_fd_sc_hd__nor2_1 _15072_ (.A(_03219_),
    .B(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand2_1 _15073_ (.A(_09348_),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__nor2_1 _15075_ (.A(_03177_),
    .B(_05472_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _15076_ (.A(_09347_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__a21oi_1 _15078_ (.A1(_03239_),
    .A2(_03242_),
    .B1(_05458_),
    .Y(_03244_));
 sky130_fd_sc_hd__or2_2 _15079_ (.A(_09348_),
    .B(_09350_),
    .X(_03245_));
 sky130_fd_sc_hd__nor3_1 _15080_ (.A(_09347_),
    .B(_09350_),
    .C(_09352_),
    .Y(_03246_));
 sky130_fd_sc_hd__nand2_1 _15081_ (.A(_03181_),
    .B(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__o211ai_1 _15082_ (.A1(_03181_),
    .A2(_03245_),
    .B1(_03190_),
    .C1(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__nor2_1 _15083_ (.A(_03181_),
    .B(_05472_),
    .Y(_03249_));
 sky130_fd_sc_hd__nor3_1 _15084_ (.A(_09347_),
    .B(_09352_),
    .C(_03245_),
    .Y(_03250_));
 sky130_fd_sc_hd__o21ai_0 _15085_ (.A1(_05461_),
    .A2(_03249_),
    .B1(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__a21oi_1 _15086_ (.A1(_03178_),
    .A2(_03175_),
    .B1(_05458_),
    .Y(_03252_));
 sky130_fd_sc_hd__nor3_1 _15088_ (.A(_09347_),
    .B(_09352_),
    .C(_03178_),
    .Y(_03254_));
 sky130_fd_sc_hd__o21ai_0 _15090_ (.A1(_03252_),
    .A2(_03254_),
    .B1(_03177_),
    .Y(_03256_));
 sky130_fd_sc_hd__nand3_1 _15091_ (.A(_03248_),
    .B(_03251_),
    .C(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__nor2_1 _15092_ (.A(_03244_),
    .B(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__a21oi_1 _15093_ (.A1(_03235_),
    .A2(_03258_),
    .B1(_05482_),
    .Y(_00754_));
 sky130_fd_sc_hd__nand2_1 _15095_ (.A(_05458_),
    .B(_05472_),
    .Y(_03260_));
 sky130_fd_sc_hd__nand2_1 _15096_ (.A(_05461_),
    .B(_03178_),
    .Y(_03261_));
 sky130_fd_sc_hd__o22ai_1 _15097_ (.A1(_05461_),
    .A2(_03260_),
    .B1(_03261_),
    .B2(_05458_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _15098_ (.A(_03179_),
    .B(_03214_),
    .Y(_03263_));
 sky130_fd_sc_hd__a21oi_1 _15099_ (.A1(_03189_),
    .A2(_03193_),
    .B1(_05472_),
    .Y(_03264_));
 sky130_fd_sc_hd__a21oi_1 _15100_ (.A1(_03250_),
    .A2(_03241_),
    .B1(_03190_),
    .Y(_03265_));
 sky130_fd_sc_hd__o22ai_1 _15101_ (.A1(_09347_),
    .A2(_03264_),
    .B1(_03265_),
    .B2(_03181_),
    .Y(_03266_));
 sky130_fd_sc_hd__a21oi_1 _15102_ (.A1(_03181_),
    .A2(_03263_),
    .B1(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__a21oi_1 _15103_ (.A1(_09348_),
    .A2(_03262_),
    .B1(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__nor2_1 _15104_ (.A(_03176_),
    .B(_03268_),
    .Y(_00755_));
 sky130_fd_sc_hd__nor2_1 _15105_ (.A(_05472_),
    .B(_03172_),
    .Y(_03269_));
 sky130_fd_sc_hd__nor2_1 _15106_ (.A(_09352_),
    .B(_03245_),
    .Y(_03270_));
 sky130_fd_sc_hd__nor2_1 _15107_ (.A(_03178_),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__nor2_1 _15108_ (.A(_05461_),
    .B(_03181_),
    .Y(_03272_));
 sky130_fd_sc_hd__o21ai_0 _15109_ (.A1(_03269_),
    .A2(_03271_),
    .B1(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__nor2_1 _15110_ (.A(_03177_),
    .B(_03181_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_1 _15111_ (.A(_03245_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__o21ai_0 _15112_ (.A1(_03183_),
    .A2(_03195_),
    .B1(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_1 _15113_ (.A(_03178_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__nor2_1 _15114_ (.A(_03183_),
    .B(_05461_),
    .Y(_03278_));
 sky130_fd_sc_hd__a211o_1 _15116_ (.A1(_09352_),
    .A2(_05461_),
    .B1(_03278_),
    .C1(_09348_),
    .X(_03280_));
 sky130_fd_sc_hd__nand2_1 _15117_ (.A(_03181_),
    .B(_03190_),
    .Y(_03281_));
 sky130_fd_sc_hd__o21ai_0 _15118_ (.A1(_03174_),
    .A2(_03281_),
    .B1(_03175_),
    .Y(_03282_));
 sky130_fd_sc_hd__a31oi_1 _15119_ (.A1(_05472_),
    .A2(_03199_),
    .A3(_03280_),
    .B1(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__a31oi_1 _15120_ (.A1(_03273_),
    .A2(_03277_),
    .A3(_03283_),
    .B1(_05482_),
    .Y(_00756_));
 sky130_fd_sc_hd__o21ai_0 _15121_ (.A1(_09348_),
    .A2(_09352_),
    .B1(_03238_),
    .Y(_03284_));
 sky130_fd_sc_hd__a21oi_1 _15122_ (.A1(_03242_),
    .A2(_03284_),
    .B1(_05458_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _15123_ (.A(_03177_),
    .B(_05472_),
    .Y(_03286_));
 sky130_fd_sc_hd__a221oi_1 _15124_ (.A1(_09347_),
    .A2(_03286_),
    .B1(_03241_),
    .B2(_09348_),
    .C1(_09352_),
    .Y(_03287_));
 sky130_fd_sc_hd__nor2_1 _15125_ (.A(_03181_),
    .B(_03178_),
    .Y(_03288_));
 sky130_fd_sc_hd__a22oi_1 _15126_ (.A1(_09352_),
    .A2(_03178_),
    .B1(_03245_),
    .B2(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__o22ai_1 _15127_ (.A1(_03181_),
    .A2(_03287_),
    .B1(_03289_),
    .B2(_05461_),
    .Y(_03290_));
 sky130_fd_sc_hd__nor2_1 _15128_ (.A(_05482_),
    .B(_03250_),
    .Y(_03291_));
 sky130_fd_sc_hd__o21ai_0 _15129_ (.A1(_03285_),
    .A2(_03290_),
    .B1(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__nand2_1 _15130_ (.A(_05476_),
    .B(_03292_),
    .Y(_00757_));
 sky130_fd_sc_hd__nor2_1 _15131_ (.A(_03177_),
    .B(_05458_),
    .Y(_03293_));
 sky130_fd_sc_hd__a21oi_1 _15132_ (.A1(_03177_),
    .A2(_03182_),
    .B1(_09350_),
    .Y(_03294_));
 sky130_fd_sc_hd__nor2_1 _15133_ (.A(_09352_),
    .B(_03199_),
    .Y(_03295_));
 sky130_fd_sc_hd__nor4_1 _15134_ (.A(_05472_),
    .B(_03293_),
    .C(_03294_),
    .D(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_1 _15135_ (.A(_09350_),
    .B(_03219_),
    .Y(_03297_));
 sky130_fd_sc_hd__nand2_1 _15136_ (.A(_09348_),
    .B(_05461_),
    .Y(_03298_));
 sky130_fd_sc_hd__a221oi_1 _15137_ (.A1(_09350_),
    .A2(_03190_),
    .B1(_03238_),
    .B2(_09347_),
    .C1(_05458_),
    .Y(_03299_));
 sky130_fd_sc_hd__a31oi_1 _15138_ (.A1(_05458_),
    .A2(_03297_),
    .A3(_03298_),
    .B1(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__nor2_1 _15139_ (.A(_03296_),
    .B(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__nor2_1 _15140_ (.A(_03176_),
    .B(_03301_),
    .Y(_00758_));
 sky130_fd_sc_hd__a22oi_1 _15141_ (.A1(_03175_),
    .A2(_03219_),
    .B1(_03237_),
    .B2(_09350_),
    .Y(_03302_));
 sky130_fd_sc_hd__nor2_1 _15142_ (.A(_03181_),
    .B(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__nand2_1 _15143_ (.A(_03193_),
    .B(_03194_),
    .Y(_03304_));
 sky130_fd_sc_hd__a221oi_1 _15144_ (.A1(_09352_),
    .A2(_03274_),
    .B1(_03304_),
    .B2(_09348_),
    .C1(_05472_),
    .Y(_03305_));
 sky130_fd_sc_hd__a221oi_1 _15145_ (.A1(_09352_),
    .A2(_03181_),
    .B1(_03272_),
    .B2(_09347_),
    .C1(_03178_),
    .Y(_03306_));
 sky130_fd_sc_hd__nor2_1 _15146_ (.A(_09347_),
    .B(_09350_),
    .Y(_03307_));
 sky130_fd_sc_hd__o32ai_1 _15147_ (.A1(_05472_),
    .A2(_03233_),
    .A3(_03307_),
    .B1(_03260_),
    .B2(_03231_),
    .Y(_03308_));
 sky130_fd_sc_hd__a21oi_1 _15148_ (.A1(_09352_),
    .A2(_03262_),
    .B1(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__o21ai_0 _15149_ (.A1(_03305_),
    .A2(_03306_),
    .B1(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__o21ai_0 _15150_ (.A1(_03303_),
    .A2(_03310_),
    .B1(_03291_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand2_1 _15151_ (.A(_05476_),
    .B(_03311_),
    .Y(_00759_));
 sky130_fd_sc_hd__nand2_1 _15152_ (.A(_09350_),
    .B(_05458_),
    .Y(_03312_));
 sky130_fd_sc_hd__a21oi_1 _15153_ (.A1(_09350_),
    .A2(_03181_),
    .B1(_09352_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _15154_ (.A(_09348_),
    .B(_03199_),
    .Y(_03314_));
 sky130_fd_sc_hd__o21ai_0 _15155_ (.A1(_03177_),
    .A2(_03313_),
    .B1(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand2_1 _15156_ (.A(_05472_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__o22ai_1 _15157_ (.A1(_03183_),
    .A2(_03286_),
    .B1(_03261_),
    .B2(_03270_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _15158_ (.A1(_05458_),
    .A2(_03317_),
    .B1(_03250_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2_1 _15159_ (.A(_09352_),
    .B(_03181_),
    .Y(_03319_));
 sky130_fd_sc_hd__o2111a_1 _15160_ (.A1(_03179_),
    .A2(_03312_),
    .B1(_03316_),
    .C1(_03318_),
    .D1(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__o21ai_0 _15161_ (.A1(_02916_),
    .A2(_03320_),
    .B1(_05476_),
    .Y(_00760_));
 sky130_fd_sc_hd__nor3_1 _15162_ (.A(_09350_),
    .B(_03181_),
    .C(_03179_),
    .Y(_03321_));
 sky130_fd_sc_hd__a21oi_1 _15163_ (.A1(_03181_),
    .A2(_03179_),
    .B1(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__nor2_1 _15164_ (.A(_03189_),
    .B(_05472_),
    .Y(_03323_));
 sky130_fd_sc_hd__a211o_1 _15165_ (.A1(_09352_),
    .A2(_03177_),
    .B1(_03323_),
    .C1(_09347_),
    .X(_03324_));
 sky130_fd_sc_hd__a21oi_1 _15166_ (.A1(_03322_),
    .A2(_03324_),
    .B1(_03285_),
    .Y(_03325_));
 sky130_fd_sc_hd__o21ai_0 _15167_ (.A1(_03176_),
    .A2(_03325_),
    .B1(_05476_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2_1 _15168_ (.A(_09352_),
    .B(_03263_),
    .Y(_03326_));
 sky130_fd_sc_hd__o21ai_0 _15169_ (.A1(_03172_),
    .A2(_03179_),
    .B1(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__a21oi_1 _15170_ (.A1(_09347_),
    .A2(_05458_),
    .B1(_09350_),
    .Y(_03328_));
 sky130_fd_sc_hd__nor2_1 _15171_ (.A(_03214_),
    .B(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__a21oi_1 _15172_ (.A1(_03181_),
    .A2(_03327_),
    .B1(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand2_1 _15173_ (.A(_09350_),
    .B(_03190_),
    .Y(_03331_));
 sky130_fd_sc_hd__nand2_1 _15174_ (.A(_03239_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand2_1 _15175_ (.A(_03181_),
    .B(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__nor2_1 _15176_ (.A(_09348_),
    .B(_09352_),
    .Y(_03334_));
 sky130_fd_sc_hd__nor2_1 _15177_ (.A(_03178_),
    .B(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__o21ai_0 _15178_ (.A1(_03323_),
    .A2(_03335_),
    .B1(_05461_),
    .Y(_03336_));
 sky130_fd_sc_hd__o21ai_0 _15179_ (.A1(_05472_),
    .A2(_03172_),
    .B1(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand2_1 _15180_ (.A(_09347_),
    .B(_03181_),
    .Y(_03338_));
 sky130_fd_sc_hd__o21ai_0 _15181_ (.A1(_03214_),
    .A2(_03338_),
    .B1(_03175_),
    .Y(_03339_));
 sky130_fd_sc_hd__a21oi_1 _15182_ (.A1(_05458_),
    .A2(_03337_),
    .B1(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__a31oi_1 _15183_ (.A1(_03330_),
    .A2(_03333_),
    .A3(_03340_),
    .B1(_05482_),
    .Y(_00762_));
 sky130_fd_sc_hd__nor2_1 _15184_ (.A(_05458_),
    .B(_05472_),
    .Y(_03341_));
 sky130_fd_sc_hd__a21oi_1 _15185_ (.A1(_09352_),
    .A2(_05472_),
    .B1(_03323_),
    .Y(_03342_));
 sky130_fd_sc_hd__o22ai_1 _15186_ (.A1(_03183_),
    .A2(_03341_),
    .B1(_03342_),
    .B2(_03181_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2_1 _15187_ (.A(_05461_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__a21oi_1 _15188_ (.A1(_09352_),
    .A2(_03178_),
    .B1(_09348_),
    .Y(_03345_));
 sky130_fd_sc_hd__nor2_1 _15189_ (.A(_05458_),
    .B(_03178_),
    .Y(_03346_));
 sky130_fd_sc_hd__o21ai_0 _15190_ (.A1(_03219_),
    .A2(_03346_),
    .B1(_09350_),
    .Y(_03347_));
 sky130_fd_sc_hd__o21a_1 _15191_ (.A1(_03194_),
    .A2(_03345_),
    .B1(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__a31oi_1 _15192_ (.A1(_03273_),
    .A2(_03344_),
    .A3(_03348_),
    .B1(_03176_),
    .Y(_00763_));
 sky130_fd_sc_hd__nor2_1 _15193_ (.A(_09348_),
    .B(_09350_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_1 _15194_ (.A(_05461_),
    .B(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__o311ai_0 _15195_ (.A1(_09347_),
    .A2(_09352_),
    .A3(_05461_),
    .B1(_03249_),
    .C1(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__o21ai_0 _15196_ (.A1(_03349_),
    .A2(_03179_),
    .B1(_03326_),
    .Y(_03352_));
 sky130_fd_sc_hd__or2_2 _15197_ (.A(_03346_),
    .B(_03249_),
    .X(_03353_));
 sky130_fd_sc_hd__o22ai_1 _15198_ (.A1(_05458_),
    .A2(_03172_),
    .B1(_03174_),
    .B2(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__a22oi_1 _15199_ (.A1(_03181_),
    .A2(_03352_),
    .B1(_03354_),
    .B2(_05461_),
    .Y(_03355_));
 sky130_fd_sc_hd__and3_1 _15200_ (.A(_03248_),
    .B(_03351_),
    .C(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__o21ai_0 _15201_ (.A1(_03176_),
    .A2(_03356_),
    .B1(_05476_),
    .Y(_00764_));
 sky130_fd_sc_hd__a21oi_1 _15202_ (.A1(_09350_),
    .A2(_03181_),
    .B1(_09348_),
    .Y(_03357_));
 sky130_fd_sc_hd__nor2_1 _15203_ (.A(_03177_),
    .B(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__a21oi_1 _15204_ (.A1(_09347_),
    .A2(_03199_),
    .B1(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__nor2_1 _15205_ (.A(_03288_),
    .B(_03334_),
    .Y(_03360_));
 sky130_fd_sc_hd__nor2_1 _15206_ (.A(_03323_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__o221a_2 _15207_ (.A1(_03178_),
    .A2(_03359_),
    .B1(_03361_),
    .B2(_05461_),
    .C1(_03309_),
    .X(_03362_));
 sky130_fd_sc_hd__o21ai_0 _15208_ (.A1(_03176_),
    .A2(_03362_),
    .B1(_05476_),
    .Y(_00765_));
 sky130_fd_sc_hd__o21ai_0 _15209_ (.A1(_09348_),
    .A2(_03214_),
    .B1(_03179_),
    .Y(_03363_));
 sky130_fd_sc_hd__and3_1 _15210_ (.A(_03183_),
    .B(_05458_),
    .C(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__a21oi_1 _15211_ (.A1(_09347_),
    .A2(_05458_),
    .B1(_09348_),
    .Y(_03365_));
 sky130_fd_sc_hd__nor2_1 _15212_ (.A(_03241_),
    .B(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__a21oi_1 _15213_ (.A1(_03281_),
    .A2(_03366_),
    .B1(_09350_),
    .Y(_03367_));
 sky130_fd_sc_hd__nor3_1 _15214_ (.A(_03176_),
    .B(_03364_),
    .C(_03367_),
    .Y(_00766_));
 sky130_fd_sc_hd__nor2_1 _15215_ (.A(_03238_),
    .B(_03312_),
    .Y(_03368_));
 sky130_fd_sc_hd__nor3_1 _15216_ (.A(_05458_),
    .B(_03263_),
    .C(_03307_),
    .Y(_03369_));
 sky130_fd_sc_hd__nor2_1 _15217_ (.A(_03346_),
    .B(_03249_),
    .Y(_03370_));
 sky130_fd_sc_hd__nand2_1 _15218_ (.A(_09352_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_1 _15219_ (.A(_09348_),
    .B(_03341_),
    .Y(_03372_));
 sky130_fd_sc_hd__a21oi_1 _15220_ (.A1(_03371_),
    .A2(_03372_),
    .B1(_05461_),
    .Y(_03373_));
 sky130_fd_sc_hd__nor3_1 _15221_ (.A(_03368_),
    .B(_03369_),
    .C(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__a21oi_1 _15222_ (.A1(_03318_),
    .A2(_03374_),
    .B1(_05482_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2_1 _15223_ (.A(_03274_),
    .B(_03246_),
    .Y(_03375_));
 sky130_fd_sc_hd__a31oi_1 _15224_ (.A1(_03177_),
    .A2(_03319_),
    .A3(_03312_),
    .B1(_05472_),
    .Y(_03376_));
 sky130_fd_sc_hd__o21ai_0 _15225_ (.A1(_09348_),
    .A2(_03375_),
    .B1(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__o21ai_0 _15226_ (.A1(_03237_),
    .A2(_03249_),
    .B1(_09347_),
    .Y(_03378_));
 sky130_fd_sc_hd__nand2_1 _15227_ (.A(_03377_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__nand2_1 _15228_ (.A(_03291_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_1 _15229_ (.A(_05476_),
    .B(_03380_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_09352_),
    .B(_03249_),
    .Y(_03381_));
 sky130_fd_sc_hd__nor2_1 _15231_ (.A(_03178_),
    .B(_03307_),
    .Y(_03382_));
 sky130_fd_sc_hd__o21ai_0 _15232_ (.A1(_09348_),
    .A2(_03382_),
    .B1(_03181_),
    .Y(_03383_));
 sky130_fd_sc_hd__a21oi_1 _15233_ (.A1(_03381_),
    .A2(_03383_),
    .B1(_03177_),
    .Y(_03384_));
 sky130_fd_sc_hd__o21ai_0 _15234_ (.A1(_09350_),
    .A2(_03177_),
    .B1(_05472_),
    .Y(_03385_));
 sky130_fd_sc_hd__o211ai_1 _15235_ (.A1(_09348_),
    .A2(_03286_),
    .B1(_03261_),
    .C1(_05458_),
    .Y(_03386_));
 sky130_fd_sc_hd__a21oi_1 _15236_ (.A1(_03183_),
    .A2(_03385_),
    .B1(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a2111oi_0 _15237_ (.A1(_03181_),
    .A2(_03352_),
    .B1(_03384_),
    .C1(_03387_),
    .D1(_03282_),
    .Y(_03388_));
 sky130_fd_sc_hd__nor2_1 _15238_ (.A(_05482_),
    .B(_03388_),
    .Y(_00769_));
 sky130_fd_sc_hd__o22ai_1 _15239_ (.A1(_03349_),
    .A2(_03179_),
    .B1(_03237_),
    .B2(_03183_),
    .Y(_03389_));
 sky130_fd_sc_hd__nand2_1 _15240_ (.A(_05458_),
    .B(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__a31oi_1 _15241_ (.A1(_03248_),
    .A2(_03330_),
    .A3(_03390_),
    .B1(_03176_),
    .Y(_00770_));
 sky130_fd_sc_hd__o21ai_0 _15242_ (.A1(_05458_),
    .A2(_03261_),
    .B1(_03199_),
    .Y(_03391_));
 sky130_fd_sc_hd__a222oi_1 _15243_ (.A1(_09350_),
    .A2(_03341_),
    .B1(_03261_),
    .B2(_09352_),
    .C1(_03391_),
    .C2(_09347_),
    .Y(_03392_));
 sky130_fd_sc_hd__a21oi_1 _15244_ (.A1(_03333_),
    .A2(_03392_),
    .B1(_03176_),
    .Y(_00771_));
 sky130_fd_sc_hd__a21oi_1 _15245_ (.A1(_09347_),
    .A2(_03181_),
    .B1(_09352_),
    .Y(_03393_));
 sky130_fd_sc_hd__o21ai_0 _15246_ (.A1(_05461_),
    .A2(_03393_),
    .B1(_03275_),
    .Y(_03394_));
 sky130_fd_sc_hd__nor2_1 _15247_ (.A(_03178_),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__a221oi_1 _15248_ (.A1(_09350_),
    .A2(_03195_),
    .B1(_03293_),
    .B2(_09352_),
    .C1(_05472_),
    .Y(_03396_));
 sky130_fd_sc_hd__o21ai_0 _15249_ (.A1(_03395_),
    .A2(_03396_),
    .B1(_03235_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _15250_ (.A(_03291_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_1 _15251_ (.A(_05476_),
    .B(_03398_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand3_1 _15252_ (.A(_03189_),
    .B(_05472_),
    .C(_03194_),
    .Y(_03399_));
 sky130_fd_sc_hd__a21oi_1 _15253_ (.A1(_03193_),
    .A2(_03399_),
    .B1(_09352_),
    .Y(_03400_));
 sky130_fd_sc_hd__a21oi_1 _15254_ (.A1(_09348_),
    .A2(_03181_),
    .B1(_09352_),
    .Y(_03401_));
 sky130_fd_sc_hd__nor2_1 _15255_ (.A(_09348_),
    .B(_03281_),
    .Y(_03402_));
 sky130_fd_sc_hd__a21oi_1 _15256_ (.A1(_03178_),
    .A2(_03401_),
    .B1(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__o221ai_1 _15257_ (.A1(_03181_),
    .A2(_03261_),
    .B1(_03403_),
    .B2(_09347_),
    .C1(_03291_),
    .Y(_03404_));
 sky130_fd_sc_hd__o21ai_0 _15258_ (.A1(_03400_),
    .A2(_03404_),
    .B1(_05476_),
    .Y(_00773_));
 sky130_fd_sc_hd__a21oi_1 _15259_ (.A1(_03312_),
    .A2(_03338_),
    .B1(_05472_),
    .Y(_03405_));
 sky130_fd_sc_hd__a21oi_1 _15260_ (.A1(_09348_),
    .A2(_03260_),
    .B1(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__nor2_1 _15261_ (.A(_03177_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__a21oi_1 _15262_ (.A1(_03338_),
    .A2(_03371_),
    .B1(_05461_),
    .Y(_03408_));
 sky130_fd_sc_hd__nor3_1 _15263_ (.A(_03303_),
    .B(_03407_),
    .C(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__nor2_1 _15264_ (.A(_03176_),
    .B(_03409_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _15265_ (.A(_09348_),
    .B(_03178_),
    .Y(_03410_));
 sky130_fd_sc_hd__a21oi_1 _15266_ (.A1(_09350_),
    .A2(_05472_),
    .B1(_09347_),
    .Y(_03411_));
 sky130_fd_sc_hd__a21oi_1 _15267_ (.A1(_03410_),
    .A2(_03411_),
    .B1(_03193_),
    .Y(_03412_));
 sky130_fd_sc_hd__nor2_1 _15268_ (.A(_03339_),
    .B(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__and3_1 _15269_ (.A(_03309_),
    .B(_03348_),
    .C(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__o21ai_0 _15270_ (.A1(_02916_),
    .A2(_03414_),
    .B1(_05476_),
    .Y(_00775_));
 sky130_fd_sc_hd__o21ai_0 _15271_ (.A1(_05461_),
    .A2(_03172_),
    .B1(_03189_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_1 _15272_ (.A(_03288_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__o21ai_0 _15273_ (.A1(_03177_),
    .A2(_03260_),
    .B1(_03179_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _15274_ (.A(_09347_),
    .B(_03263_),
    .Y(_03418_));
 sky130_fd_sc_hd__a21oi_1 _15275_ (.A1(_03297_),
    .A2(_03418_),
    .B1(_03181_),
    .Y(_03419_));
 sky130_fd_sc_hd__a211oi_1 _15276_ (.A1(_09352_),
    .A2(_03417_),
    .B1(_03419_),
    .C1(_03407_),
    .Y(_03420_));
 sky130_fd_sc_hd__a21oi_1 _15277_ (.A1(_03416_),
    .A2(_03420_),
    .B1(_03176_),
    .Y(_00776_));
 sky130_fd_sc_hd__nor2_1 _15278_ (.A(_03274_),
    .B(_03328_),
    .Y(_03421_));
 sky130_fd_sc_hd__o211ai_1 _15279_ (.A1(_09352_),
    .A2(_03421_),
    .B1(_03194_),
    .C1(_05472_),
    .Y(_03422_));
 sky130_fd_sc_hd__nor2_1 _15280_ (.A(_03282_),
    .B(_03296_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21oi_1 _15281_ (.A1(_03422_),
    .A2(_03423_),
    .B1(_05482_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _15282_ (.A(_09347_),
    .B(_05472_),
    .Y(_03424_));
 sky130_fd_sc_hd__a21oi_1 _15283_ (.A1(_03174_),
    .A2(_03424_),
    .B1(_03177_),
    .Y(_03425_));
 sky130_fd_sc_hd__a21oi_1 _15284_ (.A1(_09348_),
    .A2(_03178_),
    .B1(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _15285_ (.A(_03193_),
    .B(_03286_),
    .Y(_03427_));
 sky130_fd_sc_hd__o22ai_1 _15286_ (.A1(_03261_),
    .A2(_03312_),
    .B1(_03338_),
    .B2(_03286_),
    .Y(_03428_));
 sky130_fd_sc_hd__a21oi_1 _15287_ (.A1(_09348_),
    .A2(_03427_),
    .B1(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__o21ai_0 _15288_ (.A1(_05458_),
    .A2(_03426_),
    .B1(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__o21ai_0 _15289_ (.A1(_03250_),
    .A2(_03430_),
    .B1(_05481_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _15290_ (.A(_05476_),
    .B(_03431_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _15291_ (.A(_09352_),
    .B(_03288_),
    .Y(_03432_));
 sky130_fd_sc_hd__o21ai_0 _15292_ (.A1(_03189_),
    .A2(_03353_),
    .B1(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__o22ai_1 _15293_ (.A1(_03233_),
    .A2(_03307_),
    .B1(_03334_),
    .B2(_03199_),
    .Y(_03434_));
 sky130_fd_sc_hd__a21oi_1 _15294_ (.A1(_03319_),
    .A2(_03328_),
    .B1(_03214_),
    .Y(_03435_));
 sky130_fd_sc_hd__a221oi_1 _15295_ (.A1(_03177_),
    .A2(_03433_),
    .B1(_03434_),
    .B2(_03178_),
    .C1(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21oi_1 _15296_ (.A1(_03429_),
    .A2(_03436_),
    .B1(_03176_),
    .Y(_00779_));
 sky130_fd_sc_hd__o21ai_0 _15297_ (.A1(_09352_),
    .A2(_03178_),
    .B1(_05458_),
    .Y(_03437_));
 sky130_fd_sc_hd__o22ai_1 _15298_ (.A1(_09352_),
    .A2(_03193_),
    .B1(_03179_),
    .B2(_05458_),
    .Y(_03438_));
 sky130_fd_sc_hd__a21oi_1 _15299_ (.A1(_03189_),
    .A2(_03437_),
    .B1(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__o22ai_1 _15300_ (.A1(_03177_),
    .A2(_03370_),
    .B1(_03439_),
    .B2(_09348_),
    .Y(_03440_));
 sky130_fd_sc_hd__a21oi_1 _15301_ (.A1(_03277_),
    .A2(_03440_),
    .B1(_03176_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand2_1 _15302_ (.A(_09348_),
    .B(_03190_),
    .Y(_03441_));
 sky130_fd_sc_hd__a21oi_1 _15303_ (.A1(_03441_),
    .A2(_03418_),
    .B1(_03181_),
    .Y(_03442_));
 sky130_fd_sc_hd__a21oi_1 _15304_ (.A1(_09350_),
    .A2(_05472_),
    .B1(_03181_),
    .Y(_03443_));
 sky130_fd_sc_hd__nor2_1 _15305_ (.A(_03178_),
    .B(_03182_),
    .Y(_03444_));
 sky130_fd_sc_hd__nor3_1 _15306_ (.A(_05461_),
    .B(_03443_),
    .C(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__o21ai_0 _15307_ (.A1(_05458_),
    .A2(_03334_),
    .B1(_03183_),
    .Y(_03446_));
 sky130_fd_sc_hd__o21ai_0 _15308_ (.A1(_09348_),
    .A2(_03178_),
    .B1(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__a211oi_1 _15309_ (.A1(_03189_),
    .A2(_03447_),
    .B1(_03288_),
    .C1(_03177_),
    .Y(_03448_));
 sky130_fd_sc_hd__or4_1 _15310_ (.A(_03250_),
    .B(_03442_),
    .C(_03445_),
    .D(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__a21o_1 _15311_ (.A1(_05481_),
    .A2(_03449_),
    .B1(reset_hash),
    .X(_00781_));
 sky130_fd_sc_hd__o21ai_0 _15312_ (.A1(_03237_),
    .A2(_03341_),
    .B1(_09347_),
    .Y(_03450_));
 sky130_fd_sc_hd__nor3_1 _15313_ (.A(_09347_),
    .B(_09348_),
    .C(_09352_),
    .Y(_03451_));
 sky130_fd_sc_hd__nor2_1 _15314_ (.A(_03341_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__a21oi_1 _15315_ (.A1(_05472_),
    .A2(_03319_),
    .B1(_03177_),
    .Y(_03453_));
 sky130_fd_sc_hd__o21ai_0 _15316_ (.A1(_09350_),
    .A2(_03452_),
    .B1(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__a21oi_1 _15317_ (.A1(_03307_),
    .A2(_03249_),
    .B1(_03346_),
    .Y(_03455_));
 sky130_fd_sc_hd__o221ai_1 _15318_ (.A1(_09352_),
    .A2(_03353_),
    .B1(_03455_),
    .B2(_09348_),
    .C1(_03177_),
    .Y(_03456_));
 sky130_fd_sc_hd__a41oi_1 _15319_ (.A1(_03175_),
    .A2(_03450_),
    .A3(_03454_),
    .A4(_03456_),
    .B1(_05482_),
    .Y(_00782_));
 sky130_fd_sc_hd__o21ai_0 _15320_ (.A1(_05458_),
    .A2(_03219_),
    .B1(_09352_),
    .Y(_03457_));
 sky130_fd_sc_hd__a21oi_1 _15321_ (.A1(_03288_),
    .A2(_03278_),
    .B1(_03250_),
    .Y(_03458_));
 sky130_fd_sc_hd__a221o_1 _15322_ (.A1(_09347_),
    .A2(_03195_),
    .B1(_03293_),
    .B2(_09348_),
    .C1(_05472_),
    .X(_03459_));
 sky130_fd_sc_hd__a21oi_1 _15323_ (.A1(_09348_),
    .A2(_03177_),
    .B1(_09350_),
    .Y(_03460_));
 sky130_fd_sc_hd__o21ai_0 _15324_ (.A1(_03272_),
    .A2(_03460_),
    .B1(_05472_),
    .Y(_03461_));
 sky130_fd_sc_hd__nand2_1 _15325_ (.A(_03459_),
    .B(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__a31oi_1 _15326_ (.A1(_03457_),
    .A2(_03458_),
    .A3(_03462_),
    .B1(_05482_),
    .Y(_00783_));
 sky130_fd_sc_hd__nor2_1 _15327_ (.A(reset_hash),
    .B(_02845_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_1 _15329_ (.A(_05350_),
    .B(_07566_),
    .Y(_03464_));
 sky130_fd_sc_hd__nor2_1 _15331_ (.A(_07572_),
    .B(_03464_),
    .Y(_00785_));
 sky130_fd_sc_hd__nor2_1 _15333_ (.A(_07660_),
    .B(_03464_),
    .Y(_00786_));
 sky130_fd_sc_hd__nor2_1 _15335_ (.A(_07669_),
    .B(_03464_),
    .Y(_00787_));
 sky130_fd_sc_hd__nor2_1 _15337_ (.A(_07677_),
    .B(_03464_),
    .Y(_00788_));
 sky130_fd_sc_hd__nor2_1 _15339_ (.A(_07689_),
    .B(_03464_),
    .Y(_00789_));
 sky130_fd_sc_hd__nor2_1 _15341_ (.A(_07703_),
    .B(_03464_),
    .Y(_00790_));
 sky130_fd_sc_hd__nor2_1 _15343_ (.A(_07709_),
    .B(_03464_),
    .Y(_00791_));
 sky130_fd_sc_hd__nor2_1 _15345_ (.A(_07715_),
    .B(_03464_),
    .Y(_00792_));
 sky130_fd_sc_hd__nor2_1 _15347_ (.A(_07731_),
    .B(_03464_),
    .Y(_00793_));
 sky130_fd_sc_hd__nor2_1 _15349_ (.A(_07745_),
    .B(_03464_),
    .Y(_00794_));
 sky130_fd_sc_hd__nor2_1 _15352_ (.A(_07752_),
    .B(_03464_),
    .Y(_00795_));
 sky130_fd_sc_hd__nor2_1 _15354_ (.A(_07577_),
    .B(_03464_),
    .Y(_00796_));
 sky130_fd_sc_hd__nor2_1 _15356_ (.A(_07766_),
    .B(_03464_),
    .Y(_00797_));
 sky130_fd_sc_hd__nor2_1 _15358_ (.A(_07777_),
    .B(_03464_),
    .Y(_00798_));
 sky130_fd_sc_hd__nor2_1 _15360_ (.A(_07786_),
    .B(_03464_),
    .Y(_00799_));
 sky130_fd_sc_hd__nor2_1 _15362_ (.A(_07800_),
    .B(_03464_),
    .Y(_00800_));
 sky130_fd_sc_hd__nor2_1 _15364_ (.A(_07809_),
    .B(_03464_),
    .Y(_00801_));
 sky130_fd_sc_hd__nor2_1 _15366_ (.A(_07818_),
    .B(_03464_),
    .Y(_00802_));
 sky130_fd_sc_hd__nor2_1 _15368_ (.A(_07831_),
    .B(_03464_),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_1 _15370_ (.A(_07843_),
    .B(_03464_),
    .Y(_00804_));
 sky130_fd_sc_hd__nor2_1 _15373_ (.A(_07850_),
    .B(_03464_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand4_1 _15374_ (.A(_07852_),
    .B(_07856_),
    .C(_07857_),
    .D(_07853_),
    .Y(_03488_));
 sky130_fd_sc_hd__a31o_2 _15375_ (.A1(_07856_),
    .A2(_07857_),
    .A3(_07853_),
    .B1(_07852_),
    .X(_03489_));
 sky130_fd_sc_hd__and2_1 _15376_ (.A(\w[62][29] ),
    .B(done),
    .X(_03490_));
 sky130_fd_sc_hd__a31oi_1 _15377_ (.A1(_07591_),
    .A2(_03488_),
    .A3(_03489_),
    .B1(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__nor2_1 _15379_ (.A(_03464_),
    .B(_03491_),
    .Y(_00806_));
 sky130_fd_sc_hd__nor2_1 _15381_ (.A(_07581_),
    .B(_03464_),
    .Y(_00807_));
 sky130_fd_sc_hd__nor2_1 _15383_ (.A(_07873_),
    .B(_03464_),
    .Y(_00808_));
 sky130_fd_sc_hd__nor2_1 _15385_ (.A(_07925_),
    .B(_03464_),
    .Y(_00809_));
 sky130_fd_sc_hd__nor2_1 _15387_ (.A(_07588_),
    .B(_03464_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor2_1 _15389_ (.A(_07601_),
    .B(_03464_),
    .Y(_00811_));
 sky130_fd_sc_hd__nor2_1 _15391_ (.A(_07610_),
    .B(_03464_),
    .Y(_00812_));
 sky130_fd_sc_hd__nor2_1 _15393_ (.A(_07620_),
    .B(_03464_),
    .Y(_00813_));
 sky130_fd_sc_hd__nor2_1 _15395_ (.A(_07628_),
    .B(_03464_),
    .Y(_00814_));
 sky130_fd_sc_hd__nor2_1 _15397_ (.A(_07635_),
    .B(_03464_),
    .Y(_00815_));
 sky130_fd_sc_hd__nor2_1 _15399_ (.A(_07646_),
    .B(_03464_),
    .Y(_00816_));
 sky130_fd_sc_hd__nand2_1 _15401_ (.A(_05400_),
    .B(_07927_),
    .Y(_03504_));
 sky130_fd_sc_hd__nor2_1 _15403_ (.A(_07930_),
    .B(_03504_),
    .Y(_00817_));
 sky130_fd_sc_hd__nor2_1 _15405_ (.A(_08006_),
    .B(_03504_),
    .Y(_00818_));
 sky130_fd_sc_hd__nor2_1 _15407_ (.A(_08018_),
    .B(_03504_),
    .Y(_00819_));
 sky130_fd_sc_hd__nor2_1 _15409_ (.A(_08025_),
    .B(_03504_),
    .Y(_00820_));
 sky130_fd_sc_hd__nor2_1 _15411_ (.A(_08031_),
    .B(_03504_),
    .Y(_00821_));
 sky130_fd_sc_hd__nor2_1 _15413_ (.A(_08039_),
    .B(_03504_),
    .Y(_00822_));
 sky130_fd_sc_hd__nor2_1 _15415_ (.A(_08051_),
    .B(_03504_),
    .Y(_00823_));
 sky130_fd_sc_hd__nor2_1 _15417_ (.A(_08064_),
    .B(_03504_),
    .Y(_00824_));
 sky130_fd_sc_hd__nor2_1 _15419_ (.A(_08071_),
    .B(_03504_),
    .Y(_00825_));
 sky130_fd_sc_hd__nor2_1 _15421_ (.A(_08082_),
    .B(_03504_),
    .Y(_00826_));
 sky130_fd_sc_hd__nor2_1 _15424_ (.A(_08091_),
    .B(_03504_),
    .Y(_00827_));
 sky130_fd_sc_hd__nor2_1 _15426_ (.A(_07934_),
    .B(_03504_),
    .Y(_00828_));
 sky130_fd_sc_hd__nor2_1 _15428_ (.A(_08102_),
    .B(_03504_),
    .Y(_00829_));
 sky130_fd_sc_hd__nor2_1 _15430_ (.A(_08114_),
    .B(_03504_),
    .Y(_00830_));
 sky130_fd_sc_hd__nor2_1 _15432_ (.A(_08125_),
    .B(_03504_),
    .Y(_00831_));
 sky130_fd_sc_hd__nor2_1 _15434_ (.A(_08142_),
    .B(_03504_),
    .Y(_00832_));
 sky130_fd_sc_hd__nor2_1 _15436_ (.A(_08152_),
    .B(_03504_),
    .Y(_00833_));
 sky130_fd_sc_hd__nor2_1 _15438_ (.A(_08160_),
    .B(_03504_),
    .Y(_00834_));
 sky130_fd_sc_hd__nor2_1 _15440_ (.A(_08171_),
    .B(_03504_),
    .Y(_00835_));
 sky130_fd_sc_hd__nor2_1 _15442_ (.A(_08184_),
    .B(_03504_),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2_1 _15445_ (.A(_08204_),
    .B(_03504_),
    .Y(_00837_));
 sky130_fd_sc_hd__nor2_1 _15447_ (.A(_08209_),
    .B(_03504_),
    .Y(_00838_));
 sky130_fd_sc_hd__nor2_1 _15449_ (.A(_07937_),
    .B(_03504_),
    .Y(_00839_));
 sky130_fd_sc_hd__nor2_1 _15451_ (.A(_08221_),
    .B(_03504_),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2_1 _15453_ (.A(_08254_),
    .B(_03504_),
    .Y(_00841_));
 sky130_fd_sc_hd__nor2_1 _15455_ (.A(_07942_),
    .B(_03504_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2_1 _15457_ (.A(_07949_),
    .B(_03504_),
    .Y(_00843_));
 sky130_fd_sc_hd__nor2_1 _15459_ (.A(_07956_),
    .B(_03504_),
    .Y(_00844_));
 sky130_fd_sc_hd__nor2_1 _15461_ (.A(_07965_),
    .B(_03504_),
    .Y(_00845_));
 sky130_fd_sc_hd__nor2_1 _15463_ (.A(_07974_),
    .B(_03504_),
    .Y(_00846_));
 sky130_fd_sc_hd__nor2_1 _15465_ (.A(_07981_),
    .B(_03504_),
    .Y(_00847_));
 sky130_fd_sc_hd__nor2_1 _15467_ (.A(_07989_),
    .B(_03504_),
    .Y(_00848_));
 sky130_fd_sc_hd__nand2_1 _15468_ (.A(_05350_),
    .B(_08257_),
    .Y(_03539_));
 sky130_fd_sc_hd__nor2_1 _15470_ (.A(_07572_),
    .B(_03539_),
    .Y(_00849_));
 sky130_fd_sc_hd__nor2_1 _15471_ (.A(_07660_),
    .B(_03539_),
    .Y(_00850_));
 sky130_fd_sc_hd__nor2_1 _15472_ (.A(_07669_),
    .B(_03539_),
    .Y(_00851_));
 sky130_fd_sc_hd__nor2_1 _15473_ (.A(_07677_),
    .B(_03539_),
    .Y(_00852_));
 sky130_fd_sc_hd__nor2_1 _15474_ (.A(_07689_),
    .B(_03539_),
    .Y(_00853_));
 sky130_fd_sc_hd__nor2_1 _15475_ (.A(_07703_),
    .B(_03539_),
    .Y(_00854_));
 sky130_fd_sc_hd__nor2_1 _15476_ (.A(_07709_),
    .B(_03539_),
    .Y(_00855_));
 sky130_fd_sc_hd__nor2_1 _15477_ (.A(_07715_),
    .B(_03539_),
    .Y(_00856_));
 sky130_fd_sc_hd__nor2_1 _15478_ (.A(_07731_),
    .B(_03539_),
    .Y(_00857_));
 sky130_fd_sc_hd__nor2_1 _15479_ (.A(_07745_),
    .B(_03539_),
    .Y(_00858_));
 sky130_fd_sc_hd__nor2_1 _15481_ (.A(_07752_),
    .B(_03539_),
    .Y(_00859_));
 sky130_fd_sc_hd__nor2_1 _15482_ (.A(_07577_),
    .B(_03539_),
    .Y(_00860_));
 sky130_fd_sc_hd__nor2_1 _15483_ (.A(_07766_),
    .B(_03539_),
    .Y(_00861_));
 sky130_fd_sc_hd__nor2_1 _15484_ (.A(_07777_),
    .B(_03539_),
    .Y(_00862_));
 sky130_fd_sc_hd__nor2_1 _15485_ (.A(_07786_),
    .B(_03539_),
    .Y(_00863_));
 sky130_fd_sc_hd__nor2_1 _15486_ (.A(_07800_),
    .B(_03539_),
    .Y(_00864_));
 sky130_fd_sc_hd__nor2_1 _15487_ (.A(_07809_),
    .B(_03539_),
    .Y(_00865_));
 sky130_fd_sc_hd__nor2_1 _15488_ (.A(_07818_),
    .B(_03539_),
    .Y(_00866_));
 sky130_fd_sc_hd__nor2_1 _15489_ (.A(_07831_),
    .B(_03539_),
    .Y(_00867_));
 sky130_fd_sc_hd__nor2_1 _15490_ (.A(_07843_),
    .B(_03539_),
    .Y(_00868_));
 sky130_fd_sc_hd__nor2_1 _15492_ (.A(_07850_),
    .B(_03539_),
    .Y(_00869_));
 sky130_fd_sc_hd__nor2_1 _15493_ (.A(_03491_),
    .B(_03539_),
    .Y(_00870_));
 sky130_fd_sc_hd__nor2_1 _15494_ (.A(_07581_),
    .B(_03539_),
    .Y(_00871_));
 sky130_fd_sc_hd__nor2_1 _15495_ (.A(_07873_),
    .B(_03539_),
    .Y(_00872_));
 sky130_fd_sc_hd__nor2_1 _15496_ (.A(_07925_),
    .B(_03539_),
    .Y(_00873_));
 sky130_fd_sc_hd__nor2_1 _15497_ (.A(_07588_),
    .B(_03539_),
    .Y(_00874_));
 sky130_fd_sc_hd__nor2_1 _15498_ (.A(_07601_),
    .B(_03539_),
    .Y(_00875_));
 sky130_fd_sc_hd__nor2_1 _15499_ (.A(_07610_),
    .B(_03539_),
    .Y(_00876_));
 sky130_fd_sc_hd__nor2_1 _15500_ (.A(_07620_),
    .B(_03539_),
    .Y(_00877_));
 sky130_fd_sc_hd__nor2_1 _15501_ (.A(_07628_),
    .B(_03539_),
    .Y(_00878_));
 sky130_fd_sc_hd__nor2_1 _15502_ (.A(_07635_),
    .B(_03539_),
    .Y(_00879_));
 sky130_fd_sc_hd__nor2_1 _15503_ (.A(_07646_),
    .B(_03539_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_1 _15504_ (.A(_05400_),
    .B(_08304_),
    .Y(_03543_));
 sky130_fd_sc_hd__nor2_1 _15506_ (.A(_07930_),
    .B(_03543_),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2_1 _15507_ (.A(_08006_),
    .B(_03543_),
    .Y(_00882_));
 sky130_fd_sc_hd__nor2_1 _15508_ (.A(_08018_),
    .B(_03543_),
    .Y(_00883_));
 sky130_fd_sc_hd__nor2_1 _15509_ (.A(_08025_),
    .B(_03543_),
    .Y(_00884_));
 sky130_fd_sc_hd__nor2_1 _15510_ (.A(_08031_),
    .B(_03543_),
    .Y(_00885_));
 sky130_fd_sc_hd__nor2_1 _15511_ (.A(_08039_),
    .B(_03543_),
    .Y(_00886_));
 sky130_fd_sc_hd__nor2_1 _15512_ (.A(_08051_),
    .B(_03543_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_1 _15513_ (.A(_08064_),
    .B(_03543_),
    .Y(_00888_));
 sky130_fd_sc_hd__nor2_1 _15514_ (.A(_08071_),
    .B(_03543_),
    .Y(_00889_));
 sky130_fd_sc_hd__nor2_1 _15515_ (.A(_08082_),
    .B(_03543_),
    .Y(_00890_));
 sky130_fd_sc_hd__nor2_1 _15517_ (.A(_08091_),
    .B(_03543_),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2_1 _15518_ (.A(_07934_),
    .B(_03543_),
    .Y(_00892_));
 sky130_fd_sc_hd__nor2_1 _15519_ (.A(_08102_),
    .B(_03543_),
    .Y(_00893_));
 sky130_fd_sc_hd__nor2_1 _15520_ (.A(_08114_),
    .B(_03543_),
    .Y(_00894_));
 sky130_fd_sc_hd__nor2_1 _15521_ (.A(_08125_),
    .B(_03543_),
    .Y(_00895_));
 sky130_fd_sc_hd__nor2_1 _15522_ (.A(_08142_),
    .B(_03543_),
    .Y(_00896_));
 sky130_fd_sc_hd__nor2_1 _15523_ (.A(_08152_),
    .B(_03543_),
    .Y(_00897_));
 sky130_fd_sc_hd__nor2_1 _15524_ (.A(_08160_),
    .B(_03543_),
    .Y(_00898_));
 sky130_fd_sc_hd__nor2_1 _15525_ (.A(_08171_),
    .B(_03543_),
    .Y(_00899_));
 sky130_fd_sc_hd__nor2_1 _15526_ (.A(_08184_),
    .B(_03543_),
    .Y(_00900_));
 sky130_fd_sc_hd__nor2_1 _15528_ (.A(_08204_),
    .B(_03543_),
    .Y(_00901_));
 sky130_fd_sc_hd__nor2_1 _15529_ (.A(_08209_),
    .B(_03543_),
    .Y(_00902_));
 sky130_fd_sc_hd__nor2_1 _15530_ (.A(_07937_),
    .B(_03543_),
    .Y(_00903_));
 sky130_fd_sc_hd__nor2_1 _15531_ (.A(_08221_),
    .B(_03543_),
    .Y(_00904_));
 sky130_fd_sc_hd__nor2_1 _15532_ (.A(_08254_),
    .B(_03543_),
    .Y(_00905_));
 sky130_fd_sc_hd__nor2_1 _15533_ (.A(_07942_),
    .B(_03543_),
    .Y(_00906_));
 sky130_fd_sc_hd__nor2_1 _15534_ (.A(_07949_),
    .B(_03543_),
    .Y(_00907_));
 sky130_fd_sc_hd__nor2_1 _15535_ (.A(_07956_),
    .B(_03543_),
    .Y(_00908_));
 sky130_fd_sc_hd__nor2_1 _15536_ (.A(_07965_),
    .B(_03543_),
    .Y(_00909_));
 sky130_fd_sc_hd__nor2_1 _15537_ (.A(_07974_),
    .B(_03543_),
    .Y(_00910_));
 sky130_fd_sc_hd__nor2_1 _15538_ (.A(_07981_),
    .B(_03543_),
    .Y(_00911_));
 sky130_fd_sc_hd__nor2_1 _15539_ (.A(_07989_),
    .B(_03543_),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_1 _15540_ (.A(_05350_),
    .B(_08346_),
    .Y(_03547_));
 sky130_fd_sc_hd__nor2_1 _15542_ (.A(_07572_),
    .B(_03547_),
    .Y(_00913_));
 sky130_fd_sc_hd__nor2_1 _15543_ (.A(_07660_),
    .B(_03547_),
    .Y(_00914_));
 sky130_fd_sc_hd__nor2_1 _15544_ (.A(_07669_),
    .B(_03547_),
    .Y(_00915_));
 sky130_fd_sc_hd__nor2_1 _15545_ (.A(_07677_),
    .B(_03547_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_1 _15546_ (.A(_07689_),
    .B(_03547_),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2_1 _15547_ (.A(_07703_),
    .B(_03547_),
    .Y(_00918_));
 sky130_fd_sc_hd__nor2_1 _15548_ (.A(_07709_),
    .B(_03547_),
    .Y(_00919_));
 sky130_fd_sc_hd__nor2_1 _15549_ (.A(_07715_),
    .B(_03547_),
    .Y(_00920_));
 sky130_fd_sc_hd__nor2_1 _15550_ (.A(_07731_),
    .B(_03547_),
    .Y(_00921_));
 sky130_fd_sc_hd__nor2_1 _15551_ (.A(_07745_),
    .B(_03547_),
    .Y(_00922_));
 sky130_fd_sc_hd__nor2_1 _15553_ (.A(_07752_),
    .B(_03547_),
    .Y(_00923_));
 sky130_fd_sc_hd__nor2_1 _15554_ (.A(_07577_),
    .B(_03547_),
    .Y(_00924_));
 sky130_fd_sc_hd__nor2_1 _15555_ (.A(_07766_),
    .B(_03547_),
    .Y(_00925_));
 sky130_fd_sc_hd__nor2_1 _15556_ (.A(_07777_),
    .B(_03547_),
    .Y(_00926_));
 sky130_fd_sc_hd__nor2_1 _15557_ (.A(_07786_),
    .B(_03547_),
    .Y(_00927_));
 sky130_fd_sc_hd__nor2_1 _15558_ (.A(_07800_),
    .B(_03547_),
    .Y(_00928_));
 sky130_fd_sc_hd__nor2_1 _15559_ (.A(_07809_),
    .B(_03547_),
    .Y(_00929_));
 sky130_fd_sc_hd__nor2_1 _15560_ (.A(_07818_),
    .B(_03547_),
    .Y(_00930_));
 sky130_fd_sc_hd__nor2_1 _15561_ (.A(_07831_),
    .B(_03547_),
    .Y(_00931_));
 sky130_fd_sc_hd__nor2_1 _15562_ (.A(_07843_),
    .B(_03547_),
    .Y(_00932_));
 sky130_fd_sc_hd__nor2_1 _15564_ (.A(_07850_),
    .B(_03547_),
    .Y(_00933_));
 sky130_fd_sc_hd__nor2_1 _15565_ (.A(_03491_),
    .B(_03547_),
    .Y(_00934_));
 sky130_fd_sc_hd__nor2_1 _15566_ (.A(_07581_),
    .B(_03547_),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_1 _15567_ (.A(_07873_),
    .B(_03547_),
    .Y(_00936_));
 sky130_fd_sc_hd__nor2_1 _15568_ (.A(_07925_),
    .B(_03547_),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2_1 _15569_ (.A(_07588_),
    .B(_03547_),
    .Y(_00938_));
 sky130_fd_sc_hd__nor2_1 _15570_ (.A(_07601_),
    .B(_03547_),
    .Y(_00939_));
 sky130_fd_sc_hd__nor2_1 _15571_ (.A(_07610_),
    .B(_03547_),
    .Y(_00940_));
 sky130_fd_sc_hd__nor2_1 _15572_ (.A(_07620_),
    .B(_03547_),
    .Y(_00941_));
 sky130_fd_sc_hd__nor2_1 _15573_ (.A(_07628_),
    .B(_03547_),
    .Y(_00942_));
 sky130_fd_sc_hd__nor2_1 _15574_ (.A(_07635_),
    .B(_03547_),
    .Y(_00943_));
 sky130_fd_sc_hd__nor2_1 _15575_ (.A(_07646_),
    .B(_03547_),
    .Y(_00944_));
 sky130_fd_sc_hd__nand2_1 _15576_ (.A(_05400_),
    .B(_08390_),
    .Y(_03551_));
 sky130_fd_sc_hd__nor2_1 _15578_ (.A(_07930_),
    .B(_03551_),
    .Y(_00945_));
 sky130_fd_sc_hd__nor2_1 _15579_ (.A(_08006_),
    .B(_03551_),
    .Y(_00946_));
 sky130_fd_sc_hd__nor2_1 _15580_ (.A(_08018_),
    .B(_03551_),
    .Y(_00947_));
 sky130_fd_sc_hd__nor2_1 _15581_ (.A(_08025_),
    .B(_03551_),
    .Y(_00948_));
 sky130_fd_sc_hd__nor2_1 _15582_ (.A(_08031_),
    .B(_03551_),
    .Y(_00949_));
 sky130_fd_sc_hd__nor2_1 _15583_ (.A(_08039_),
    .B(_03551_),
    .Y(_00950_));
 sky130_fd_sc_hd__nor2_1 _15584_ (.A(_08051_),
    .B(_03551_),
    .Y(_00951_));
 sky130_fd_sc_hd__nor2_1 _15585_ (.A(_08064_),
    .B(_03551_),
    .Y(_00952_));
 sky130_fd_sc_hd__nor2_1 _15586_ (.A(_08071_),
    .B(_03551_),
    .Y(_00953_));
 sky130_fd_sc_hd__nor2_1 _15587_ (.A(_08082_),
    .B(_03551_),
    .Y(_00954_));
 sky130_fd_sc_hd__nor2_1 _15589_ (.A(_08091_),
    .B(_03551_),
    .Y(_00955_));
 sky130_fd_sc_hd__nor2_1 _15590_ (.A(_07934_),
    .B(_03551_),
    .Y(_00956_));
 sky130_fd_sc_hd__nor2_1 _15591_ (.A(_08102_),
    .B(_03551_),
    .Y(_00957_));
 sky130_fd_sc_hd__nor2_1 _15592_ (.A(_08114_),
    .B(_03551_),
    .Y(_00958_));
 sky130_fd_sc_hd__nor2_1 _15593_ (.A(_08125_),
    .B(_03551_),
    .Y(_00959_));
 sky130_fd_sc_hd__nor2_1 _15594_ (.A(_08142_),
    .B(_03551_),
    .Y(_00960_));
 sky130_fd_sc_hd__nor2_1 _15595_ (.A(_08152_),
    .B(_03551_),
    .Y(_00961_));
 sky130_fd_sc_hd__nor2_1 _15596_ (.A(_08160_),
    .B(_03551_),
    .Y(_00962_));
 sky130_fd_sc_hd__nor2_1 _15597_ (.A(_08171_),
    .B(_03551_),
    .Y(_00963_));
 sky130_fd_sc_hd__nor2_1 _15598_ (.A(_08184_),
    .B(_03551_),
    .Y(_00964_));
 sky130_fd_sc_hd__nor2_1 _15600_ (.A(_08204_),
    .B(_03551_),
    .Y(_00965_));
 sky130_fd_sc_hd__nor2_1 _15601_ (.A(_08209_),
    .B(_03551_),
    .Y(_00966_));
 sky130_fd_sc_hd__nor2_1 _15602_ (.A(_07937_),
    .B(_03551_),
    .Y(_00967_));
 sky130_fd_sc_hd__nor2_1 _15603_ (.A(_08221_),
    .B(_03551_),
    .Y(_00968_));
 sky130_fd_sc_hd__nor2_1 _15604_ (.A(_08254_),
    .B(_03551_),
    .Y(_00969_));
 sky130_fd_sc_hd__nor2_1 _15605_ (.A(_07942_),
    .B(_03551_),
    .Y(_00970_));
 sky130_fd_sc_hd__nor2_1 _15606_ (.A(_07949_),
    .B(_03551_),
    .Y(_00971_));
 sky130_fd_sc_hd__nor2_1 _15607_ (.A(_07956_),
    .B(_03551_),
    .Y(_00972_));
 sky130_fd_sc_hd__nor2_1 _15608_ (.A(_07965_),
    .B(_03551_),
    .Y(_00973_));
 sky130_fd_sc_hd__nor2_1 _15609_ (.A(_07974_),
    .B(_03551_),
    .Y(_00974_));
 sky130_fd_sc_hd__nor2_1 _15610_ (.A(_07981_),
    .B(_03551_),
    .Y(_00975_));
 sky130_fd_sc_hd__nor2_1 _15611_ (.A(_07989_),
    .B(_03551_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_1 _15612_ (.A(_05350_),
    .B(_08431_),
    .Y(_03555_));
 sky130_fd_sc_hd__nor2_1 _15614_ (.A(_07572_),
    .B(_03555_),
    .Y(_00977_));
 sky130_fd_sc_hd__nor2_1 _15615_ (.A(_07660_),
    .B(_03555_),
    .Y(_00978_));
 sky130_fd_sc_hd__nor2_1 _15616_ (.A(_07669_),
    .B(_03555_),
    .Y(_00979_));
 sky130_fd_sc_hd__nor2_1 _15617_ (.A(_07677_),
    .B(_03555_),
    .Y(_00980_));
 sky130_fd_sc_hd__nor2_1 _15618_ (.A(_07689_),
    .B(_03555_),
    .Y(_00981_));
 sky130_fd_sc_hd__nor2_1 _15619_ (.A(_07703_),
    .B(_03555_),
    .Y(_00982_));
 sky130_fd_sc_hd__nor2_1 _15620_ (.A(_07709_),
    .B(_03555_),
    .Y(_00983_));
 sky130_fd_sc_hd__nor2_1 _15621_ (.A(_07715_),
    .B(_03555_),
    .Y(_00984_));
 sky130_fd_sc_hd__nor2_1 _15622_ (.A(_07731_),
    .B(_03555_),
    .Y(_00985_));
 sky130_fd_sc_hd__nor2_1 _15623_ (.A(_07745_),
    .B(_03555_),
    .Y(_00986_));
 sky130_fd_sc_hd__nor2_1 _15625_ (.A(_07752_),
    .B(_03555_),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _15626_ (.A(_07577_),
    .B(_03555_),
    .Y(_00988_));
 sky130_fd_sc_hd__nor2_1 _15627_ (.A(_07766_),
    .B(_03555_),
    .Y(_00989_));
 sky130_fd_sc_hd__nor2_1 _15628_ (.A(_07777_),
    .B(_03555_),
    .Y(_00990_));
 sky130_fd_sc_hd__nor2_1 _15629_ (.A(_07786_),
    .B(_03555_),
    .Y(_00991_));
 sky130_fd_sc_hd__nor2_1 _15630_ (.A(_07800_),
    .B(_03555_),
    .Y(_00992_));
 sky130_fd_sc_hd__nor2_1 _15631_ (.A(_07809_),
    .B(_03555_),
    .Y(_00993_));
 sky130_fd_sc_hd__nor2_1 _15632_ (.A(_07818_),
    .B(_03555_),
    .Y(_00994_));
 sky130_fd_sc_hd__nor2_1 _15633_ (.A(_07831_),
    .B(_03555_),
    .Y(_00995_));
 sky130_fd_sc_hd__nor2_1 _15634_ (.A(_07843_),
    .B(_03555_),
    .Y(_00996_));
 sky130_fd_sc_hd__nor2_1 _15636_ (.A(_07850_),
    .B(_03555_),
    .Y(_00997_));
 sky130_fd_sc_hd__nor2_1 _15637_ (.A(_03491_),
    .B(_03555_),
    .Y(_00998_));
 sky130_fd_sc_hd__nor2_1 _15638_ (.A(_07581_),
    .B(_03555_),
    .Y(_00999_));
 sky130_fd_sc_hd__nor2_1 _15639_ (.A(_07873_),
    .B(_03555_),
    .Y(_01000_));
 sky130_fd_sc_hd__nor2_1 _15640_ (.A(_07925_),
    .B(_03555_),
    .Y(_01001_));
 sky130_fd_sc_hd__nor2_1 _15641_ (.A(_07588_),
    .B(_03555_),
    .Y(_01002_));
 sky130_fd_sc_hd__nor2_1 _15642_ (.A(_07601_),
    .B(_03555_),
    .Y(_01003_));
 sky130_fd_sc_hd__nor2_1 _15643_ (.A(_07610_),
    .B(_03555_),
    .Y(_01004_));
 sky130_fd_sc_hd__nor2_1 _15644_ (.A(_07620_),
    .B(_03555_),
    .Y(_01005_));
 sky130_fd_sc_hd__nor2_1 _15645_ (.A(_07628_),
    .B(_03555_),
    .Y(_01006_));
 sky130_fd_sc_hd__nor2_1 _15646_ (.A(_07635_),
    .B(_03555_),
    .Y(_01007_));
 sky130_fd_sc_hd__nor2_1 _15647_ (.A(_07646_),
    .B(_03555_),
    .Y(_01008_));
 sky130_fd_sc_hd__or3_1 _15648_ (.A(reset),
    .B(_05399_),
    .C(_05409_),
    .X(_03559_));
 sky130_fd_sc_hd__nor2_1 _15651_ (.A(_07930_),
    .B(_03559_),
    .Y(_01009_));
 sky130_fd_sc_hd__nor2_1 _15652_ (.A(_08006_),
    .B(_03559_),
    .Y(_01010_));
 sky130_fd_sc_hd__nor2_1 _15653_ (.A(_08018_),
    .B(_03559_),
    .Y(_01011_));
 sky130_fd_sc_hd__nor2_1 _15654_ (.A(_08025_),
    .B(_03559_),
    .Y(_01012_));
 sky130_fd_sc_hd__nor2_1 _15655_ (.A(_08031_),
    .B(_03559_),
    .Y(_01013_));
 sky130_fd_sc_hd__nor2_1 _15656_ (.A(_08039_),
    .B(_03559_),
    .Y(_01014_));
 sky130_fd_sc_hd__nor2_1 _15657_ (.A(_08051_),
    .B(_03559_),
    .Y(_01015_));
 sky130_fd_sc_hd__nor2_1 _15658_ (.A(_08064_),
    .B(_03559_),
    .Y(_01016_));
 sky130_fd_sc_hd__nor2_1 _15659_ (.A(_08071_),
    .B(_03559_),
    .Y(_01017_));
 sky130_fd_sc_hd__nor2_1 _15660_ (.A(_08082_),
    .B(_03559_),
    .Y(_01018_));
 sky130_fd_sc_hd__nor2_1 _15662_ (.A(_08091_),
    .B(_03559_),
    .Y(_01019_));
 sky130_fd_sc_hd__nor2_1 _15663_ (.A(_07934_),
    .B(_03559_),
    .Y(_01020_));
 sky130_fd_sc_hd__nor2_1 _15664_ (.A(_08102_),
    .B(_03559_),
    .Y(_01021_));
 sky130_fd_sc_hd__nor2_1 _15665_ (.A(_08114_),
    .B(_03559_),
    .Y(_01022_));
 sky130_fd_sc_hd__nor2_1 _15666_ (.A(_08125_),
    .B(_03559_),
    .Y(_01023_));
 sky130_fd_sc_hd__nor2_1 _15667_ (.A(_08142_),
    .B(_03559_),
    .Y(_01024_));
 sky130_fd_sc_hd__nor2_1 _15668_ (.A(_08152_),
    .B(_03559_),
    .Y(_01025_));
 sky130_fd_sc_hd__nor2_1 _15669_ (.A(_08160_),
    .B(_03559_),
    .Y(_01026_));
 sky130_fd_sc_hd__nor2_1 _15670_ (.A(_08171_),
    .B(_03559_),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2_1 _15671_ (.A(_08184_),
    .B(_03559_),
    .Y(_01028_));
 sky130_fd_sc_hd__nor2_1 _15673_ (.A(_08204_),
    .B(_03559_),
    .Y(_01029_));
 sky130_fd_sc_hd__nor2_1 _15674_ (.A(_08209_),
    .B(_03559_),
    .Y(_01030_));
 sky130_fd_sc_hd__nor2_1 _15675_ (.A(_07937_),
    .B(_03559_),
    .Y(_01031_));
 sky130_fd_sc_hd__nor2_1 _15676_ (.A(_08221_),
    .B(_03559_),
    .Y(_01032_));
 sky130_fd_sc_hd__nor2_1 _15677_ (.A(_08254_),
    .B(_03559_),
    .Y(_01033_));
 sky130_fd_sc_hd__nor2_1 _15678_ (.A(_07942_),
    .B(_03559_),
    .Y(_01034_));
 sky130_fd_sc_hd__nor2_1 _15679_ (.A(_07949_),
    .B(_03559_),
    .Y(_01035_));
 sky130_fd_sc_hd__nor2_1 _15680_ (.A(_07956_),
    .B(_03559_),
    .Y(_01036_));
 sky130_fd_sc_hd__nor2_1 _15681_ (.A(_07965_),
    .B(_03559_),
    .Y(_01037_));
 sky130_fd_sc_hd__nor2_1 _15682_ (.A(_07974_),
    .B(_03559_),
    .Y(_01038_));
 sky130_fd_sc_hd__nor2_1 _15683_ (.A(_07981_),
    .B(_03559_),
    .Y(_01039_));
 sky130_fd_sc_hd__nor2_1 _15684_ (.A(_07989_),
    .B(_03559_),
    .Y(_01040_));
 sky130_fd_sc_hd__nand2_1 _15685_ (.A(_05356_),
    .B(_07566_),
    .Y(_03564_));
 sky130_fd_sc_hd__nor2_1 _15687_ (.A(_07572_),
    .B(_03564_),
    .Y(_01041_));
 sky130_fd_sc_hd__nor2_1 _15688_ (.A(_07660_),
    .B(_03564_),
    .Y(_01042_));
 sky130_fd_sc_hd__nor2_1 _15689_ (.A(_07669_),
    .B(_03564_),
    .Y(_01043_));
 sky130_fd_sc_hd__nor2_1 _15690_ (.A(_07677_),
    .B(_03564_),
    .Y(_01044_));
 sky130_fd_sc_hd__nor2_1 _15691_ (.A(_07689_),
    .B(_03564_),
    .Y(_01045_));
 sky130_fd_sc_hd__nor2_1 _15692_ (.A(_07703_),
    .B(_03564_),
    .Y(_01046_));
 sky130_fd_sc_hd__nor2_1 _15693_ (.A(_07709_),
    .B(_03564_),
    .Y(_01047_));
 sky130_fd_sc_hd__nor2_1 _15694_ (.A(_07715_),
    .B(_03564_),
    .Y(_01048_));
 sky130_fd_sc_hd__nor2_1 _15695_ (.A(_07731_),
    .B(_03564_),
    .Y(_01049_));
 sky130_fd_sc_hd__nor2_1 _15696_ (.A(_07745_),
    .B(_03564_),
    .Y(_01050_));
 sky130_fd_sc_hd__nor2_1 _15698_ (.A(_07752_),
    .B(_03564_),
    .Y(_01051_));
 sky130_fd_sc_hd__nor2_1 _15699_ (.A(_07577_),
    .B(_03564_),
    .Y(_01052_));
 sky130_fd_sc_hd__nor2_1 _15700_ (.A(_07766_),
    .B(_03564_),
    .Y(_01053_));
 sky130_fd_sc_hd__nor2_1 _15701_ (.A(_07777_),
    .B(_03564_),
    .Y(_01054_));
 sky130_fd_sc_hd__nor2_1 _15702_ (.A(_07786_),
    .B(_03564_),
    .Y(_01055_));
 sky130_fd_sc_hd__nor2_1 _15703_ (.A(_07800_),
    .B(_03564_),
    .Y(_01056_));
 sky130_fd_sc_hd__nor2_1 _15704_ (.A(_07809_),
    .B(_03564_),
    .Y(_01057_));
 sky130_fd_sc_hd__nor2_1 _15705_ (.A(_07818_),
    .B(_03564_),
    .Y(_01058_));
 sky130_fd_sc_hd__nor2_1 _15706_ (.A(_07831_),
    .B(_03564_),
    .Y(_01059_));
 sky130_fd_sc_hd__nor2_1 _15707_ (.A(_07843_),
    .B(_03564_),
    .Y(_01060_));
 sky130_fd_sc_hd__nor2_1 _15709_ (.A(_07850_),
    .B(_03564_),
    .Y(_01061_));
 sky130_fd_sc_hd__nor2_1 _15710_ (.A(_03491_),
    .B(_03564_),
    .Y(_01062_));
 sky130_fd_sc_hd__nor2_1 _15711_ (.A(_07581_),
    .B(_03564_),
    .Y(_01063_));
 sky130_fd_sc_hd__nor2_1 _15712_ (.A(_07873_),
    .B(_03564_),
    .Y(_01064_));
 sky130_fd_sc_hd__nor2_1 _15713_ (.A(_07925_),
    .B(_03564_),
    .Y(_01065_));
 sky130_fd_sc_hd__nor2_1 _15714_ (.A(_07588_),
    .B(_03564_),
    .Y(_01066_));
 sky130_fd_sc_hd__nor2_1 _15715_ (.A(_07601_),
    .B(_03564_),
    .Y(_01067_));
 sky130_fd_sc_hd__nor2_1 _15716_ (.A(_07610_),
    .B(_03564_),
    .Y(_01068_));
 sky130_fd_sc_hd__nor2_1 _15717_ (.A(_07620_),
    .B(_03564_),
    .Y(_01069_));
 sky130_fd_sc_hd__nor2_1 _15718_ (.A(_07628_),
    .B(_03564_),
    .Y(_01070_));
 sky130_fd_sc_hd__nor2_1 _15719_ (.A(_07635_),
    .B(_03564_),
    .Y(_01071_));
 sky130_fd_sc_hd__nor2_1 _15720_ (.A(_07646_),
    .B(_03564_),
    .Y(_01072_));
 sky130_fd_sc_hd__nand2_1 _15721_ (.A(_05411_),
    .B(_07927_),
    .Y(_03568_));
 sky130_fd_sc_hd__nor2_1 _15723_ (.A(_07930_),
    .B(_03568_),
    .Y(_01073_));
 sky130_fd_sc_hd__nor2_1 _15724_ (.A(_08006_),
    .B(_03568_),
    .Y(_01074_));
 sky130_fd_sc_hd__nor2_1 _15725_ (.A(_08018_),
    .B(_03568_),
    .Y(_01075_));
 sky130_fd_sc_hd__nor2_1 _15726_ (.A(_08025_),
    .B(_03568_),
    .Y(_01076_));
 sky130_fd_sc_hd__nor2_1 _15727_ (.A(_08031_),
    .B(_03568_),
    .Y(_01077_));
 sky130_fd_sc_hd__nor2_1 _15728_ (.A(_08039_),
    .B(_03568_),
    .Y(_01078_));
 sky130_fd_sc_hd__nor2_1 _15729_ (.A(_08051_),
    .B(_03568_),
    .Y(_01079_));
 sky130_fd_sc_hd__nor2_1 _15730_ (.A(_08064_),
    .B(_03568_),
    .Y(_01080_));
 sky130_fd_sc_hd__nor2_1 _15731_ (.A(_08071_),
    .B(_03568_),
    .Y(_01081_));
 sky130_fd_sc_hd__nor2_1 _15732_ (.A(_08082_),
    .B(_03568_),
    .Y(_01082_));
 sky130_fd_sc_hd__nor2_1 _15734_ (.A(_08091_),
    .B(_03568_),
    .Y(_01083_));
 sky130_fd_sc_hd__nor2_1 _15735_ (.A(_07934_),
    .B(_03568_),
    .Y(_01084_));
 sky130_fd_sc_hd__nor2_1 _15736_ (.A(_08102_),
    .B(_03568_),
    .Y(_01085_));
 sky130_fd_sc_hd__nor2_1 _15737_ (.A(_08114_),
    .B(_03568_),
    .Y(_01086_));
 sky130_fd_sc_hd__nor2_1 _15738_ (.A(_08125_),
    .B(_03568_),
    .Y(_01087_));
 sky130_fd_sc_hd__nor2_1 _15739_ (.A(_08142_),
    .B(_03568_),
    .Y(_01088_));
 sky130_fd_sc_hd__nor2_1 _15740_ (.A(_08152_),
    .B(_03568_),
    .Y(_01089_));
 sky130_fd_sc_hd__nor2_1 _15741_ (.A(_08160_),
    .B(_03568_),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _15742_ (.A(_08171_),
    .B(_03568_),
    .Y(_01091_));
 sky130_fd_sc_hd__nor2_1 _15743_ (.A(_08184_),
    .B(_03568_),
    .Y(_01092_));
 sky130_fd_sc_hd__nor2_1 _15745_ (.A(_08204_),
    .B(_03568_),
    .Y(_01093_));
 sky130_fd_sc_hd__nor2_1 _15746_ (.A(_08209_),
    .B(_03568_),
    .Y(_01094_));
 sky130_fd_sc_hd__nor2_1 _15747_ (.A(_07937_),
    .B(_03568_),
    .Y(_01095_));
 sky130_fd_sc_hd__nor2_1 _15748_ (.A(_08221_),
    .B(_03568_),
    .Y(_01096_));
 sky130_fd_sc_hd__nor2_1 _15749_ (.A(_08254_),
    .B(_03568_),
    .Y(_01097_));
 sky130_fd_sc_hd__nor2_1 _15750_ (.A(_07942_),
    .B(_03568_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_1 _15751_ (.A(_07949_),
    .B(_03568_),
    .Y(_01099_));
 sky130_fd_sc_hd__nor2_1 _15752_ (.A(_07956_),
    .B(_03568_),
    .Y(_01100_));
 sky130_fd_sc_hd__nor2_1 _15753_ (.A(_07965_),
    .B(_03568_),
    .Y(_01101_));
 sky130_fd_sc_hd__nor2_1 _15754_ (.A(_07974_),
    .B(_03568_),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_1 _15755_ (.A(_07981_),
    .B(_03568_),
    .Y(_01103_));
 sky130_fd_sc_hd__nor2_1 _15756_ (.A(_07989_),
    .B(_03568_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _15757_ (.A(_05356_),
    .B(_08257_),
    .Y(_03572_));
 sky130_fd_sc_hd__nor2_1 _15759_ (.A(_07572_),
    .B(_03572_),
    .Y(_01105_));
 sky130_fd_sc_hd__nor2_1 _15760_ (.A(_07660_),
    .B(_03572_),
    .Y(_01106_));
 sky130_fd_sc_hd__nor2_1 _15761_ (.A(_07669_),
    .B(_03572_),
    .Y(_01107_));
 sky130_fd_sc_hd__nor2_1 _15762_ (.A(_07677_),
    .B(_03572_),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _15763_ (.A(_07689_),
    .B(_03572_),
    .Y(_01109_));
 sky130_fd_sc_hd__nor2_1 _15764_ (.A(_07703_),
    .B(_03572_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(_07709_),
    .B(_03572_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_1 _15766_ (.A(_07715_),
    .B(_03572_),
    .Y(_01112_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_07731_),
    .B(_03572_),
    .Y(_01113_));
 sky130_fd_sc_hd__nor2_1 _15768_ (.A(_07745_),
    .B(_03572_),
    .Y(_01114_));
 sky130_fd_sc_hd__nor2_1 _15770_ (.A(_07752_),
    .B(_03572_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _15771_ (.A(_07577_),
    .B(_03572_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor2_1 _15772_ (.A(_07766_),
    .B(_03572_),
    .Y(_01117_));
 sky130_fd_sc_hd__nor2_1 _15773_ (.A(_07777_),
    .B(_03572_),
    .Y(_01118_));
 sky130_fd_sc_hd__nor2_1 _15774_ (.A(_07786_),
    .B(_03572_),
    .Y(_01119_));
 sky130_fd_sc_hd__nor2_1 _15775_ (.A(_07800_),
    .B(_03572_),
    .Y(_01120_));
 sky130_fd_sc_hd__nor2_1 _15776_ (.A(_07809_),
    .B(_03572_),
    .Y(_01121_));
 sky130_fd_sc_hd__nor2_1 _15777_ (.A(_07818_),
    .B(_03572_),
    .Y(_01122_));
 sky130_fd_sc_hd__nor2_1 _15778_ (.A(_07831_),
    .B(_03572_),
    .Y(_01123_));
 sky130_fd_sc_hd__nor2_1 _15779_ (.A(_07843_),
    .B(_03572_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _15781_ (.A(_07850_),
    .B(_03572_),
    .Y(_01125_));
 sky130_fd_sc_hd__nor2_1 _15782_ (.A(_03491_),
    .B(_03572_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_1 _15783_ (.A(_07581_),
    .B(_03572_),
    .Y(_01127_));
 sky130_fd_sc_hd__nor2_1 _15784_ (.A(_07873_),
    .B(_03572_),
    .Y(_01128_));
 sky130_fd_sc_hd__nor2_1 _15785_ (.A(_07925_),
    .B(_03572_),
    .Y(_01129_));
 sky130_fd_sc_hd__nor2_1 _15786_ (.A(_07588_),
    .B(_03572_),
    .Y(_01130_));
 sky130_fd_sc_hd__nor2_1 _15787_ (.A(_07601_),
    .B(_03572_),
    .Y(_01131_));
 sky130_fd_sc_hd__nor2_1 _15788_ (.A(_07610_),
    .B(_03572_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_1 _15789_ (.A(_07620_),
    .B(_03572_),
    .Y(_01133_));
 sky130_fd_sc_hd__nor2_1 _15790_ (.A(_07628_),
    .B(_03572_),
    .Y(_01134_));
 sky130_fd_sc_hd__nor2_1 _15791_ (.A(_07635_),
    .B(_03572_),
    .Y(_01135_));
 sky130_fd_sc_hd__nor2_1 _15792_ (.A(_07646_),
    .B(_03572_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand2_1 _15793_ (.A(_05411_),
    .B(_08304_),
    .Y(_03576_));
 sky130_fd_sc_hd__nor2_1 _15795_ (.A(_07930_),
    .B(_03576_),
    .Y(_01137_));
 sky130_fd_sc_hd__nor2_1 _15796_ (.A(_08006_),
    .B(_03576_),
    .Y(_01138_));
 sky130_fd_sc_hd__nor2_1 _15797_ (.A(_08018_),
    .B(_03576_),
    .Y(_01139_));
 sky130_fd_sc_hd__nor2_1 _15798_ (.A(_08025_),
    .B(_03576_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _15799_ (.A(_08031_),
    .B(_03576_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _15800_ (.A(_08039_),
    .B(_03576_),
    .Y(_01142_));
 sky130_fd_sc_hd__nor2_1 _15801_ (.A(_08051_),
    .B(_03576_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_1 _15802_ (.A(_08064_),
    .B(_03576_),
    .Y(_01144_));
 sky130_fd_sc_hd__nor2_1 _15803_ (.A(_08071_),
    .B(_03576_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _15804_ (.A(_08082_),
    .B(_03576_),
    .Y(_01146_));
 sky130_fd_sc_hd__nor2_1 _15806_ (.A(_08091_),
    .B(_03576_),
    .Y(_01147_));
 sky130_fd_sc_hd__nor2_1 _15807_ (.A(_07934_),
    .B(_03576_),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_1 _15808_ (.A(_08102_),
    .B(_03576_),
    .Y(_01149_));
 sky130_fd_sc_hd__nor2_1 _15809_ (.A(_08114_),
    .B(_03576_),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_1 _15810_ (.A(_08125_),
    .B(_03576_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _15811_ (.A(_08142_),
    .B(_03576_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor2_1 _15812_ (.A(_08152_),
    .B(_03576_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor2_1 _15813_ (.A(_08160_),
    .B(_03576_),
    .Y(_01154_));
 sky130_fd_sc_hd__nor2_1 _15814_ (.A(_08171_),
    .B(_03576_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _15815_ (.A(_08184_),
    .B(_03576_),
    .Y(_01156_));
 sky130_fd_sc_hd__nor2_1 _15817_ (.A(_08204_),
    .B(_03576_),
    .Y(_01157_));
 sky130_fd_sc_hd__nor2_1 _15818_ (.A(_08209_),
    .B(_03576_),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _15819_ (.A(_07937_),
    .B(_03576_),
    .Y(_01159_));
 sky130_fd_sc_hd__nor2_1 _15820_ (.A(_08221_),
    .B(_03576_),
    .Y(_01160_));
 sky130_fd_sc_hd__nor2_1 _15821_ (.A(_08254_),
    .B(_03576_),
    .Y(_01161_));
 sky130_fd_sc_hd__nor2_1 _15822_ (.A(_07942_),
    .B(_03576_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_1 _15823_ (.A(_07949_),
    .B(_03576_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_1 _15824_ (.A(_07956_),
    .B(_03576_),
    .Y(_01164_));
 sky130_fd_sc_hd__nor2_1 _15825_ (.A(_07965_),
    .B(_03576_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _15826_ (.A(_07974_),
    .B(_03576_),
    .Y(_01166_));
 sky130_fd_sc_hd__nor2_1 _15827_ (.A(_07981_),
    .B(_03576_),
    .Y(_01167_));
 sky130_fd_sc_hd__nor2_1 _15828_ (.A(_07989_),
    .B(_03576_),
    .Y(_01168_));
 sky130_fd_sc_hd__nand2_1 _15829_ (.A(_05356_),
    .B(_08346_),
    .Y(_03580_));
 sky130_fd_sc_hd__nor2_1 _15831_ (.A(_07572_),
    .B(_03580_),
    .Y(_01169_));
 sky130_fd_sc_hd__nor2_1 _15832_ (.A(_07660_),
    .B(_03580_),
    .Y(_01170_));
 sky130_fd_sc_hd__nor2_1 _15833_ (.A(_07669_),
    .B(_03580_),
    .Y(_01171_));
 sky130_fd_sc_hd__nor2_1 _15834_ (.A(_07677_),
    .B(_03580_),
    .Y(_01172_));
 sky130_fd_sc_hd__nor2_1 _15835_ (.A(_07689_),
    .B(_03580_),
    .Y(_01173_));
 sky130_fd_sc_hd__nor2_1 _15836_ (.A(_07703_),
    .B(_03580_),
    .Y(_01174_));
 sky130_fd_sc_hd__nor2_1 _15837_ (.A(_07709_),
    .B(_03580_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor2_1 _15838_ (.A(_07715_),
    .B(_03580_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2_1 _15839_ (.A(_07731_),
    .B(_03580_),
    .Y(_01177_));
 sky130_fd_sc_hd__nor2_1 _15840_ (.A(_07745_),
    .B(_03580_),
    .Y(_01178_));
 sky130_fd_sc_hd__nor2_1 _15842_ (.A(_07752_),
    .B(_03580_),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_1 _15843_ (.A(_07577_),
    .B(_03580_),
    .Y(_01180_));
 sky130_fd_sc_hd__nor2_1 _15844_ (.A(_07766_),
    .B(_03580_),
    .Y(_01181_));
 sky130_fd_sc_hd__nor2_1 _15845_ (.A(_07777_),
    .B(_03580_),
    .Y(_01182_));
 sky130_fd_sc_hd__nor2_1 _15846_ (.A(_07786_),
    .B(_03580_),
    .Y(_01183_));
 sky130_fd_sc_hd__nor2_1 _15847_ (.A(_07800_),
    .B(_03580_),
    .Y(_01184_));
 sky130_fd_sc_hd__nor2_1 _15848_ (.A(_07809_),
    .B(_03580_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_1 _15849_ (.A(_07818_),
    .B(_03580_),
    .Y(_01186_));
 sky130_fd_sc_hd__nor2_1 _15850_ (.A(_07831_),
    .B(_03580_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_1 _15851_ (.A(_07843_),
    .B(_03580_),
    .Y(_01188_));
 sky130_fd_sc_hd__nor2_1 _15853_ (.A(_07850_),
    .B(_03580_),
    .Y(_01189_));
 sky130_fd_sc_hd__nor2_1 _15854_ (.A(_03491_),
    .B(_03580_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _15855_ (.A(_07581_),
    .B(_03580_),
    .Y(_01191_));
 sky130_fd_sc_hd__nor2_1 _15856_ (.A(_07873_),
    .B(_03580_),
    .Y(_01192_));
 sky130_fd_sc_hd__nor2_1 _15857_ (.A(_07925_),
    .B(_03580_),
    .Y(_01193_));
 sky130_fd_sc_hd__nor2_1 _15858_ (.A(_07588_),
    .B(_03580_),
    .Y(_01194_));
 sky130_fd_sc_hd__nor2_1 _15859_ (.A(_07601_),
    .B(_03580_),
    .Y(_01195_));
 sky130_fd_sc_hd__nor2_1 _15860_ (.A(_07610_),
    .B(_03580_),
    .Y(_01196_));
 sky130_fd_sc_hd__nor2_1 _15861_ (.A(_07620_),
    .B(_03580_),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_1 _15862_ (.A(_07628_),
    .B(_03580_),
    .Y(_01198_));
 sky130_fd_sc_hd__nor2_1 _15863_ (.A(_07635_),
    .B(_03580_),
    .Y(_01199_));
 sky130_fd_sc_hd__nor2_1 _15864_ (.A(_07646_),
    .B(_03580_),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _15865_ (.A(_05411_),
    .B(_08390_),
    .Y(_03584_));
 sky130_fd_sc_hd__nor2_1 _15867_ (.A(_07930_),
    .B(_03584_),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _15868_ (.A(_08006_),
    .B(_03584_),
    .Y(_01202_));
 sky130_fd_sc_hd__nor2_1 _15869_ (.A(_08018_),
    .B(_03584_),
    .Y(_01203_));
 sky130_fd_sc_hd__nor2_1 _15870_ (.A(_08025_),
    .B(_03584_),
    .Y(_01204_));
 sky130_fd_sc_hd__nor2_1 _15871_ (.A(_08031_),
    .B(_03584_),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_1 _15872_ (.A(_08039_),
    .B(_03584_),
    .Y(_01206_));
 sky130_fd_sc_hd__nor2_1 _15873_ (.A(_08051_),
    .B(_03584_),
    .Y(_01207_));
 sky130_fd_sc_hd__nor2_1 _15874_ (.A(_08064_),
    .B(_03584_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _15875_ (.A(_08071_),
    .B(_03584_),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_1 _15876_ (.A(_08082_),
    .B(_03584_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor2_1 _15878_ (.A(_08091_),
    .B(_03584_),
    .Y(_01211_));
 sky130_fd_sc_hd__nor2_1 _15879_ (.A(_07934_),
    .B(_03584_),
    .Y(_01212_));
 sky130_fd_sc_hd__nor2_1 _15880_ (.A(_08102_),
    .B(_03584_),
    .Y(_01213_));
 sky130_fd_sc_hd__nor2_1 _15881_ (.A(_08114_),
    .B(_03584_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_1 _15882_ (.A(_08125_),
    .B(_03584_),
    .Y(_01215_));
 sky130_fd_sc_hd__nor2_1 _15883_ (.A(_08142_),
    .B(_03584_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_1 _15884_ (.A(_08152_),
    .B(_03584_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _15885_ (.A(_08160_),
    .B(_03584_),
    .Y(_01218_));
 sky130_fd_sc_hd__nor2_1 _15886_ (.A(_08171_),
    .B(_03584_),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_1 _15887_ (.A(_08184_),
    .B(_03584_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor2_1 _15889_ (.A(_08204_),
    .B(_03584_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _15890_ (.A(_08209_),
    .B(_03584_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_1 _15891_ (.A(_07937_),
    .B(_03584_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_1 _15892_ (.A(_08221_),
    .B(_03584_),
    .Y(_01224_));
 sky130_fd_sc_hd__nor2_1 _15893_ (.A(_08254_),
    .B(_03584_),
    .Y(_01225_));
 sky130_fd_sc_hd__nor2_1 _15894_ (.A(_07942_),
    .B(_03584_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _15895_ (.A(_07949_),
    .B(_03584_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor2_1 _15896_ (.A(_07956_),
    .B(_03584_),
    .Y(_01228_));
 sky130_fd_sc_hd__nor2_1 _15897_ (.A(_07965_),
    .B(_03584_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_1 _15898_ (.A(_07974_),
    .B(_03584_),
    .Y(_01230_));
 sky130_fd_sc_hd__nor2_1 _15899_ (.A(_07981_),
    .B(_03584_),
    .Y(_01231_));
 sky130_fd_sc_hd__nor2_1 _15900_ (.A(_07989_),
    .B(_03584_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_1 _15901_ (.A(_05356_),
    .B(_08431_),
    .Y(_03588_));
 sky130_fd_sc_hd__nor2_1 _15903_ (.A(_07572_),
    .B(_03588_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_1 _15904_ (.A(_07660_),
    .B(_03588_),
    .Y(_01234_));
 sky130_fd_sc_hd__nor2_1 _15905_ (.A(_07669_),
    .B(_03588_),
    .Y(_01235_));
 sky130_fd_sc_hd__nor2_1 _15906_ (.A(_07677_),
    .B(_03588_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_1 _15907_ (.A(_07689_),
    .B(_03588_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _15908_ (.A(_07703_),
    .B(_03588_),
    .Y(_01238_));
 sky130_fd_sc_hd__nor2_1 _15909_ (.A(_07709_),
    .B(_03588_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _15910_ (.A(_07715_),
    .B(_03588_),
    .Y(_01240_));
 sky130_fd_sc_hd__nor2_1 _15911_ (.A(_07731_),
    .B(_03588_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_1 _15912_ (.A(_07745_),
    .B(_03588_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_1 _15914_ (.A(_07752_),
    .B(_03588_),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _15915_ (.A(_07577_),
    .B(_03588_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _15916_ (.A(_07766_),
    .B(_03588_),
    .Y(_01245_));
 sky130_fd_sc_hd__nor2_1 _15917_ (.A(_07777_),
    .B(_03588_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _15918_ (.A(_07786_),
    .B(_03588_),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_1 _15919_ (.A(_07800_),
    .B(_03588_),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _15920_ (.A(_07809_),
    .B(_03588_),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_1 _15921_ (.A(_07818_),
    .B(_03588_),
    .Y(_01250_));
 sky130_fd_sc_hd__nor2_1 _15922_ (.A(_07831_),
    .B(_03588_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor2_1 _15923_ (.A(_07843_),
    .B(_03588_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _15925_ (.A(_07850_),
    .B(_03588_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor2_1 _15926_ (.A(_03491_),
    .B(_03588_),
    .Y(_01254_));
 sky130_fd_sc_hd__nor2_1 _15927_ (.A(_07581_),
    .B(_03588_),
    .Y(_01255_));
 sky130_fd_sc_hd__nor2_1 _15928_ (.A(_07873_),
    .B(_03588_),
    .Y(_01256_));
 sky130_fd_sc_hd__nor2_1 _15929_ (.A(_07925_),
    .B(_03588_),
    .Y(_01257_));
 sky130_fd_sc_hd__nor2_1 _15930_ (.A(_07588_),
    .B(_03588_),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _15931_ (.A(_07601_),
    .B(_03588_),
    .Y(_01259_));
 sky130_fd_sc_hd__nor2_1 _15932_ (.A(_07610_),
    .B(_03588_),
    .Y(_01260_));
 sky130_fd_sc_hd__nor2_1 _15933_ (.A(_07620_),
    .B(_03588_),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_1 _15934_ (.A(_07628_),
    .B(_03588_),
    .Y(_01262_));
 sky130_fd_sc_hd__nor2_1 _15935_ (.A(_07635_),
    .B(_03588_),
    .Y(_01263_));
 sky130_fd_sc_hd__nor2_1 _15936_ (.A(_07646_),
    .B(_03588_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand2_1 _15937_ (.A(_05411_),
    .B(_08803_),
    .Y(_03592_));
 sky130_fd_sc_hd__nor2_1 _15939_ (.A(_07930_),
    .B(_03592_),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _15940_ (.A(_08006_),
    .B(_03592_),
    .Y(_01266_));
 sky130_fd_sc_hd__nor2_1 _15941_ (.A(_08018_),
    .B(_03592_),
    .Y(_01267_));
 sky130_fd_sc_hd__nor2_1 _15942_ (.A(_08025_),
    .B(_03592_),
    .Y(_01268_));
 sky130_fd_sc_hd__nor2_1 _15943_ (.A(_08031_),
    .B(_03592_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_1 _15944_ (.A(_08039_),
    .B(_03592_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _15945_ (.A(_08051_),
    .B(_03592_),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_1 _15946_ (.A(_08064_),
    .B(_03592_),
    .Y(_01272_));
 sky130_fd_sc_hd__nor2_1 _15947_ (.A(_08071_),
    .B(_03592_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor2_1 _15948_ (.A(_08082_),
    .B(_03592_),
    .Y(_01274_));
 sky130_fd_sc_hd__nor2_1 _15950_ (.A(_08091_),
    .B(_03592_),
    .Y(_01275_));
 sky130_fd_sc_hd__nor2_1 _15951_ (.A(_07934_),
    .B(_03592_),
    .Y(_01276_));
 sky130_fd_sc_hd__nor2_1 _15952_ (.A(_08102_),
    .B(_03592_),
    .Y(_01277_));
 sky130_fd_sc_hd__nor2_1 _15953_ (.A(_08114_),
    .B(_03592_),
    .Y(_01278_));
 sky130_fd_sc_hd__nor2_1 _15954_ (.A(_08125_),
    .B(_03592_),
    .Y(_01279_));
 sky130_fd_sc_hd__nor2_1 _15955_ (.A(_08142_),
    .B(_03592_),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_1 _15956_ (.A(_08152_),
    .B(_03592_),
    .Y(_01281_));
 sky130_fd_sc_hd__nor2_1 _15957_ (.A(_08160_),
    .B(_03592_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor2_1 _15958_ (.A(_08171_),
    .B(_03592_),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_1 _15959_ (.A(_08184_),
    .B(_03592_),
    .Y(_01284_));
 sky130_fd_sc_hd__nor2_1 _15961_ (.A(_08204_),
    .B(_03592_),
    .Y(_01285_));
 sky130_fd_sc_hd__nor2_1 _15962_ (.A(_08209_),
    .B(_03592_),
    .Y(_01286_));
 sky130_fd_sc_hd__nor2_1 _15963_ (.A(_07937_),
    .B(_03592_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_1 _15964_ (.A(_08221_),
    .B(_03592_),
    .Y(_01288_));
 sky130_fd_sc_hd__nor2_1 _15965_ (.A(_08254_),
    .B(_03592_),
    .Y(_01289_));
 sky130_fd_sc_hd__nor2_1 _15966_ (.A(_07942_),
    .B(_03592_),
    .Y(_01290_));
 sky130_fd_sc_hd__nor2_1 _15967_ (.A(_07949_),
    .B(_03592_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_1 _15968_ (.A(_07956_),
    .B(_03592_),
    .Y(_01292_));
 sky130_fd_sc_hd__nor2_1 _15969_ (.A(_07965_),
    .B(_03592_),
    .Y(_01293_));
 sky130_fd_sc_hd__nor2_1 _15970_ (.A(_07974_),
    .B(_03592_),
    .Y(_01294_));
 sky130_fd_sc_hd__nor2_1 _15971_ (.A(_07981_),
    .B(_03592_),
    .Y(_01295_));
 sky130_fd_sc_hd__nor2_1 _15972_ (.A(_07989_),
    .B(_03592_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand2_1 _15973_ (.A(_05364_),
    .B(_07566_),
    .Y(_03596_));
 sky130_fd_sc_hd__nor2_1 _15975_ (.A(_07572_),
    .B(_03596_),
    .Y(_01297_));
 sky130_fd_sc_hd__nor2_1 _15976_ (.A(_07660_),
    .B(_03596_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_1 _15977_ (.A(_07669_),
    .B(_03596_),
    .Y(_01299_));
 sky130_fd_sc_hd__nor2_1 _15978_ (.A(_07677_),
    .B(_03596_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _15979_ (.A(_07689_),
    .B(_03596_),
    .Y(_01301_));
 sky130_fd_sc_hd__nor2_1 _15980_ (.A(_07703_),
    .B(_03596_),
    .Y(_01302_));
 sky130_fd_sc_hd__nor2_1 _15981_ (.A(_07709_),
    .B(_03596_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_1 _15982_ (.A(_07715_),
    .B(_03596_),
    .Y(_01304_));
 sky130_fd_sc_hd__nor2_1 _15983_ (.A(_07731_),
    .B(_03596_),
    .Y(_01305_));
 sky130_fd_sc_hd__nor2_1 _15984_ (.A(_07745_),
    .B(_03596_),
    .Y(_01306_));
 sky130_fd_sc_hd__nor2_1 _15986_ (.A(_07752_),
    .B(_03596_),
    .Y(_01307_));
 sky130_fd_sc_hd__nor2_1 _15987_ (.A(_07577_),
    .B(_03596_),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_1 _15988_ (.A(_07766_),
    .B(_03596_),
    .Y(_01309_));
 sky130_fd_sc_hd__nor2_1 _15989_ (.A(_07777_),
    .B(_03596_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor2_1 _15990_ (.A(_07786_),
    .B(_03596_),
    .Y(_01311_));
 sky130_fd_sc_hd__nor2_1 _15991_ (.A(_07800_),
    .B(_03596_),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _15992_ (.A(_07809_),
    .B(_03596_),
    .Y(_01313_));
 sky130_fd_sc_hd__nor2_1 _15993_ (.A(_07818_),
    .B(_03596_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_1 _15994_ (.A(_07831_),
    .B(_03596_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2_1 _15995_ (.A(_07843_),
    .B(_03596_),
    .Y(_01316_));
 sky130_fd_sc_hd__nor2_1 _15997_ (.A(_07850_),
    .B(_03596_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_1 _15998_ (.A(_03491_),
    .B(_03596_),
    .Y(_01318_));
 sky130_fd_sc_hd__nor2_1 _15999_ (.A(_07581_),
    .B(_03596_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_1 _16000_ (.A(_07873_),
    .B(_03596_),
    .Y(_01320_));
 sky130_fd_sc_hd__nor2_1 _16001_ (.A(_07925_),
    .B(_03596_),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2_1 _16002_ (.A(_07588_),
    .B(_03596_),
    .Y(_01322_));
 sky130_fd_sc_hd__nor2_1 _16003_ (.A(_07601_),
    .B(_03596_),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2_1 _16004_ (.A(_07610_),
    .B(_03596_),
    .Y(_01324_));
 sky130_fd_sc_hd__nor2_1 _16005_ (.A(_07620_),
    .B(_03596_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_1 _16006_ (.A(_07628_),
    .B(_03596_),
    .Y(_01326_));
 sky130_fd_sc_hd__nor2_1 _16007_ (.A(_07635_),
    .B(_03596_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_1 _16008_ (.A(_07646_),
    .B(_03596_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _16009_ (.A(_05417_),
    .B(_07927_),
    .Y(_03600_));
 sky130_fd_sc_hd__nor2_1 _16011_ (.A(_07930_),
    .B(_03600_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _16012_ (.A(_08006_),
    .B(_03600_),
    .Y(_01330_));
 sky130_fd_sc_hd__nor2_1 _16013_ (.A(_08018_),
    .B(_03600_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2_1 _16014_ (.A(_08025_),
    .B(_03600_),
    .Y(_01332_));
 sky130_fd_sc_hd__nor2_1 _16015_ (.A(_08031_),
    .B(_03600_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2_1 _16016_ (.A(_08039_),
    .B(_03600_),
    .Y(_01334_));
 sky130_fd_sc_hd__nor2_1 _16017_ (.A(_08051_),
    .B(_03600_),
    .Y(_01335_));
 sky130_fd_sc_hd__nor2_1 _16018_ (.A(_08064_),
    .B(_03600_),
    .Y(_01336_));
 sky130_fd_sc_hd__nor2_1 _16019_ (.A(_08071_),
    .B(_03600_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2_1 _16020_ (.A(_08082_),
    .B(_03600_),
    .Y(_01338_));
 sky130_fd_sc_hd__nor2_1 _16022_ (.A(_08091_),
    .B(_03600_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2_1 _16023_ (.A(_07934_),
    .B(_03600_),
    .Y(_01340_));
 sky130_fd_sc_hd__nor2_1 _16024_ (.A(_08102_),
    .B(_03600_),
    .Y(_01341_));
 sky130_fd_sc_hd__nor2_1 _16025_ (.A(_08114_),
    .B(_03600_),
    .Y(_01342_));
 sky130_fd_sc_hd__nor2_1 _16026_ (.A(_08125_),
    .B(_03600_),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_1 _16027_ (.A(_08142_),
    .B(_03600_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _16028_ (.A(_08152_),
    .B(_03600_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _16029_ (.A(_08160_),
    .B(_03600_),
    .Y(_01346_));
 sky130_fd_sc_hd__nor2_1 _16030_ (.A(_08171_),
    .B(_03600_),
    .Y(_01347_));
 sky130_fd_sc_hd__nor2_1 _16031_ (.A(_08184_),
    .B(_03600_),
    .Y(_01348_));
 sky130_fd_sc_hd__nor2_1 _16033_ (.A(_08204_),
    .B(_03600_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2_1 _16034_ (.A(_08209_),
    .B(_03600_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor2_1 _16035_ (.A(_07937_),
    .B(_03600_),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2_1 _16036_ (.A(_08221_),
    .B(_03600_),
    .Y(_01352_));
 sky130_fd_sc_hd__nor2_1 _16037_ (.A(_08254_),
    .B(_03600_),
    .Y(_01353_));
 sky130_fd_sc_hd__nor2_1 _16038_ (.A(_07942_),
    .B(_03600_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor2_1 _16039_ (.A(_07949_),
    .B(_03600_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2_1 _16040_ (.A(_07956_),
    .B(_03600_),
    .Y(_01356_));
 sky130_fd_sc_hd__nor2_1 _16041_ (.A(_07965_),
    .B(_03600_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_1 _16042_ (.A(_07974_),
    .B(_03600_),
    .Y(_01358_));
 sky130_fd_sc_hd__nor2_1 _16043_ (.A(_07981_),
    .B(_03600_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _16044_ (.A(_07989_),
    .B(_03600_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(_05364_),
    .B(_08257_),
    .Y(_03604_));
 sky130_fd_sc_hd__nor2_1 _16047_ (.A(_07572_),
    .B(_03604_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2_1 _16048_ (.A(_07660_),
    .B(_03604_),
    .Y(_01362_));
 sky130_fd_sc_hd__nor2_1 _16049_ (.A(_07669_),
    .B(_03604_),
    .Y(_01363_));
 sky130_fd_sc_hd__nor2_1 _16050_ (.A(_07677_),
    .B(_03604_),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_1 _16051_ (.A(_07689_),
    .B(_03604_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_1 _16052_ (.A(_07703_),
    .B(_03604_),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_1 _16053_ (.A(_07709_),
    .B(_03604_),
    .Y(_01367_));
 sky130_fd_sc_hd__nor2_1 _16054_ (.A(_07715_),
    .B(_03604_),
    .Y(_01368_));
 sky130_fd_sc_hd__nor2_1 _16055_ (.A(_07731_),
    .B(_03604_),
    .Y(_01369_));
 sky130_fd_sc_hd__nor2_1 _16056_ (.A(_07745_),
    .B(_03604_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _16058_ (.A(_07752_),
    .B(_03604_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_1 _16059_ (.A(_07577_),
    .B(_03604_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_1 _16060_ (.A(_07766_),
    .B(_03604_),
    .Y(_01373_));
 sky130_fd_sc_hd__nor2_1 _16061_ (.A(_07777_),
    .B(_03604_),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_1 _16062_ (.A(_07786_),
    .B(_03604_),
    .Y(_01375_));
 sky130_fd_sc_hd__nor2_1 _16063_ (.A(_07800_),
    .B(_03604_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _16064_ (.A(_07809_),
    .B(_03604_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _16065_ (.A(_07818_),
    .B(_03604_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_1 _16066_ (.A(_07831_),
    .B(_03604_),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_1 _16067_ (.A(_07843_),
    .B(_03604_),
    .Y(_01380_));
 sky130_fd_sc_hd__nor2_1 _16069_ (.A(_07850_),
    .B(_03604_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _16070_ (.A(_03491_),
    .B(_03604_),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_1 _16071_ (.A(_07581_),
    .B(_03604_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _16072_ (.A(_07873_),
    .B(_03604_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_1 _16073_ (.A(_07925_),
    .B(_03604_),
    .Y(_01385_));
 sky130_fd_sc_hd__nor2_1 _16074_ (.A(_07588_),
    .B(_03604_),
    .Y(_01386_));
 sky130_fd_sc_hd__nor2_1 _16075_ (.A(_07601_),
    .B(_03604_),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_1 _16076_ (.A(_07610_),
    .B(_03604_),
    .Y(_01388_));
 sky130_fd_sc_hd__nor2_1 _16077_ (.A(_07620_),
    .B(_03604_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _16078_ (.A(_07628_),
    .B(_03604_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_1 _16079_ (.A(_07635_),
    .B(_03604_),
    .Y(_01391_));
 sky130_fd_sc_hd__nor2_1 _16080_ (.A(_07646_),
    .B(_03604_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(_05417_),
    .B(_08304_),
    .Y(_03608_));
 sky130_fd_sc_hd__nor2_1 _16083_ (.A(_07930_),
    .B(_03608_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _16084_ (.A(_08006_),
    .B(_03608_),
    .Y(_01394_));
 sky130_fd_sc_hd__nor2_1 _16085_ (.A(_08018_),
    .B(_03608_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2_1 _16086_ (.A(_08025_),
    .B(_03608_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _16087_ (.A(_08031_),
    .B(_03608_),
    .Y(_01397_));
 sky130_fd_sc_hd__nor2_1 _16088_ (.A(_08039_),
    .B(_03608_),
    .Y(_01398_));
 sky130_fd_sc_hd__nor2_1 _16089_ (.A(_08051_),
    .B(_03608_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor2_1 _16090_ (.A(_08064_),
    .B(_03608_),
    .Y(_01400_));
 sky130_fd_sc_hd__nor2_1 _16091_ (.A(_08071_),
    .B(_03608_),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_1 _16092_ (.A(_08082_),
    .B(_03608_),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_1 _16094_ (.A(_08091_),
    .B(_03608_),
    .Y(_01403_));
 sky130_fd_sc_hd__nor2_1 _16095_ (.A(_07934_),
    .B(_03608_),
    .Y(_01404_));
 sky130_fd_sc_hd__nor2_1 _16096_ (.A(_08102_),
    .B(_03608_),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _16097_ (.A(_08114_),
    .B(_03608_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _16098_ (.A(_08125_),
    .B(_03608_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _16099_ (.A(_08142_),
    .B(_03608_),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_1 _16100_ (.A(_08152_),
    .B(_03608_),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_1 _16101_ (.A(_08160_),
    .B(_03608_),
    .Y(_01410_));
 sky130_fd_sc_hd__nor2_1 _16102_ (.A(_08171_),
    .B(_03608_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor2_1 _16103_ (.A(_08184_),
    .B(_03608_),
    .Y(_01412_));
 sky130_fd_sc_hd__nor2_1 _16105_ (.A(_08204_),
    .B(_03608_),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_1 _16106_ (.A(_08209_),
    .B(_03608_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _16107_ (.A(_07937_),
    .B(_03608_),
    .Y(_01415_));
 sky130_fd_sc_hd__nor2_1 _16108_ (.A(_08221_),
    .B(_03608_),
    .Y(_01416_));
 sky130_fd_sc_hd__nor2_1 _16109_ (.A(_08254_),
    .B(_03608_),
    .Y(_01417_));
 sky130_fd_sc_hd__nor2_1 _16110_ (.A(_07942_),
    .B(_03608_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _16111_ (.A(_07949_),
    .B(_03608_),
    .Y(_01419_));
 sky130_fd_sc_hd__nor2_1 _16112_ (.A(_07956_),
    .B(_03608_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_1 _16113_ (.A(_07965_),
    .B(_03608_),
    .Y(_01421_));
 sky130_fd_sc_hd__nor2_1 _16114_ (.A(_07974_),
    .B(_03608_),
    .Y(_01422_));
 sky130_fd_sc_hd__nor2_1 _16115_ (.A(_07981_),
    .B(_03608_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _16116_ (.A(_07989_),
    .B(_03608_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand2_1 _16118_ (.A(_05364_),
    .B(_08346_),
    .Y(_03613_));
 sky130_fd_sc_hd__nor2_1 _16120_ (.A(_07572_),
    .B(_03613_),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_1 _16122_ (.A(_07660_),
    .B(_03613_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_1 _16124_ (.A(_07669_),
    .B(_03613_),
    .Y(_01427_));
 sky130_fd_sc_hd__nor2_1 _16126_ (.A(_07677_),
    .B(_03613_),
    .Y(_01428_));
 sky130_fd_sc_hd__nor2_1 _16128_ (.A(_07689_),
    .B(_03613_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _16130_ (.A(_07703_),
    .B(_03613_),
    .Y(_01430_));
 sky130_fd_sc_hd__nor2_1 _16132_ (.A(_07709_),
    .B(_03613_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_1 _16134_ (.A(_07715_),
    .B(_03613_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_1 _16136_ (.A(_07731_),
    .B(_03613_),
    .Y(_01433_));
 sky130_fd_sc_hd__nor2_1 _16138_ (.A(_07745_),
    .B(_03613_),
    .Y(_01434_));
 sky130_fd_sc_hd__nor2_1 _16141_ (.A(_07752_),
    .B(_03613_),
    .Y(_01435_));
 sky130_fd_sc_hd__nor2_1 _16143_ (.A(_07577_),
    .B(_03613_),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_1 _16145_ (.A(_07766_),
    .B(_03613_),
    .Y(_01437_));
 sky130_fd_sc_hd__nor2_1 _16147_ (.A(_07777_),
    .B(_03613_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _16149_ (.A(_07786_),
    .B(_03613_),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_1 _16151_ (.A(_07800_),
    .B(_03613_),
    .Y(_01440_));
 sky130_fd_sc_hd__nor2_1 _16153_ (.A(_07809_),
    .B(_03613_),
    .Y(_01441_));
 sky130_fd_sc_hd__nor2_1 _16155_ (.A(_07818_),
    .B(_03613_),
    .Y(_01442_));
 sky130_fd_sc_hd__nor2_1 _16157_ (.A(_07831_),
    .B(_03613_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2_1 _16159_ (.A(_07843_),
    .B(_03613_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _16162_ (.A(_07850_),
    .B(_03613_),
    .Y(_01445_));
 sky130_fd_sc_hd__nor2_1 _16164_ (.A(_03491_),
    .B(_03613_),
    .Y(_01446_));
 sky130_fd_sc_hd__nor2_1 _16166_ (.A(_07581_),
    .B(_03613_),
    .Y(_01447_));
 sky130_fd_sc_hd__nor2_1 _16168_ (.A(_07873_),
    .B(_03613_),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_1 _16170_ (.A(_07925_),
    .B(_03613_),
    .Y(_01449_));
 sky130_fd_sc_hd__nor2_1 _16172_ (.A(_07588_),
    .B(_03613_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _16174_ (.A(_07601_),
    .B(_03613_),
    .Y(_01451_));
 sky130_fd_sc_hd__nor2_1 _16176_ (.A(_07610_),
    .B(_03613_),
    .Y(_01452_));
 sky130_fd_sc_hd__nor2_1 _16178_ (.A(_07620_),
    .B(_03613_),
    .Y(_01453_));
 sky130_fd_sc_hd__nor2_1 _16180_ (.A(_07628_),
    .B(_03613_),
    .Y(_01454_));
 sky130_fd_sc_hd__nor2_1 _16182_ (.A(_07635_),
    .B(_03613_),
    .Y(_01455_));
 sky130_fd_sc_hd__nor2_1 _16184_ (.A(_07646_),
    .B(_03613_),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_1 _16186_ (.A(_05417_),
    .B(_08390_),
    .Y(_03649_));
 sky130_fd_sc_hd__nor2_1 _16188_ (.A(_07930_),
    .B(_03649_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor2_1 _16190_ (.A(_08006_),
    .B(_03649_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_1 _16192_ (.A(_08018_),
    .B(_03649_),
    .Y(_01459_));
 sky130_fd_sc_hd__nor2_1 _16194_ (.A(_08025_),
    .B(_03649_),
    .Y(_01460_));
 sky130_fd_sc_hd__nor2_1 _16196_ (.A(_08031_),
    .B(_03649_),
    .Y(_01461_));
 sky130_fd_sc_hd__nor2_1 _16198_ (.A(_08039_),
    .B(_03649_),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_1 _16200_ (.A(_08051_),
    .B(_03649_),
    .Y(_01463_));
 sky130_fd_sc_hd__nor2_1 _16202_ (.A(_08064_),
    .B(_03649_),
    .Y(_01464_));
 sky130_fd_sc_hd__nor2_1 _16204_ (.A(_08071_),
    .B(_03649_),
    .Y(_01465_));
 sky130_fd_sc_hd__nor2_1 _16206_ (.A(_08082_),
    .B(_03649_),
    .Y(_01466_));
 sky130_fd_sc_hd__nor2_1 _16209_ (.A(_08091_),
    .B(_03649_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _16211_ (.A(_07934_),
    .B(_03649_),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_1 _16213_ (.A(_08102_),
    .B(_03649_),
    .Y(_01469_));
 sky130_fd_sc_hd__nor2_1 _16215_ (.A(_08114_),
    .B(_03649_),
    .Y(_01470_));
 sky130_fd_sc_hd__nor2_1 _16217_ (.A(_08125_),
    .B(_03649_),
    .Y(_01471_));
 sky130_fd_sc_hd__nor2_1 _16219_ (.A(_08142_),
    .B(_03649_),
    .Y(_01472_));
 sky130_fd_sc_hd__nor2_1 _16221_ (.A(_08152_),
    .B(_03649_),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_1 _16223_ (.A(_08160_),
    .B(_03649_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor2_1 _16225_ (.A(_08171_),
    .B(_03649_),
    .Y(_01475_));
 sky130_fd_sc_hd__nor2_1 _16227_ (.A(_08184_),
    .B(_03649_),
    .Y(_01476_));
 sky130_fd_sc_hd__nor2_1 _16230_ (.A(_08204_),
    .B(_03649_),
    .Y(_01477_));
 sky130_fd_sc_hd__nor2_1 _16232_ (.A(_08209_),
    .B(_03649_),
    .Y(_01478_));
 sky130_fd_sc_hd__nor2_1 _16234_ (.A(_07937_),
    .B(_03649_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_1 _16236_ (.A(_08221_),
    .B(_03649_),
    .Y(_01480_));
 sky130_fd_sc_hd__nor2_1 _16238_ (.A(_08254_),
    .B(_03649_),
    .Y(_01481_));
 sky130_fd_sc_hd__nor2_1 _16240_ (.A(_07942_),
    .B(_03649_),
    .Y(_01482_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(_07949_),
    .B(_03649_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _16244_ (.A(_07956_),
    .B(_03649_),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_1 _16246_ (.A(_07965_),
    .B(_03649_),
    .Y(_01485_));
 sky130_fd_sc_hd__nor2_1 _16248_ (.A(_07974_),
    .B(_03649_),
    .Y(_01486_));
 sky130_fd_sc_hd__nor2_1 _16250_ (.A(_07981_),
    .B(_03649_),
    .Y(_01487_));
 sky130_fd_sc_hd__nor2_1 _16252_ (.A(_07989_),
    .B(_03649_),
    .Y(_01488_));
 sky130_fd_sc_hd__nand2_1 _16253_ (.A(_05364_),
    .B(_08431_),
    .Y(_03684_));
 sky130_fd_sc_hd__nor2_1 _16255_ (.A(_07572_),
    .B(_03684_),
    .Y(_01489_));
 sky130_fd_sc_hd__nor2_1 _16256_ (.A(_07660_),
    .B(_03684_),
    .Y(_01490_));
 sky130_fd_sc_hd__nor2_1 _16257_ (.A(_07669_),
    .B(_03684_),
    .Y(_01491_));
 sky130_fd_sc_hd__nor2_1 _16258_ (.A(_07677_),
    .B(_03684_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_1 _16259_ (.A(_07689_),
    .B(_03684_),
    .Y(_01493_));
 sky130_fd_sc_hd__nor2_1 _16260_ (.A(_07703_),
    .B(_03684_),
    .Y(_01494_));
 sky130_fd_sc_hd__nor2_1 _16261_ (.A(_07709_),
    .B(_03684_),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_1 _16262_ (.A(_07715_),
    .B(_03684_),
    .Y(_01496_));
 sky130_fd_sc_hd__nor2_1 _16263_ (.A(_07731_),
    .B(_03684_),
    .Y(_01497_));
 sky130_fd_sc_hd__nor2_1 _16264_ (.A(_07745_),
    .B(_03684_),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_1 _16266_ (.A(_07752_),
    .B(_03684_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _16267_ (.A(_07577_),
    .B(_03684_),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_1 _16268_ (.A(_07766_),
    .B(_03684_),
    .Y(_01501_));
 sky130_fd_sc_hd__nor2_1 _16269_ (.A(_07777_),
    .B(_03684_),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _16270_ (.A(_07786_),
    .B(_03684_),
    .Y(_01503_));
 sky130_fd_sc_hd__nor2_1 _16271_ (.A(_07800_),
    .B(_03684_),
    .Y(_01504_));
 sky130_fd_sc_hd__nor2_1 _16272_ (.A(_07809_),
    .B(_03684_),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_1 _16273_ (.A(_07818_),
    .B(_03684_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_1 _16274_ (.A(_07831_),
    .B(_03684_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_1 _16275_ (.A(_07843_),
    .B(_03684_),
    .Y(_01508_));
 sky130_fd_sc_hd__nor2_1 _16277_ (.A(_07850_),
    .B(_03684_),
    .Y(_01509_));
 sky130_fd_sc_hd__nor2_1 _16278_ (.A(_03491_),
    .B(_03684_),
    .Y(_01510_));
 sky130_fd_sc_hd__nor2_1 _16279_ (.A(_07581_),
    .B(_03684_),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_1 _16280_ (.A(_07873_),
    .B(_03684_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_1 _16281_ (.A(_07925_),
    .B(_03684_),
    .Y(_01513_));
 sky130_fd_sc_hd__nor2_1 _16282_ (.A(_07588_),
    .B(_03684_),
    .Y(_01514_));
 sky130_fd_sc_hd__nor2_1 _16283_ (.A(_07601_),
    .B(_03684_),
    .Y(_01515_));
 sky130_fd_sc_hd__nor2_1 _16284_ (.A(_07610_),
    .B(_03684_),
    .Y(_01516_));
 sky130_fd_sc_hd__nor2_1 _16285_ (.A(_07620_),
    .B(_03684_),
    .Y(_01517_));
 sky130_fd_sc_hd__nor2_1 _16286_ (.A(_07628_),
    .B(_03684_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor2_1 _16287_ (.A(_07635_),
    .B(_03684_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor2_1 _16288_ (.A(_07646_),
    .B(_03684_),
    .Y(_01520_));
 sky130_fd_sc_hd__nand3_1 _16289_ (.A(_09567_),
    .B(\count_2[5] ),
    .C(_08476_),
    .Y(_03688_));
 sky130_fd_sc_hd__nor2_1 _16291_ (.A(_07930_),
    .B(_03688_),
    .Y(_01521_));
 sky130_fd_sc_hd__nor2_1 _16292_ (.A(_08006_),
    .B(_03688_),
    .Y(_01522_));
 sky130_fd_sc_hd__nor2_1 _16293_ (.A(_08018_),
    .B(_03688_),
    .Y(_01523_));
 sky130_fd_sc_hd__nor2_1 _16294_ (.A(_08025_),
    .B(_03688_),
    .Y(_01524_));
 sky130_fd_sc_hd__nor2_1 _16295_ (.A(_08031_),
    .B(_03688_),
    .Y(_01525_));
 sky130_fd_sc_hd__nor2_1 _16296_ (.A(_08039_),
    .B(_03688_),
    .Y(_01526_));
 sky130_fd_sc_hd__nor2_1 _16297_ (.A(_08051_),
    .B(_03688_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _16298_ (.A(_08064_),
    .B(_03688_),
    .Y(_01528_));
 sky130_fd_sc_hd__nor2_1 _16299_ (.A(_08071_),
    .B(_03688_),
    .Y(_01529_));
 sky130_fd_sc_hd__nor2_1 _16300_ (.A(_08082_),
    .B(_03688_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _16302_ (.A(_08091_),
    .B(_03688_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _16303_ (.A(_07934_),
    .B(_03688_),
    .Y(_01532_));
 sky130_fd_sc_hd__nor2_1 _16304_ (.A(_08102_),
    .B(_03688_),
    .Y(_01533_));
 sky130_fd_sc_hd__nor2_1 _16305_ (.A(_08114_),
    .B(_03688_),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _16306_ (.A(_08125_),
    .B(_03688_),
    .Y(_01535_));
 sky130_fd_sc_hd__nor2_1 _16307_ (.A(_08142_),
    .B(_03688_),
    .Y(_01536_));
 sky130_fd_sc_hd__nor2_1 _16308_ (.A(_08152_),
    .B(_03688_),
    .Y(_01537_));
 sky130_fd_sc_hd__nor2_1 _16309_ (.A(_08160_),
    .B(_03688_),
    .Y(_01538_));
 sky130_fd_sc_hd__nor2_1 _16310_ (.A(_08171_),
    .B(_03688_),
    .Y(_01539_));
 sky130_fd_sc_hd__nor2_1 _16311_ (.A(_08184_),
    .B(_03688_),
    .Y(_01540_));
 sky130_fd_sc_hd__nor2_1 _16313_ (.A(_08204_),
    .B(_03688_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _16314_ (.A(_08209_),
    .B(_03688_),
    .Y(_01542_));
 sky130_fd_sc_hd__nor2_1 _16315_ (.A(_07937_),
    .B(_03688_),
    .Y(_01543_));
 sky130_fd_sc_hd__nor2_1 _16316_ (.A(_08221_),
    .B(_03688_),
    .Y(_01544_));
 sky130_fd_sc_hd__nor2_1 _16317_ (.A(_08254_),
    .B(_03688_),
    .Y(_01545_));
 sky130_fd_sc_hd__nor2_1 _16318_ (.A(_07942_),
    .B(_03688_),
    .Y(_01546_));
 sky130_fd_sc_hd__nor2_1 _16319_ (.A(_07949_),
    .B(_03688_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_1 _16320_ (.A(_07956_),
    .B(_03688_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _16321_ (.A(_07965_),
    .B(_03688_),
    .Y(_01549_));
 sky130_fd_sc_hd__nor2_1 _16322_ (.A(_07974_),
    .B(_03688_),
    .Y(_01550_));
 sky130_fd_sc_hd__nor2_1 _16323_ (.A(_07981_),
    .B(_03688_),
    .Y(_01551_));
 sky130_fd_sc_hd__nor2_1 _16324_ (.A(_07989_),
    .B(_03688_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand2_1 _16325_ (.A(_05369_),
    .B(_07566_),
    .Y(_03692_));
 sky130_fd_sc_hd__nor2_1 _16327_ (.A(_07572_),
    .B(_03692_),
    .Y(_01553_));
 sky130_fd_sc_hd__nor2_1 _16328_ (.A(_07660_),
    .B(_03692_),
    .Y(_01554_));
 sky130_fd_sc_hd__nor2_1 _16329_ (.A(_07669_),
    .B(_03692_),
    .Y(_01555_));
 sky130_fd_sc_hd__nor2_1 _16330_ (.A(_07677_),
    .B(_03692_),
    .Y(_01556_));
 sky130_fd_sc_hd__nor2_1 _16331_ (.A(_07689_),
    .B(_03692_),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2_1 _16332_ (.A(_07703_),
    .B(_03692_),
    .Y(_01558_));
 sky130_fd_sc_hd__nor2_1 _16333_ (.A(_07709_),
    .B(_03692_),
    .Y(_01559_));
 sky130_fd_sc_hd__nor2_1 _16334_ (.A(_07715_),
    .B(_03692_),
    .Y(_01560_));
 sky130_fd_sc_hd__nor2_1 _16335_ (.A(_07731_),
    .B(_03692_),
    .Y(_01561_));
 sky130_fd_sc_hd__nor2_1 _16336_ (.A(_07745_),
    .B(_03692_),
    .Y(_01562_));
 sky130_fd_sc_hd__nor2_1 _16338_ (.A(_07752_),
    .B(_03692_),
    .Y(_01563_));
 sky130_fd_sc_hd__nor2_1 _16339_ (.A(_07577_),
    .B(_03692_),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_1 _16340_ (.A(_07766_),
    .B(_03692_),
    .Y(_01565_));
 sky130_fd_sc_hd__nor2_1 _16341_ (.A(_07777_),
    .B(_03692_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_1 _16342_ (.A(_07786_),
    .B(_03692_),
    .Y(_01567_));
 sky130_fd_sc_hd__nor2_1 _16343_ (.A(_07800_),
    .B(_03692_),
    .Y(_01568_));
 sky130_fd_sc_hd__nor2_1 _16344_ (.A(_07809_),
    .B(_03692_),
    .Y(_01569_));
 sky130_fd_sc_hd__nor2_1 _16345_ (.A(_07818_),
    .B(_03692_),
    .Y(_01570_));
 sky130_fd_sc_hd__nor2_1 _16346_ (.A(_07831_),
    .B(_03692_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_1 _16347_ (.A(_07843_),
    .B(_03692_),
    .Y(_01572_));
 sky130_fd_sc_hd__nor2_1 _16349_ (.A(_07850_),
    .B(_03692_),
    .Y(_01573_));
 sky130_fd_sc_hd__nor2_1 _16350_ (.A(_03491_),
    .B(_03692_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor2_1 _16351_ (.A(_07581_),
    .B(_03692_),
    .Y(_01575_));
 sky130_fd_sc_hd__nor2_1 _16352_ (.A(_07873_),
    .B(_03692_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _16353_ (.A(_07925_),
    .B(_03692_),
    .Y(_01577_));
 sky130_fd_sc_hd__nor2_1 _16354_ (.A(_07588_),
    .B(_03692_),
    .Y(_01578_));
 sky130_fd_sc_hd__nor2_1 _16355_ (.A(_07601_),
    .B(_03692_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _16356_ (.A(_07610_),
    .B(_03692_),
    .Y(_01580_));
 sky130_fd_sc_hd__nor2_1 _16357_ (.A(_07620_),
    .B(_03692_),
    .Y(_01581_));
 sky130_fd_sc_hd__nor2_1 _16358_ (.A(_07628_),
    .B(_03692_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_1 _16359_ (.A(_07635_),
    .B(_03692_),
    .Y(_01583_));
 sky130_fd_sc_hd__nor2_1 _16360_ (.A(_07646_),
    .B(_03692_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _16361_ (.A(_05424_),
    .B(_07927_),
    .Y(_03696_));
 sky130_fd_sc_hd__nor2_1 _16363_ (.A(_07930_),
    .B(_03696_),
    .Y(_01585_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_08006_),
    .B(_03696_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor2_1 _16365_ (.A(_08018_),
    .B(_03696_),
    .Y(_01587_));
 sky130_fd_sc_hd__nor2_1 _16366_ (.A(_08025_),
    .B(_03696_),
    .Y(_01588_));
 sky130_fd_sc_hd__nor2_1 _16367_ (.A(_08031_),
    .B(_03696_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_1 _16368_ (.A(_08039_),
    .B(_03696_),
    .Y(_01590_));
 sky130_fd_sc_hd__nor2_1 _16369_ (.A(_08051_),
    .B(_03696_),
    .Y(_01591_));
 sky130_fd_sc_hd__nor2_1 _16370_ (.A(_08064_),
    .B(_03696_),
    .Y(_01592_));
 sky130_fd_sc_hd__nor2_1 _16371_ (.A(_08071_),
    .B(_03696_),
    .Y(_01593_));
 sky130_fd_sc_hd__nor2_1 _16372_ (.A(_08082_),
    .B(_03696_),
    .Y(_01594_));
 sky130_fd_sc_hd__nor2_1 _16374_ (.A(_08091_),
    .B(_03696_),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_1 _16375_ (.A(_07934_),
    .B(_03696_),
    .Y(_01596_));
 sky130_fd_sc_hd__nor2_1 _16376_ (.A(_08102_),
    .B(_03696_),
    .Y(_01597_));
 sky130_fd_sc_hd__nor2_1 _16377_ (.A(_08114_),
    .B(_03696_),
    .Y(_01598_));
 sky130_fd_sc_hd__nor2_1 _16378_ (.A(_08125_),
    .B(_03696_),
    .Y(_01599_));
 sky130_fd_sc_hd__nor2_1 _16379_ (.A(_08142_),
    .B(_03696_),
    .Y(_01600_));
 sky130_fd_sc_hd__nor2_1 _16380_ (.A(_08152_),
    .B(_03696_),
    .Y(_01601_));
 sky130_fd_sc_hd__nor2_1 _16381_ (.A(_08160_),
    .B(_03696_),
    .Y(_01602_));
 sky130_fd_sc_hd__nor2_1 _16382_ (.A(_08171_),
    .B(_03696_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _16383_ (.A(_08184_),
    .B(_03696_),
    .Y(_01604_));
 sky130_fd_sc_hd__nor2_1 _16385_ (.A(_08204_),
    .B(_03696_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _16386_ (.A(_08209_),
    .B(_03696_),
    .Y(_01606_));
 sky130_fd_sc_hd__nor2_1 _16387_ (.A(_07937_),
    .B(_03696_),
    .Y(_01607_));
 sky130_fd_sc_hd__nor2_1 _16388_ (.A(_08221_),
    .B(_03696_),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_1 _16389_ (.A(_08254_),
    .B(_03696_),
    .Y(_01609_));
 sky130_fd_sc_hd__nor2_1 _16390_ (.A(_07942_),
    .B(_03696_),
    .Y(_01610_));
 sky130_fd_sc_hd__nor2_1 _16391_ (.A(_07949_),
    .B(_03696_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_1 _16392_ (.A(_07956_),
    .B(_03696_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_1 _16393_ (.A(_07965_),
    .B(_03696_),
    .Y(_01613_));
 sky130_fd_sc_hd__nor2_1 _16394_ (.A(_07974_),
    .B(_03696_),
    .Y(_01614_));
 sky130_fd_sc_hd__nor2_1 _16395_ (.A(_07981_),
    .B(_03696_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_1 _16396_ (.A(_07989_),
    .B(_03696_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _16397_ (.A(_05369_),
    .B(_08257_),
    .Y(_03700_));
 sky130_fd_sc_hd__nor2_1 _16399_ (.A(_07572_),
    .B(_03700_),
    .Y(_01617_));
 sky130_fd_sc_hd__nor2_1 _16400_ (.A(_07660_),
    .B(_03700_),
    .Y(_01618_));
 sky130_fd_sc_hd__nor2_1 _16401_ (.A(_07669_),
    .B(_03700_),
    .Y(_01619_));
 sky130_fd_sc_hd__nor2_1 _16402_ (.A(_07677_),
    .B(_03700_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _16403_ (.A(_07689_),
    .B(_03700_),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_1 _16404_ (.A(_07703_),
    .B(_03700_),
    .Y(_01622_));
 sky130_fd_sc_hd__nor2_1 _16405_ (.A(_07709_),
    .B(_03700_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_1 _16406_ (.A(_07715_),
    .B(_03700_),
    .Y(_01624_));
 sky130_fd_sc_hd__nor2_1 _16407_ (.A(_07731_),
    .B(_03700_),
    .Y(_01625_));
 sky130_fd_sc_hd__nor2_1 _16408_ (.A(_07745_),
    .B(_03700_),
    .Y(_01626_));
 sky130_fd_sc_hd__nor2_1 _16410_ (.A(_07752_),
    .B(_03700_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _16411_ (.A(_07577_),
    .B(_03700_),
    .Y(_01628_));
 sky130_fd_sc_hd__nor2_1 _16412_ (.A(_07766_),
    .B(_03700_),
    .Y(_01629_));
 sky130_fd_sc_hd__nor2_1 _16413_ (.A(_07777_),
    .B(_03700_),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_1 _16414_ (.A(_07786_),
    .B(_03700_),
    .Y(_01631_));
 sky130_fd_sc_hd__nor2_1 _16415_ (.A(_07800_),
    .B(_03700_),
    .Y(_01632_));
 sky130_fd_sc_hd__nor2_1 _16416_ (.A(_07809_),
    .B(_03700_),
    .Y(_01633_));
 sky130_fd_sc_hd__nor2_1 _16417_ (.A(_07818_),
    .B(_03700_),
    .Y(_01634_));
 sky130_fd_sc_hd__nor2_1 _16418_ (.A(_07831_),
    .B(_03700_),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_1 _16419_ (.A(_07843_),
    .B(_03700_),
    .Y(_01636_));
 sky130_fd_sc_hd__nor2_1 _16421_ (.A(_07850_),
    .B(_03700_),
    .Y(_01637_));
 sky130_fd_sc_hd__nor2_1 _16422_ (.A(_03491_),
    .B(_03700_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor2_1 _16423_ (.A(_07581_),
    .B(_03700_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_1 _16424_ (.A(_07873_),
    .B(_03700_),
    .Y(_01640_));
 sky130_fd_sc_hd__nor2_1 _16425_ (.A(_07925_),
    .B(_03700_),
    .Y(_01641_));
 sky130_fd_sc_hd__nor2_1 _16426_ (.A(_07588_),
    .B(_03700_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor2_1 _16427_ (.A(_07601_),
    .B(_03700_),
    .Y(_01643_));
 sky130_fd_sc_hd__nor2_1 _16428_ (.A(_07610_),
    .B(_03700_),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _16429_ (.A(_07620_),
    .B(_03700_),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_1 _16430_ (.A(_07628_),
    .B(_03700_),
    .Y(_01646_));
 sky130_fd_sc_hd__nor2_1 _16431_ (.A(_07635_),
    .B(_03700_),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_1 _16432_ (.A(_07646_),
    .B(_03700_),
    .Y(_01648_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(_05424_),
    .B(_08304_),
    .Y(_03704_));
 sky130_fd_sc_hd__nor2_1 _16435_ (.A(_07930_),
    .B(_03704_),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_1 _16436_ (.A(_08006_),
    .B(_03704_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _16437_ (.A(_08018_),
    .B(_03704_),
    .Y(_01651_));
 sky130_fd_sc_hd__nor2_1 _16438_ (.A(_08025_),
    .B(_03704_),
    .Y(_01652_));
 sky130_fd_sc_hd__nor2_1 _16439_ (.A(_08031_),
    .B(_03704_),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _16440_ (.A(_08039_),
    .B(_03704_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_1 _16441_ (.A(_08051_),
    .B(_03704_),
    .Y(_01655_));
 sky130_fd_sc_hd__nor2_1 _16442_ (.A(_08064_),
    .B(_03704_),
    .Y(_01656_));
 sky130_fd_sc_hd__nor2_1 _16443_ (.A(_08071_),
    .B(_03704_),
    .Y(_01657_));
 sky130_fd_sc_hd__nor2_1 _16444_ (.A(_08082_),
    .B(_03704_),
    .Y(_01658_));
 sky130_fd_sc_hd__nor2_1 _16446_ (.A(_08091_),
    .B(_03704_),
    .Y(_01659_));
 sky130_fd_sc_hd__nor2_1 _16447_ (.A(_07934_),
    .B(_03704_),
    .Y(_01660_));
 sky130_fd_sc_hd__nor2_1 _16448_ (.A(_08102_),
    .B(_03704_),
    .Y(_01661_));
 sky130_fd_sc_hd__nor2_1 _16449_ (.A(_08114_),
    .B(_03704_),
    .Y(_01662_));
 sky130_fd_sc_hd__nor2_1 _16450_ (.A(_08125_),
    .B(_03704_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor2_1 _16451_ (.A(_08142_),
    .B(_03704_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_1 _16452_ (.A(_08152_),
    .B(_03704_),
    .Y(_01665_));
 sky130_fd_sc_hd__nor2_1 _16453_ (.A(_08160_),
    .B(_03704_),
    .Y(_01666_));
 sky130_fd_sc_hd__nor2_1 _16454_ (.A(_08171_),
    .B(_03704_),
    .Y(_01667_));
 sky130_fd_sc_hd__nor2_1 _16455_ (.A(_08184_),
    .B(_03704_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _16457_ (.A(_08204_),
    .B(_03704_),
    .Y(_01669_));
 sky130_fd_sc_hd__nor2_1 _16458_ (.A(_08209_),
    .B(_03704_),
    .Y(_01670_));
 sky130_fd_sc_hd__nor2_1 _16459_ (.A(_07937_),
    .B(_03704_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_1 _16460_ (.A(_08221_),
    .B(_03704_),
    .Y(_01672_));
 sky130_fd_sc_hd__nor2_1 _16461_ (.A(_08254_),
    .B(_03704_),
    .Y(_01673_));
 sky130_fd_sc_hd__nor2_1 _16462_ (.A(_07942_),
    .B(_03704_),
    .Y(_01674_));
 sky130_fd_sc_hd__nor2_1 _16463_ (.A(_07949_),
    .B(_03704_),
    .Y(_01675_));
 sky130_fd_sc_hd__nor2_1 _16464_ (.A(_07956_),
    .B(_03704_),
    .Y(_01676_));
 sky130_fd_sc_hd__nor2_1 _16465_ (.A(_07965_),
    .B(_03704_),
    .Y(_01677_));
 sky130_fd_sc_hd__nor2_1 _16466_ (.A(_07974_),
    .B(_03704_),
    .Y(_01678_));
 sky130_fd_sc_hd__nor2_1 _16467_ (.A(_07981_),
    .B(_03704_),
    .Y(_01679_));
 sky130_fd_sc_hd__nor2_1 _16468_ (.A(_07989_),
    .B(_03704_),
    .Y(_01680_));
 sky130_fd_sc_hd__nand2_1 _16469_ (.A(_05369_),
    .B(_08346_),
    .Y(_03708_));
 sky130_fd_sc_hd__nor2_1 _16471_ (.A(_07572_),
    .B(_03708_),
    .Y(_01681_));
 sky130_fd_sc_hd__nor2_1 _16472_ (.A(_07660_),
    .B(_03708_),
    .Y(_01682_));
 sky130_fd_sc_hd__nor2_1 _16473_ (.A(_07669_),
    .B(_03708_),
    .Y(_01683_));
 sky130_fd_sc_hd__nor2_1 _16474_ (.A(_07677_),
    .B(_03708_),
    .Y(_01684_));
 sky130_fd_sc_hd__nor2_1 _16475_ (.A(_07689_),
    .B(_03708_),
    .Y(_01685_));
 sky130_fd_sc_hd__nor2_1 _16476_ (.A(_07703_),
    .B(_03708_),
    .Y(_01686_));
 sky130_fd_sc_hd__nor2_1 _16477_ (.A(_07709_),
    .B(_03708_),
    .Y(_01687_));
 sky130_fd_sc_hd__nor2_1 _16478_ (.A(_07715_),
    .B(_03708_),
    .Y(_01688_));
 sky130_fd_sc_hd__nor2_1 _16479_ (.A(_07731_),
    .B(_03708_),
    .Y(_01689_));
 sky130_fd_sc_hd__nor2_1 _16480_ (.A(_07745_),
    .B(_03708_),
    .Y(_01690_));
 sky130_fd_sc_hd__nor2_1 _16482_ (.A(_07752_),
    .B(_03708_),
    .Y(_01691_));
 sky130_fd_sc_hd__nor2_1 _16483_ (.A(_07577_),
    .B(_03708_),
    .Y(_01692_));
 sky130_fd_sc_hd__nor2_1 _16484_ (.A(_07766_),
    .B(_03708_),
    .Y(_01693_));
 sky130_fd_sc_hd__nor2_1 _16485_ (.A(_07777_),
    .B(_03708_),
    .Y(_01694_));
 sky130_fd_sc_hd__nor2_1 _16486_ (.A(_07786_),
    .B(_03708_),
    .Y(_01695_));
 sky130_fd_sc_hd__nor2_1 _16487_ (.A(_07800_),
    .B(_03708_),
    .Y(_01696_));
 sky130_fd_sc_hd__nor2_1 _16488_ (.A(_07809_),
    .B(_03708_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_1 _16489_ (.A(_07818_),
    .B(_03708_),
    .Y(_01698_));
 sky130_fd_sc_hd__nor2_1 _16490_ (.A(_07831_),
    .B(_03708_),
    .Y(_01699_));
 sky130_fd_sc_hd__nor2_1 _16491_ (.A(_07843_),
    .B(_03708_),
    .Y(_01700_));
 sky130_fd_sc_hd__nor2_1 _16493_ (.A(_07850_),
    .B(_03708_),
    .Y(_01701_));
 sky130_fd_sc_hd__nor2_1 _16494_ (.A(_03491_),
    .B(_03708_),
    .Y(_01702_));
 sky130_fd_sc_hd__nor2_1 _16495_ (.A(_07581_),
    .B(_03708_),
    .Y(_01703_));
 sky130_fd_sc_hd__nor2_1 _16496_ (.A(_07873_),
    .B(_03708_),
    .Y(_01704_));
 sky130_fd_sc_hd__nor2_1 _16497_ (.A(_07925_),
    .B(_03708_),
    .Y(_01705_));
 sky130_fd_sc_hd__nor2_1 _16498_ (.A(_07588_),
    .B(_03708_),
    .Y(_01706_));
 sky130_fd_sc_hd__nor2_1 _16499_ (.A(_07601_),
    .B(_03708_),
    .Y(_01707_));
 sky130_fd_sc_hd__nor2_1 _16500_ (.A(_07610_),
    .B(_03708_),
    .Y(_01708_));
 sky130_fd_sc_hd__nor2_1 _16501_ (.A(_07620_),
    .B(_03708_),
    .Y(_01709_));
 sky130_fd_sc_hd__nor2_1 _16502_ (.A(_07628_),
    .B(_03708_),
    .Y(_01710_));
 sky130_fd_sc_hd__nor2_1 _16503_ (.A(_07635_),
    .B(_03708_),
    .Y(_01711_));
 sky130_fd_sc_hd__nor2_1 _16504_ (.A(_07646_),
    .B(_03708_),
    .Y(_01712_));
 sky130_fd_sc_hd__nand2_1 _16505_ (.A(_05424_),
    .B(_08390_),
    .Y(_03712_));
 sky130_fd_sc_hd__nor2_1 _16507_ (.A(_07930_),
    .B(_03712_),
    .Y(_01713_));
 sky130_fd_sc_hd__nor2_1 _16508_ (.A(_08006_),
    .B(_03712_),
    .Y(_01714_));
 sky130_fd_sc_hd__nor2_1 _16509_ (.A(_08018_),
    .B(_03712_),
    .Y(_01715_));
 sky130_fd_sc_hd__nor2_1 _16510_ (.A(_08025_),
    .B(_03712_),
    .Y(_01716_));
 sky130_fd_sc_hd__nor2_1 _16511_ (.A(_08031_),
    .B(_03712_),
    .Y(_01717_));
 sky130_fd_sc_hd__nor2_1 _16512_ (.A(_08039_),
    .B(_03712_),
    .Y(_01718_));
 sky130_fd_sc_hd__nor2_1 _16513_ (.A(_08051_),
    .B(_03712_),
    .Y(_01719_));
 sky130_fd_sc_hd__nor2_1 _16514_ (.A(_08064_),
    .B(_03712_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor2_1 _16515_ (.A(_08071_),
    .B(_03712_),
    .Y(_01721_));
 sky130_fd_sc_hd__nor2_1 _16516_ (.A(_08082_),
    .B(_03712_),
    .Y(_01722_));
 sky130_fd_sc_hd__nor2_1 _16518_ (.A(_08091_),
    .B(_03712_),
    .Y(_01723_));
 sky130_fd_sc_hd__nor2_1 _16519_ (.A(_07934_),
    .B(_03712_),
    .Y(_01724_));
 sky130_fd_sc_hd__nor2_1 _16520_ (.A(_08102_),
    .B(_03712_),
    .Y(_01725_));
 sky130_fd_sc_hd__nor2_1 _16521_ (.A(_08114_),
    .B(_03712_),
    .Y(_01726_));
 sky130_fd_sc_hd__nor2_1 _16522_ (.A(_08125_),
    .B(_03712_),
    .Y(_01727_));
 sky130_fd_sc_hd__nor2_1 _16523_ (.A(_08142_),
    .B(_03712_),
    .Y(_01728_));
 sky130_fd_sc_hd__nor2_1 _16524_ (.A(_08152_),
    .B(_03712_),
    .Y(_01729_));
 sky130_fd_sc_hd__nor2_1 _16525_ (.A(_08160_),
    .B(_03712_),
    .Y(_01730_));
 sky130_fd_sc_hd__nor2_1 _16526_ (.A(_08171_),
    .B(_03712_),
    .Y(_01731_));
 sky130_fd_sc_hd__nor2_1 _16527_ (.A(_08184_),
    .B(_03712_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_1 _16529_ (.A(_08204_),
    .B(_03712_),
    .Y(_01733_));
 sky130_fd_sc_hd__nor2_1 _16530_ (.A(_08209_),
    .B(_03712_),
    .Y(_01734_));
 sky130_fd_sc_hd__nor2_1 _16531_ (.A(_07937_),
    .B(_03712_),
    .Y(_01735_));
 sky130_fd_sc_hd__nor2_1 _16532_ (.A(_08221_),
    .B(_03712_),
    .Y(_01736_));
 sky130_fd_sc_hd__nor2_1 _16533_ (.A(_08254_),
    .B(_03712_),
    .Y(_01737_));
 sky130_fd_sc_hd__nor2_1 _16534_ (.A(_07942_),
    .B(_03712_),
    .Y(_01738_));
 sky130_fd_sc_hd__nor2_1 _16535_ (.A(_07949_),
    .B(_03712_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _16536_ (.A(_07956_),
    .B(_03712_),
    .Y(_01740_));
 sky130_fd_sc_hd__nor2_1 _16537_ (.A(_07965_),
    .B(_03712_),
    .Y(_01741_));
 sky130_fd_sc_hd__nor2_1 _16538_ (.A(_07974_),
    .B(_03712_),
    .Y(_01742_));
 sky130_fd_sc_hd__nor2_1 _16539_ (.A(_07981_),
    .B(_03712_),
    .Y(_01743_));
 sky130_fd_sc_hd__nor2_1 _16540_ (.A(_07989_),
    .B(_03712_),
    .Y(_01744_));
 sky130_fd_sc_hd__nand2_1 _16541_ (.A(_05369_),
    .B(_08431_),
    .Y(_03716_));
 sky130_fd_sc_hd__nor2_1 _16543_ (.A(_07572_),
    .B(_03716_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor2_1 _16544_ (.A(_07660_),
    .B(_03716_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _16545_ (.A(_07669_),
    .B(_03716_),
    .Y(_01747_));
 sky130_fd_sc_hd__nor2_1 _16546_ (.A(_07677_),
    .B(_03716_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _16547_ (.A(_07689_),
    .B(_03716_),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_1 _16548_ (.A(_07703_),
    .B(_03716_),
    .Y(_01750_));
 sky130_fd_sc_hd__nor2_1 _16549_ (.A(_07709_),
    .B(_03716_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor2_1 _16550_ (.A(_07715_),
    .B(_03716_),
    .Y(_01752_));
 sky130_fd_sc_hd__nor2_1 _16551_ (.A(_07731_),
    .B(_03716_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_1 _16552_ (.A(_07745_),
    .B(_03716_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _16554_ (.A(_07752_),
    .B(_03716_),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_1 _16555_ (.A(_07577_),
    .B(_03716_),
    .Y(_01756_));
 sky130_fd_sc_hd__nor2_1 _16556_ (.A(_07766_),
    .B(_03716_),
    .Y(_01757_));
 sky130_fd_sc_hd__nor2_1 _16557_ (.A(_07777_),
    .B(_03716_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _16558_ (.A(_07786_),
    .B(_03716_),
    .Y(_01759_));
 sky130_fd_sc_hd__nor2_1 _16559_ (.A(_07800_),
    .B(_03716_),
    .Y(_01760_));
 sky130_fd_sc_hd__nor2_1 _16560_ (.A(_07809_),
    .B(_03716_),
    .Y(_01761_));
 sky130_fd_sc_hd__nor2_1 _16561_ (.A(_07818_),
    .B(_03716_),
    .Y(_01762_));
 sky130_fd_sc_hd__nor2_1 _16562_ (.A(_07831_),
    .B(_03716_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _16563_ (.A(_07843_),
    .B(_03716_),
    .Y(_01764_));
 sky130_fd_sc_hd__nor2_1 _16565_ (.A(_07850_),
    .B(_03716_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_1 _16566_ (.A(_03491_),
    .B(_03716_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor2_1 _16567_ (.A(_07581_),
    .B(_03716_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _16568_ (.A(_07873_),
    .B(_03716_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _16569_ (.A(_07925_),
    .B(_03716_),
    .Y(_01769_));
 sky130_fd_sc_hd__nor2_1 _16570_ (.A(_07588_),
    .B(_03716_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor2_1 _16571_ (.A(_07601_),
    .B(_03716_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _16572_ (.A(_07610_),
    .B(_03716_),
    .Y(_01772_));
 sky130_fd_sc_hd__nor2_1 _16573_ (.A(_07620_),
    .B(_03716_),
    .Y(_01773_));
 sky130_fd_sc_hd__nor2_1 _16574_ (.A(_07628_),
    .B(_03716_),
    .Y(_01774_));
 sky130_fd_sc_hd__nor2_1 _16575_ (.A(_07635_),
    .B(_03716_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _16576_ (.A(_07646_),
    .B(_03716_),
    .Y(_01776_));
 sky130_fd_sc_hd__nand2_1 _16577_ (.A(_05424_),
    .B(_08803_),
    .Y(_03720_));
 sky130_fd_sc_hd__nor2_1 _16579_ (.A(_07930_),
    .B(_03720_),
    .Y(_01777_));
 sky130_fd_sc_hd__nor2_1 _16580_ (.A(_08006_),
    .B(_03720_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _16581_ (.A(_08018_),
    .B(_03720_),
    .Y(_01779_));
 sky130_fd_sc_hd__nor2_1 _16582_ (.A(_08025_),
    .B(_03720_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _16583_ (.A(_08031_),
    .B(_03720_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _16584_ (.A(_08039_),
    .B(_03720_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor2_1 _16585_ (.A(_08051_),
    .B(_03720_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_1 _16586_ (.A(_08064_),
    .B(_03720_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _16587_ (.A(_08071_),
    .B(_03720_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _16588_ (.A(_08082_),
    .B(_03720_),
    .Y(_01786_));
 sky130_fd_sc_hd__nor2_1 _16590_ (.A(_08091_),
    .B(_03720_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _16591_ (.A(_07934_),
    .B(_03720_),
    .Y(_01788_));
 sky130_fd_sc_hd__nor2_1 _16592_ (.A(_08102_),
    .B(_03720_),
    .Y(_01789_));
 sky130_fd_sc_hd__nor2_1 _16593_ (.A(_08114_),
    .B(_03720_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor2_1 _16594_ (.A(_08125_),
    .B(_03720_),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _16595_ (.A(_08142_),
    .B(_03720_),
    .Y(_01792_));
 sky130_fd_sc_hd__nor2_1 _16596_ (.A(_08152_),
    .B(_03720_),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _16597_ (.A(_08160_),
    .B(_03720_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _16598_ (.A(_08171_),
    .B(_03720_),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_1 _16599_ (.A(_08184_),
    .B(_03720_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _16601_ (.A(_08204_),
    .B(_03720_),
    .Y(_01797_));
 sky130_fd_sc_hd__nor2_1 _16602_ (.A(_08209_),
    .B(_03720_),
    .Y(_01798_));
 sky130_fd_sc_hd__nor2_1 _16603_ (.A(_07937_),
    .B(_03720_),
    .Y(_01799_));
 sky130_fd_sc_hd__nor2_1 _16604_ (.A(_08221_),
    .B(_03720_),
    .Y(_01800_));
 sky130_fd_sc_hd__nor2_1 _16605_ (.A(_08254_),
    .B(_03720_),
    .Y(_01801_));
 sky130_fd_sc_hd__nor2_1 _16606_ (.A(_07942_),
    .B(_03720_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _16607_ (.A(_07949_),
    .B(_03720_),
    .Y(_01803_));
 sky130_fd_sc_hd__nor2_1 _16608_ (.A(_07956_),
    .B(_03720_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _16609_ (.A(_07965_),
    .B(_03720_),
    .Y(_01805_));
 sky130_fd_sc_hd__nor2_1 _16610_ (.A(_07974_),
    .B(_03720_),
    .Y(_01806_));
 sky130_fd_sc_hd__nor2_1 _16611_ (.A(_07981_),
    .B(_03720_),
    .Y(_01807_));
 sky130_fd_sc_hd__nor2_1 _16612_ (.A(_07989_),
    .B(_03720_),
    .Y(_01808_));
 sky130_fd_sc_hd__nand2_1 _16613_ (.A(_05376_),
    .B(_07566_),
    .Y(_03724_));
 sky130_fd_sc_hd__nor2_1 _16615_ (.A(_07572_),
    .B(_03724_),
    .Y(_01809_));
 sky130_fd_sc_hd__nor2_1 _16616_ (.A(_07660_),
    .B(_03724_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _16617_ (.A(_07669_),
    .B(_03724_),
    .Y(_01811_));
 sky130_fd_sc_hd__nor2_1 _16618_ (.A(_07677_),
    .B(_03724_),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_1 _16619_ (.A(_07689_),
    .B(_03724_),
    .Y(_01813_));
 sky130_fd_sc_hd__nor2_1 _16620_ (.A(_07703_),
    .B(_03724_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_1 _16621_ (.A(_07709_),
    .B(_03724_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _16622_ (.A(_07715_),
    .B(_03724_),
    .Y(_01816_));
 sky130_fd_sc_hd__nor2_1 _16623_ (.A(_07731_),
    .B(_03724_),
    .Y(_01817_));
 sky130_fd_sc_hd__nor2_1 _16624_ (.A(_07745_),
    .B(_03724_),
    .Y(_01818_));
 sky130_fd_sc_hd__nor2_1 _16626_ (.A(_07752_),
    .B(_03724_),
    .Y(_01819_));
 sky130_fd_sc_hd__nor2_1 _16627_ (.A(_07577_),
    .B(_03724_),
    .Y(_01820_));
 sky130_fd_sc_hd__nor2_1 _16628_ (.A(_07766_),
    .B(_03724_),
    .Y(_01821_));
 sky130_fd_sc_hd__nor2_1 _16629_ (.A(_07777_),
    .B(_03724_),
    .Y(_01822_));
 sky130_fd_sc_hd__nor2_1 _16630_ (.A(_07786_),
    .B(_03724_),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_1 _16631_ (.A(_07800_),
    .B(_03724_),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _16632_ (.A(_07809_),
    .B(_03724_),
    .Y(_01825_));
 sky130_fd_sc_hd__nor2_1 _16633_ (.A(_07818_),
    .B(_03724_),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _16634_ (.A(_07831_),
    .B(_03724_),
    .Y(_01827_));
 sky130_fd_sc_hd__nor2_1 _16635_ (.A(_07843_),
    .B(_03724_),
    .Y(_01828_));
 sky130_fd_sc_hd__nor2_1 _16637_ (.A(_07850_),
    .B(_03724_),
    .Y(_01829_));
 sky130_fd_sc_hd__nor2_1 _16638_ (.A(_03491_),
    .B(_03724_),
    .Y(_01830_));
 sky130_fd_sc_hd__nor2_1 _16639_ (.A(_07581_),
    .B(_03724_),
    .Y(_01831_));
 sky130_fd_sc_hd__nor2_1 _16640_ (.A(_07873_),
    .B(_03724_),
    .Y(_01832_));
 sky130_fd_sc_hd__nor2_1 _16641_ (.A(_07925_),
    .B(_03724_),
    .Y(_01833_));
 sky130_fd_sc_hd__nor2_1 _16642_ (.A(_07588_),
    .B(_03724_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _16643_ (.A(_07601_),
    .B(_03724_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor2_1 _16644_ (.A(_07610_),
    .B(_03724_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _16645_ (.A(_07620_),
    .B(_03724_),
    .Y(_01837_));
 sky130_fd_sc_hd__nor2_1 _16646_ (.A(_07628_),
    .B(_03724_),
    .Y(_01838_));
 sky130_fd_sc_hd__nor2_1 _16647_ (.A(_07635_),
    .B(_03724_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _16648_ (.A(_07646_),
    .B(_03724_),
    .Y(_01840_));
 sky130_fd_sc_hd__nand2_1 _16649_ (.A(_05431_),
    .B(_07927_),
    .Y(_03728_));
 sky130_fd_sc_hd__nor2_1 _16651_ (.A(_07930_),
    .B(_03728_),
    .Y(_01841_));
 sky130_fd_sc_hd__nor2_1 _16652_ (.A(_08006_),
    .B(_03728_),
    .Y(_01842_));
 sky130_fd_sc_hd__nor2_1 _16653_ (.A(_08018_),
    .B(_03728_),
    .Y(_01843_));
 sky130_fd_sc_hd__nor2_1 _16654_ (.A(_08025_),
    .B(_03728_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _16655_ (.A(_08031_),
    .B(_03728_),
    .Y(_01845_));
 sky130_fd_sc_hd__nor2_1 _16656_ (.A(_08039_),
    .B(_03728_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_1 _16657_ (.A(_08051_),
    .B(_03728_),
    .Y(_01847_));
 sky130_fd_sc_hd__nor2_1 _16658_ (.A(_08064_),
    .B(_03728_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_1 _16659_ (.A(_08071_),
    .B(_03728_),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _16660_ (.A(_08082_),
    .B(_03728_),
    .Y(_01850_));
 sky130_fd_sc_hd__nor2_1 _16662_ (.A(_08091_),
    .B(_03728_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor2_1 _16663_ (.A(_07934_),
    .B(_03728_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _16664_ (.A(_08102_),
    .B(_03728_),
    .Y(_01853_));
 sky130_fd_sc_hd__nor2_1 _16665_ (.A(_08114_),
    .B(_03728_),
    .Y(_01854_));
 sky130_fd_sc_hd__nor2_1 _16666_ (.A(_08125_),
    .B(_03728_),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_1 _16667_ (.A(_08142_),
    .B(_03728_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _16668_ (.A(_08152_),
    .B(_03728_),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _16669_ (.A(_08160_),
    .B(_03728_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _16670_ (.A(_08171_),
    .B(_03728_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _16671_ (.A(_08184_),
    .B(_03728_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor2_1 _16673_ (.A(_08204_),
    .B(_03728_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _16674_ (.A(_08209_),
    .B(_03728_),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_1 _16675_ (.A(_07937_),
    .B(_03728_),
    .Y(_01863_));
 sky130_fd_sc_hd__nor2_1 _16676_ (.A(_08221_),
    .B(_03728_),
    .Y(_01864_));
 sky130_fd_sc_hd__nor2_1 _16677_ (.A(_08254_),
    .B(_03728_),
    .Y(_01865_));
 sky130_fd_sc_hd__nor2_1 _16678_ (.A(_07942_),
    .B(_03728_),
    .Y(_01866_));
 sky130_fd_sc_hd__nor2_1 _16679_ (.A(_07949_),
    .B(_03728_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor2_1 _16680_ (.A(_07956_),
    .B(_03728_),
    .Y(_01868_));
 sky130_fd_sc_hd__nor2_1 _16681_ (.A(_07965_),
    .B(_03728_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _16682_ (.A(_07974_),
    .B(_03728_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _16683_ (.A(_07981_),
    .B(_03728_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _16684_ (.A(_07989_),
    .B(_03728_),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_1 _16685_ (.A(_05376_),
    .B(_08257_),
    .Y(_03732_));
 sky130_fd_sc_hd__nor2_1 _16687_ (.A(_07572_),
    .B(_03732_),
    .Y(_01873_));
 sky130_fd_sc_hd__nor2_1 _16688_ (.A(_07660_),
    .B(_03732_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _16689_ (.A(_07669_),
    .B(_03732_),
    .Y(_01875_));
 sky130_fd_sc_hd__nor2_1 _16690_ (.A(_07677_),
    .B(_03732_),
    .Y(_01876_));
 sky130_fd_sc_hd__nor2_1 _16691_ (.A(_07689_),
    .B(_03732_),
    .Y(_01877_));
 sky130_fd_sc_hd__nor2_1 _16692_ (.A(_07703_),
    .B(_03732_),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _16693_ (.A(_07709_),
    .B(_03732_),
    .Y(_01879_));
 sky130_fd_sc_hd__nor2_1 _16694_ (.A(_07715_),
    .B(_03732_),
    .Y(_01880_));
 sky130_fd_sc_hd__nor2_1 _16695_ (.A(_07731_),
    .B(_03732_),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_1 _16696_ (.A(_07745_),
    .B(_03732_),
    .Y(_01882_));
 sky130_fd_sc_hd__nor2_1 _16698_ (.A(_07752_),
    .B(_03732_),
    .Y(_01883_));
 sky130_fd_sc_hd__nor2_1 _16699_ (.A(_07577_),
    .B(_03732_),
    .Y(_01884_));
 sky130_fd_sc_hd__nor2_1 _16700_ (.A(_07766_),
    .B(_03732_),
    .Y(_01885_));
 sky130_fd_sc_hd__nor2_1 _16701_ (.A(_07777_),
    .B(_03732_),
    .Y(_01886_));
 sky130_fd_sc_hd__nor2_1 _16702_ (.A(_07786_),
    .B(_03732_),
    .Y(_01887_));
 sky130_fd_sc_hd__nor2_1 _16703_ (.A(_07800_),
    .B(_03732_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor2_1 _16704_ (.A(_07809_),
    .B(_03732_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor2_1 _16705_ (.A(_07818_),
    .B(_03732_),
    .Y(_01890_));
 sky130_fd_sc_hd__nor2_1 _16706_ (.A(_07831_),
    .B(_03732_),
    .Y(_01891_));
 sky130_fd_sc_hd__nor2_1 _16707_ (.A(_07843_),
    .B(_03732_),
    .Y(_01892_));
 sky130_fd_sc_hd__nor2_1 _16709_ (.A(_07850_),
    .B(_03732_),
    .Y(_01893_));
 sky130_fd_sc_hd__nor2_1 _16710_ (.A(_03491_),
    .B(_03732_),
    .Y(_01894_));
 sky130_fd_sc_hd__nor2_1 _16711_ (.A(_07581_),
    .B(_03732_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _16712_ (.A(_07873_),
    .B(_03732_),
    .Y(_01896_));
 sky130_fd_sc_hd__nor2_1 _16713_ (.A(_07925_),
    .B(_03732_),
    .Y(_01897_));
 sky130_fd_sc_hd__nor2_1 _16714_ (.A(_07588_),
    .B(_03732_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _16715_ (.A(_07601_),
    .B(_03732_),
    .Y(_01899_));
 sky130_fd_sc_hd__nor2_1 _16716_ (.A(_07610_),
    .B(_03732_),
    .Y(_01900_));
 sky130_fd_sc_hd__nor2_1 _16717_ (.A(_07620_),
    .B(_03732_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _16718_ (.A(_07628_),
    .B(_03732_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _16719_ (.A(_07635_),
    .B(_03732_),
    .Y(_01903_));
 sky130_fd_sc_hd__nor2_1 _16720_ (.A(_07646_),
    .B(_03732_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _16721_ (.A(_05431_),
    .B(_08304_),
    .Y(_03736_));
 sky130_fd_sc_hd__nor2_1 _16723_ (.A(_07930_),
    .B(_03736_),
    .Y(_01905_));
 sky130_fd_sc_hd__nor2_1 _16724_ (.A(_08006_),
    .B(_03736_),
    .Y(_01906_));
 sky130_fd_sc_hd__nor2_1 _16725_ (.A(_08018_),
    .B(_03736_),
    .Y(_01907_));
 sky130_fd_sc_hd__nor2_1 _16726_ (.A(_08025_),
    .B(_03736_),
    .Y(_01908_));
 sky130_fd_sc_hd__nor2_1 _16727_ (.A(_08031_),
    .B(_03736_),
    .Y(_01909_));
 sky130_fd_sc_hd__nor2_1 _16728_ (.A(_08039_),
    .B(_03736_),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _16729_ (.A(_08051_),
    .B(_03736_),
    .Y(_01911_));
 sky130_fd_sc_hd__nor2_1 _16730_ (.A(_08064_),
    .B(_03736_),
    .Y(_01912_));
 sky130_fd_sc_hd__nor2_1 _16731_ (.A(_08071_),
    .B(_03736_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_08082_),
    .B(_03736_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _16734_ (.A(_08091_),
    .B(_03736_),
    .Y(_01915_));
 sky130_fd_sc_hd__nor2_1 _16735_ (.A(_07934_),
    .B(_03736_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _16736_ (.A(_08102_),
    .B(_03736_),
    .Y(_01917_));
 sky130_fd_sc_hd__nor2_1 _16737_ (.A(_08114_),
    .B(_03736_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _16738_ (.A(_08125_),
    .B(_03736_),
    .Y(_01919_));
 sky130_fd_sc_hd__nor2_1 _16739_ (.A(_08142_),
    .B(_03736_),
    .Y(_01920_));
 sky130_fd_sc_hd__nor2_1 _16740_ (.A(_08152_),
    .B(_03736_),
    .Y(_01921_));
 sky130_fd_sc_hd__nor2_1 _16741_ (.A(_08160_),
    .B(_03736_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _16742_ (.A(_08171_),
    .B(_03736_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_1 _16743_ (.A(_08184_),
    .B(_03736_),
    .Y(_01924_));
 sky130_fd_sc_hd__nor2_1 _16745_ (.A(_08204_),
    .B(_03736_),
    .Y(_01925_));
 sky130_fd_sc_hd__nor2_1 _16746_ (.A(_08209_),
    .B(_03736_),
    .Y(_01926_));
 sky130_fd_sc_hd__nor2_1 _16747_ (.A(_07937_),
    .B(_03736_),
    .Y(_01927_));
 sky130_fd_sc_hd__nor2_1 _16748_ (.A(_08221_),
    .B(_03736_),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _16749_ (.A(_08254_),
    .B(_03736_),
    .Y(_01929_));
 sky130_fd_sc_hd__nor2_1 _16750_ (.A(_07942_),
    .B(_03736_),
    .Y(_01930_));
 sky130_fd_sc_hd__nor2_1 _16751_ (.A(_07949_),
    .B(_03736_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _16752_ (.A(_07956_),
    .B(_03736_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_1 _16753_ (.A(_07965_),
    .B(_03736_),
    .Y(_01933_));
 sky130_fd_sc_hd__nor2_1 _16754_ (.A(_07974_),
    .B(_03736_),
    .Y(_01934_));
 sky130_fd_sc_hd__nor2_1 _16755_ (.A(_07981_),
    .B(_03736_),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_1 _16756_ (.A(_07989_),
    .B(_03736_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_1 _16757_ (.A(_05376_),
    .B(_08346_),
    .Y(_03740_));
 sky130_fd_sc_hd__nor2_1 _16759_ (.A(_07572_),
    .B(_03740_),
    .Y(_01937_));
 sky130_fd_sc_hd__nor2_1 _16760_ (.A(_07660_),
    .B(_03740_),
    .Y(_01938_));
 sky130_fd_sc_hd__nor2_1 _16761_ (.A(_07669_),
    .B(_03740_),
    .Y(_01939_));
 sky130_fd_sc_hd__nor2_1 _16762_ (.A(_07677_),
    .B(_03740_),
    .Y(_01940_));
 sky130_fd_sc_hd__nor2_1 _16763_ (.A(_07689_),
    .B(_03740_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor2_1 _16764_ (.A(_07703_),
    .B(_03740_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_1 _16765_ (.A(_07709_),
    .B(_03740_),
    .Y(_01943_));
 sky130_fd_sc_hd__nor2_1 _16766_ (.A(_07715_),
    .B(_03740_),
    .Y(_01944_));
 sky130_fd_sc_hd__nor2_1 _16767_ (.A(_07731_),
    .B(_03740_),
    .Y(_01945_));
 sky130_fd_sc_hd__nor2_1 _16768_ (.A(_07745_),
    .B(_03740_),
    .Y(_01946_));
 sky130_fd_sc_hd__nor2_1 _16770_ (.A(_07752_),
    .B(_03740_),
    .Y(_01947_));
 sky130_fd_sc_hd__nor2_1 _16771_ (.A(_07577_),
    .B(_03740_),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_1 _16772_ (.A(_07766_),
    .B(_03740_),
    .Y(_01949_));
 sky130_fd_sc_hd__nor2_1 _16773_ (.A(_07777_),
    .B(_03740_),
    .Y(_01950_));
 sky130_fd_sc_hd__nor2_1 _16774_ (.A(_07786_),
    .B(_03740_),
    .Y(_01951_));
 sky130_fd_sc_hd__nor2_1 _16775_ (.A(_07800_),
    .B(_03740_),
    .Y(_01952_));
 sky130_fd_sc_hd__nor2_1 _16776_ (.A(_07809_),
    .B(_03740_),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _16777_ (.A(_07818_),
    .B(_03740_),
    .Y(_01954_));
 sky130_fd_sc_hd__nor2_1 _16778_ (.A(_07831_),
    .B(_03740_),
    .Y(_01955_));
 sky130_fd_sc_hd__nor2_1 _16779_ (.A(_07843_),
    .B(_03740_),
    .Y(_01956_));
 sky130_fd_sc_hd__nor2_1 _16781_ (.A(_07850_),
    .B(_03740_),
    .Y(_01957_));
 sky130_fd_sc_hd__nor2_1 _16782_ (.A(_03491_),
    .B(_03740_),
    .Y(_01958_));
 sky130_fd_sc_hd__nor2_1 _16783_ (.A(_07581_),
    .B(_03740_),
    .Y(_01959_));
 sky130_fd_sc_hd__nor2_1 _16784_ (.A(_07873_),
    .B(_03740_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2_1 _16785_ (.A(_07925_),
    .B(_03740_),
    .Y(_01961_));
 sky130_fd_sc_hd__nor2_1 _16786_ (.A(_07588_),
    .B(_03740_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _16787_ (.A(_07601_),
    .B(_03740_),
    .Y(_01963_));
 sky130_fd_sc_hd__nor2_1 _16788_ (.A(_07610_),
    .B(_03740_),
    .Y(_01964_));
 sky130_fd_sc_hd__nor2_1 _16789_ (.A(_07620_),
    .B(_03740_),
    .Y(_01965_));
 sky130_fd_sc_hd__nor2_1 _16790_ (.A(_07628_),
    .B(_03740_),
    .Y(_01966_));
 sky130_fd_sc_hd__nor2_1 _16791_ (.A(_07635_),
    .B(_03740_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _16792_ (.A(_07646_),
    .B(_03740_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _16793_ (.A(_05431_),
    .B(_08390_),
    .Y(_03744_));
 sky130_fd_sc_hd__nor2_1 _16795_ (.A(_07930_),
    .B(_03744_),
    .Y(_01969_));
 sky130_fd_sc_hd__nor2_1 _16796_ (.A(_08006_),
    .B(_03744_),
    .Y(_01970_));
 sky130_fd_sc_hd__nor2_1 _16797_ (.A(_08018_),
    .B(_03744_),
    .Y(_01971_));
 sky130_fd_sc_hd__nor2_1 _16798_ (.A(_08025_),
    .B(_03744_),
    .Y(_01972_));
 sky130_fd_sc_hd__nor2_1 _16799_ (.A(_08031_),
    .B(_03744_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_1 _16800_ (.A(_08039_),
    .B(_03744_),
    .Y(_01974_));
 sky130_fd_sc_hd__nor2_1 _16801_ (.A(_08051_),
    .B(_03744_),
    .Y(_01975_));
 sky130_fd_sc_hd__nor2_1 _16802_ (.A(_08064_),
    .B(_03744_),
    .Y(_01976_));
 sky130_fd_sc_hd__nor2_1 _16803_ (.A(_08071_),
    .B(_03744_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_1 _16804_ (.A(_08082_),
    .B(_03744_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _16806_ (.A(_08091_),
    .B(_03744_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _16807_ (.A(_07934_),
    .B(_03744_),
    .Y(_01980_));
 sky130_fd_sc_hd__nor2_1 _16808_ (.A(_08102_),
    .B(_03744_),
    .Y(_01981_));
 sky130_fd_sc_hd__nor2_1 _16809_ (.A(_08114_),
    .B(_03744_),
    .Y(_01982_));
 sky130_fd_sc_hd__nor2_1 _16810_ (.A(_08125_),
    .B(_03744_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _16811_ (.A(_08142_),
    .B(_03744_),
    .Y(_01984_));
 sky130_fd_sc_hd__nor2_1 _16812_ (.A(_08152_),
    .B(_03744_),
    .Y(_01985_));
 sky130_fd_sc_hd__nor2_1 _16813_ (.A(_08160_),
    .B(_03744_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_1 _16814_ (.A(_08171_),
    .B(_03744_),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2_1 _16815_ (.A(_08184_),
    .B(_03744_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor2_1 _16817_ (.A(_08204_),
    .B(_03744_),
    .Y(_01989_));
 sky130_fd_sc_hd__nor2_1 _16818_ (.A(_08209_),
    .B(_03744_),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_1 _16819_ (.A(_07937_),
    .B(_03744_),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_1 _16820_ (.A(_08221_),
    .B(_03744_),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _16821_ (.A(_08254_),
    .B(_03744_),
    .Y(_01993_));
 sky130_fd_sc_hd__nor2_1 _16822_ (.A(_07942_),
    .B(_03744_),
    .Y(_01994_));
 sky130_fd_sc_hd__nor2_1 _16823_ (.A(_07949_),
    .B(_03744_),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_1 _16824_ (.A(_07956_),
    .B(_03744_),
    .Y(_01996_));
 sky130_fd_sc_hd__nor2_1 _16825_ (.A(_07965_),
    .B(_03744_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _16826_ (.A(_07974_),
    .B(_03744_),
    .Y(_01998_));
 sky130_fd_sc_hd__nor2_1 _16827_ (.A(_07981_),
    .B(_03744_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor2_1 _16828_ (.A(_07989_),
    .B(_03744_),
    .Y(_02000_));
 sky130_fd_sc_hd__nand2_1 _16829_ (.A(_05376_),
    .B(_08431_),
    .Y(_03748_));
 sky130_fd_sc_hd__nor2_1 _16831_ (.A(_07572_),
    .B(_03748_),
    .Y(_02001_));
 sky130_fd_sc_hd__nor2_1 _16832_ (.A(_07660_),
    .B(_03748_),
    .Y(_02002_));
 sky130_fd_sc_hd__nor2_1 _16833_ (.A(_07669_),
    .B(_03748_),
    .Y(_02003_));
 sky130_fd_sc_hd__nor2_1 _16834_ (.A(_07677_),
    .B(_03748_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_1 _16835_ (.A(_07689_),
    .B(_03748_),
    .Y(_02005_));
 sky130_fd_sc_hd__nor2_1 _16836_ (.A(_07703_),
    .B(_03748_),
    .Y(_02006_));
 sky130_fd_sc_hd__nor2_1 _16837_ (.A(_07709_),
    .B(_03748_),
    .Y(_02007_));
 sky130_fd_sc_hd__nor2_1 _16838_ (.A(_07715_),
    .B(_03748_),
    .Y(_02008_));
 sky130_fd_sc_hd__nor2_1 _16839_ (.A(_07731_),
    .B(_03748_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _16840_ (.A(_07745_),
    .B(_03748_),
    .Y(_02010_));
 sky130_fd_sc_hd__nor2_1 _16842_ (.A(_07752_),
    .B(_03748_),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _16843_ (.A(_07577_),
    .B(_03748_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_1 _16844_ (.A(_07766_),
    .B(_03748_),
    .Y(_02013_));
 sky130_fd_sc_hd__nor2_1 _16845_ (.A(_07777_),
    .B(_03748_),
    .Y(_02014_));
 sky130_fd_sc_hd__nor2_1 _16846_ (.A(_07786_),
    .B(_03748_),
    .Y(_02015_));
 sky130_fd_sc_hd__nor2_1 _16847_ (.A(_07800_),
    .B(_03748_),
    .Y(_02016_));
 sky130_fd_sc_hd__nor2_1 _16848_ (.A(_07809_),
    .B(_03748_),
    .Y(_02017_));
 sky130_fd_sc_hd__nor2_1 _16849_ (.A(_07818_),
    .B(_03748_),
    .Y(_02018_));
 sky130_fd_sc_hd__nor2_1 _16850_ (.A(_07831_),
    .B(_03748_),
    .Y(_02019_));
 sky130_fd_sc_hd__nor2_1 _16851_ (.A(_07843_),
    .B(_03748_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _16853_ (.A(_07850_),
    .B(_03748_),
    .Y(_02021_));
 sky130_fd_sc_hd__nor2_1 _16854_ (.A(_03491_),
    .B(_03748_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_1 _16855_ (.A(_07581_),
    .B(_03748_),
    .Y(_02023_));
 sky130_fd_sc_hd__nor2_1 _16856_ (.A(_07873_),
    .B(_03748_),
    .Y(_02024_));
 sky130_fd_sc_hd__nor2_1 _16857_ (.A(_07925_),
    .B(_03748_),
    .Y(_02025_));
 sky130_fd_sc_hd__nor2_1 _16858_ (.A(_07588_),
    .B(_03748_),
    .Y(_02026_));
 sky130_fd_sc_hd__nor2_1 _16859_ (.A(_07601_),
    .B(_03748_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _16860_ (.A(_07610_),
    .B(_03748_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _16861_ (.A(_07620_),
    .B(_03748_),
    .Y(_02029_));
 sky130_fd_sc_hd__nor2_1 _16862_ (.A(_07628_),
    .B(_03748_),
    .Y(_02030_));
 sky130_fd_sc_hd__nor2_1 _16863_ (.A(_07635_),
    .B(_03748_),
    .Y(_02031_));
 sky130_fd_sc_hd__nor2_1 _16864_ (.A(_07646_),
    .B(_03748_),
    .Y(_02032_));
 sky130_fd_sc_hd__or3_1 _16865_ (.A(reset),
    .B(_05422_),
    .C(_05399_),
    .X(_03752_));
 sky130_fd_sc_hd__nor2_1 _16868_ (.A(_07930_),
    .B(_03752_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_1 _16869_ (.A(_08006_),
    .B(_03752_),
    .Y(_02034_));
 sky130_fd_sc_hd__nor2_1 _16870_ (.A(_08018_),
    .B(_03752_),
    .Y(_02035_));
 sky130_fd_sc_hd__nor2_1 _16871_ (.A(_08025_),
    .B(_03752_),
    .Y(_02036_));
 sky130_fd_sc_hd__nor2_1 _16872_ (.A(_08031_),
    .B(_03752_),
    .Y(_02037_));
 sky130_fd_sc_hd__nor2_1 _16873_ (.A(_08039_),
    .B(_03752_),
    .Y(_02038_));
 sky130_fd_sc_hd__nor2_1 _16874_ (.A(_08051_),
    .B(_03752_),
    .Y(_02039_));
 sky130_fd_sc_hd__nor2_1 _16875_ (.A(_08064_),
    .B(_03752_),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _16876_ (.A(_08071_),
    .B(_03752_),
    .Y(_02041_));
 sky130_fd_sc_hd__nor2_1 _16877_ (.A(_08082_),
    .B(_03752_),
    .Y(_02042_));
 sky130_fd_sc_hd__nor2_1 _16879_ (.A(_08091_),
    .B(_03752_),
    .Y(_02043_));
 sky130_fd_sc_hd__nor2_1 _16880_ (.A(_07934_),
    .B(_03752_),
    .Y(_02044_));
 sky130_fd_sc_hd__nor2_1 _16881_ (.A(_08102_),
    .B(_03752_),
    .Y(_02045_));
 sky130_fd_sc_hd__nor2_1 _16882_ (.A(_08114_),
    .B(_03752_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_1 _16883_ (.A(_08125_),
    .B(_03752_),
    .Y(_02047_));
 sky130_fd_sc_hd__nor2_1 _16884_ (.A(_08142_),
    .B(_03752_),
    .Y(_02048_));
 sky130_fd_sc_hd__nor2_1 _16885_ (.A(_08152_),
    .B(_03752_),
    .Y(_02049_));
 sky130_fd_sc_hd__nor2_1 _16886_ (.A(_08160_),
    .B(_03752_),
    .Y(_02050_));
 sky130_fd_sc_hd__nor2_1 _16887_ (.A(_08171_),
    .B(_03752_),
    .Y(_02051_));
 sky130_fd_sc_hd__nor2_1 _16888_ (.A(_08184_),
    .B(_03752_),
    .Y(_02052_));
 sky130_fd_sc_hd__nor2_1 _16890_ (.A(_08204_),
    .B(_03752_),
    .Y(_02053_));
 sky130_fd_sc_hd__nor2_1 _16891_ (.A(_08209_),
    .B(_03752_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _16892_ (.A(_07937_),
    .B(_03752_),
    .Y(_02055_));
 sky130_fd_sc_hd__nor2_1 _16893_ (.A(_08221_),
    .B(_03752_),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_1 _16894_ (.A(_08254_),
    .B(_03752_),
    .Y(_02057_));
 sky130_fd_sc_hd__nor2_1 _16895_ (.A(_07942_),
    .B(_03752_),
    .Y(_02058_));
 sky130_fd_sc_hd__nor2_1 _16896_ (.A(_07949_),
    .B(_03752_),
    .Y(_02059_));
 sky130_fd_sc_hd__nor2_1 _16897_ (.A(_07956_),
    .B(_03752_),
    .Y(_02060_));
 sky130_fd_sc_hd__nor2_1 _16898_ (.A(_07965_),
    .B(_03752_),
    .Y(_02061_));
 sky130_fd_sc_hd__nor2_1 _16899_ (.A(_07974_),
    .B(_03752_),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _16900_ (.A(_07981_),
    .B(_03752_),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_1 _16901_ (.A(_07989_),
    .B(_03752_),
    .Y(_02064_));
 sky130_fd_sc_hd__nand2_1 _16902_ (.A(_05383_),
    .B(_07566_),
    .Y(_03757_));
 sky130_fd_sc_hd__nor2_1 _16904_ (.A(_07572_),
    .B(_03757_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor2_1 _16905_ (.A(_07660_),
    .B(_03757_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _16906_ (.A(_07669_),
    .B(_03757_),
    .Y(_02067_));
 sky130_fd_sc_hd__nor2_1 _16907_ (.A(_07677_),
    .B(_03757_),
    .Y(_02068_));
 sky130_fd_sc_hd__nor2_1 _16908_ (.A(_07689_),
    .B(_03757_),
    .Y(_02069_));
 sky130_fd_sc_hd__nor2_1 _16909_ (.A(_07703_),
    .B(_03757_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_1 _16910_ (.A(_07709_),
    .B(_03757_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_1 _16911_ (.A(_07715_),
    .B(_03757_),
    .Y(_02072_));
 sky130_fd_sc_hd__nor2_1 _16912_ (.A(_07731_),
    .B(_03757_),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_1 _16913_ (.A(_07745_),
    .B(_03757_),
    .Y(_02074_));
 sky130_fd_sc_hd__nor2_1 _16915_ (.A(_07752_),
    .B(_03757_),
    .Y(_02075_));
 sky130_fd_sc_hd__nor2_1 _16916_ (.A(_07577_),
    .B(_03757_),
    .Y(_02076_));
 sky130_fd_sc_hd__nor2_1 _16917_ (.A(_07766_),
    .B(_03757_),
    .Y(_02077_));
 sky130_fd_sc_hd__nor2_1 _16918_ (.A(_07777_),
    .B(_03757_),
    .Y(_02078_));
 sky130_fd_sc_hd__nor2_1 _16919_ (.A(_07786_),
    .B(_03757_),
    .Y(_02079_));
 sky130_fd_sc_hd__nor2_1 _16920_ (.A(_07800_),
    .B(_03757_),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _16921_ (.A(_07809_),
    .B(_03757_),
    .Y(_02081_));
 sky130_fd_sc_hd__nor2_1 _16922_ (.A(_07818_),
    .B(_03757_),
    .Y(_02082_));
 sky130_fd_sc_hd__nor2_1 _16923_ (.A(_07831_),
    .B(_03757_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_1 _16924_ (.A(_07843_),
    .B(_03757_),
    .Y(_02084_));
 sky130_fd_sc_hd__nor2_1 _16926_ (.A(_07850_),
    .B(_03757_),
    .Y(_02085_));
 sky130_fd_sc_hd__nor2_1 _16927_ (.A(_03491_),
    .B(_03757_),
    .Y(_02086_));
 sky130_fd_sc_hd__nor2_1 _16928_ (.A(_07581_),
    .B(_03757_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor2_1 _16929_ (.A(_07873_),
    .B(_03757_),
    .Y(_02088_));
 sky130_fd_sc_hd__nor2_1 _16930_ (.A(_07925_),
    .B(_03757_),
    .Y(_02089_));
 sky130_fd_sc_hd__nor2_1 _16931_ (.A(_07588_),
    .B(_03757_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _16932_ (.A(_07601_),
    .B(_03757_),
    .Y(_02091_));
 sky130_fd_sc_hd__nor2_1 _16933_ (.A(_07610_),
    .B(_03757_),
    .Y(_02092_));
 sky130_fd_sc_hd__nor2_1 _16934_ (.A(_07620_),
    .B(_03757_),
    .Y(_02093_));
 sky130_fd_sc_hd__nor2_1 _16935_ (.A(_07628_),
    .B(_03757_),
    .Y(_02094_));
 sky130_fd_sc_hd__nor2_1 _16936_ (.A(_07635_),
    .B(_03757_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor2_1 _16937_ (.A(_07646_),
    .B(_03757_),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_1 _16938_ (.A(_05436_),
    .B(_07927_),
    .Y(_03761_));
 sky130_fd_sc_hd__nor2_1 _16940_ (.A(_07930_),
    .B(_03761_),
    .Y(_02097_));
 sky130_fd_sc_hd__nor2_1 _16941_ (.A(_08006_),
    .B(_03761_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_1 _16942_ (.A(_08018_),
    .B(_03761_),
    .Y(_02099_));
 sky130_fd_sc_hd__nor2_1 _16943_ (.A(_08025_),
    .B(_03761_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_1 _16944_ (.A(_08031_),
    .B(_03761_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor2_1 _16945_ (.A(_08039_),
    .B(_03761_),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _16946_ (.A(_08051_),
    .B(_03761_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _16947_ (.A(_08064_),
    .B(_03761_),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _16948_ (.A(_08071_),
    .B(_03761_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _16949_ (.A(_08082_),
    .B(_03761_),
    .Y(_02106_));
 sky130_fd_sc_hd__nor2_1 _16951_ (.A(_08091_),
    .B(_03761_),
    .Y(_02107_));
 sky130_fd_sc_hd__nor2_1 _16952_ (.A(_07934_),
    .B(_03761_),
    .Y(_02108_));
 sky130_fd_sc_hd__nor2_1 _16953_ (.A(_08102_),
    .B(_03761_),
    .Y(_02109_));
 sky130_fd_sc_hd__nor2_1 _16954_ (.A(_08114_),
    .B(_03761_),
    .Y(_02110_));
 sky130_fd_sc_hd__nor2_1 _16955_ (.A(_08125_),
    .B(_03761_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor2_1 _16956_ (.A(_08142_),
    .B(_03761_),
    .Y(_02112_));
 sky130_fd_sc_hd__nor2_1 _16957_ (.A(_08152_),
    .B(_03761_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor2_1 _16958_ (.A(_08160_),
    .B(_03761_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _16959_ (.A(_08171_),
    .B(_03761_),
    .Y(_02115_));
 sky130_fd_sc_hd__nor2_1 _16960_ (.A(_08184_),
    .B(_03761_),
    .Y(_02116_));
 sky130_fd_sc_hd__nor2_1 _16962_ (.A(_08204_),
    .B(_03761_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _16963_ (.A(_08209_),
    .B(_03761_),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_1 _16964_ (.A(_07937_),
    .B(_03761_),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _16965_ (.A(_08221_),
    .B(_03761_),
    .Y(_02120_));
 sky130_fd_sc_hd__nor2_1 _16966_ (.A(_08254_),
    .B(_03761_),
    .Y(_02121_));
 sky130_fd_sc_hd__nor2_1 _16967_ (.A(_07942_),
    .B(_03761_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _16968_ (.A(_07949_),
    .B(_03761_),
    .Y(_02123_));
 sky130_fd_sc_hd__nor2_1 _16969_ (.A(_07956_),
    .B(_03761_),
    .Y(_02124_));
 sky130_fd_sc_hd__nor2_1 _16970_ (.A(_07965_),
    .B(_03761_),
    .Y(_02125_));
 sky130_fd_sc_hd__nor2_1 _16971_ (.A(_07974_),
    .B(_03761_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor2_1 _16972_ (.A(_07981_),
    .B(_03761_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _16973_ (.A(_07989_),
    .B(_03761_),
    .Y(_02128_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(_05383_),
    .B(_08257_),
    .Y(_03765_));
 sky130_fd_sc_hd__nor2_1 _16976_ (.A(_07572_),
    .B(_03765_),
    .Y(_02129_));
 sky130_fd_sc_hd__nor2_1 _16977_ (.A(_07660_),
    .B(_03765_),
    .Y(_02130_));
 sky130_fd_sc_hd__nor2_1 _16978_ (.A(_07669_),
    .B(_03765_),
    .Y(_02131_));
 sky130_fd_sc_hd__nor2_1 _16979_ (.A(_07677_),
    .B(_03765_),
    .Y(_02132_));
 sky130_fd_sc_hd__nor2_1 _16980_ (.A(_07689_),
    .B(_03765_),
    .Y(_02133_));
 sky130_fd_sc_hd__nor2_1 _16981_ (.A(_07703_),
    .B(_03765_),
    .Y(_02134_));
 sky130_fd_sc_hd__nor2_1 _16982_ (.A(_07709_),
    .B(_03765_),
    .Y(_02135_));
 sky130_fd_sc_hd__nor2_1 _16983_ (.A(_07715_),
    .B(_03765_),
    .Y(_02136_));
 sky130_fd_sc_hd__nor2_1 _16984_ (.A(_07731_),
    .B(_03765_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _16985_ (.A(_07745_),
    .B(_03765_),
    .Y(_02138_));
 sky130_fd_sc_hd__nor2_1 _16987_ (.A(_07752_),
    .B(_03765_),
    .Y(_02139_));
 sky130_fd_sc_hd__nor2_1 _16988_ (.A(_07577_),
    .B(_03765_),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2_1 _16989_ (.A(_07766_),
    .B(_03765_),
    .Y(_02141_));
 sky130_fd_sc_hd__nor2_1 _16990_ (.A(_07777_),
    .B(_03765_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _16991_ (.A(_07786_),
    .B(_03765_),
    .Y(_02143_));
 sky130_fd_sc_hd__nor2_1 _16992_ (.A(_07800_),
    .B(_03765_),
    .Y(_02144_));
 sky130_fd_sc_hd__nor2_1 _16993_ (.A(_07809_),
    .B(_03765_),
    .Y(_02145_));
 sky130_fd_sc_hd__nor2_1 _16994_ (.A(_07818_),
    .B(_03765_),
    .Y(_02146_));
 sky130_fd_sc_hd__nor2_1 _16995_ (.A(_07831_),
    .B(_03765_),
    .Y(_02147_));
 sky130_fd_sc_hd__nor2_1 _16996_ (.A(_07843_),
    .B(_03765_),
    .Y(_02148_));
 sky130_fd_sc_hd__nor2_1 _16998_ (.A(_07850_),
    .B(_03765_),
    .Y(_02149_));
 sky130_fd_sc_hd__nor2_1 _16999_ (.A(_03491_),
    .B(_03765_),
    .Y(_02150_));
 sky130_fd_sc_hd__nor2_1 _17000_ (.A(_07581_),
    .B(_03765_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_1 _17001_ (.A(_07873_),
    .B(_03765_),
    .Y(_02152_));
 sky130_fd_sc_hd__nor2_1 _17002_ (.A(_07925_),
    .B(_03765_),
    .Y(_02153_));
 sky130_fd_sc_hd__nor2_1 _17003_ (.A(_07588_),
    .B(_03765_),
    .Y(_02154_));
 sky130_fd_sc_hd__nor2_1 _17004_ (.A(_07601_),
    .B(_03765_),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _17005_ (.A(_07610_),
    .B(_03765_),
    .Y(_02156_));
 sky130_fd_sc_hd__nor2_1 _17006_ (.A(_07620_),
    .B(_03765_),
    .Y(_02157_));
 sky130_fd_sc_hd__nor2_1 _17007_ (.A(_07628_),
    .B(_03765_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _17008_ (.A(_07635_),
    .B(_03765_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _17009_ (.A(_07646_),
    .B(_03765_),
    .Y(_02160_));
 sky130_fd_sc_hd__nand2_1 _17010_ (.A(_05436_),
    .B(_08304_),
    .Y(_03769_));
 sky130_fd_sc_hd__nor2_1 _17012_ (.A(_07930_),
    .B(_03769_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_1 _17013_ (.A(_08006_),
    .B(_03769_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _17014_ (.A(_08018_),
    .B(_03769_),
    .Y(_02163_));
 sky130_fd_sc_hd__nor2_1 _17015_ (.A(_08025_),
    .B(_03769_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _17016_ (.A(_08031_),
    .B(_03769_),
    .Y(_02165_));
 sky130_fd_sc_hd__nor2_1 _17017_ (.A(_08039_),
    .B(_03769_),
    .Y(_02166_));
 sky130_fd_sc_hd__nor2_1 _17018_ (.A(_08051_),
    .B(_03769_),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _17019_ (.A(_08064_),
    .B(_03769_),
    .Y(_02168_));
 sky130_fd_sc_hd__nor2_1 _17020_ (.A(_08071_),
    .B(_03769_),
    .Y(_02169_));
 sky130_fd_sc_hd__nor2_1 _17021_ (.A(_08082_),
    .B(_03769_),
    .Y(_02170_));
 sky130_fd_sc_hd__nor2_1 _17023_ (.A(_08091_),
    .B(_03769_),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_1 _17024_ (.A(_07934_),
    .B(_03769_),
    .Y(_02172_));
 sky130_fd_sc_hd__nor2_1 _17025_ (.A(_08102_),
    .B(_03769_),
    .Y(_02173_));
 sky130_fd_sc_hd__nor2_1 _17026_ (.A(_08114_),
    .B(_03769_),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_1 _17027_ (.A(_08125_),
    .B(_03769_),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _17028_ (.A(_08142_),
    .B(_03769_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _17029_ (.A(_08152_),
    .B(_03769_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _17030_ (.A(_08160_),
    .B(_03769_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _17031_ (.A(_08171_),
    .B(_03769_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_1 _17032_ (.A(_08184_),
    .B(_03769_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _17034_ (.A(_08204_),
    .B(_03769_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_1 _17035_ (.A(_08209_),
    .B(_03769_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_1 _17036_ (.A(_07937_),
    .B(_03769_),
    .Y(_02183_));
 sky130_fd_sc_hd__nor2_1 _17037_ (.A(_08221_),
    .B(_03769_),
    .Y(_02184_));
 sky130_fd_sc_hd__nor2_1 _17038_ (.A(_08254_),
    .B(_03769_),
    .Y(_02185_));
 sky130_fd_sc_hd__nor2_1 _17039_ (.A(_07942_),
    .B(_03769_),
    .Y(_02186_));
 sky130_fd_sc_hd__nor2_1 _17040_ (.A(_07949_),
    .B(_03769_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _17041_ (.A(_07956_),
    .B(_03769_),
    .Y(_02188_));
 sky130_fd_sc_hd__nor2_1 _17042_ (.A(_07965_),
    .B(_03769_),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _17043_ (.A(_07974_),
    .B(_03769_),
    .Y(_02190_));
 sky130_fd_sc_hd__nor2_1 _17044_ (.A(_07981_),
    .B(_03769_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _17045_ (.A(_07989_),
    .B(_03769_),
    .Y(_02192_));
 sky130_fd_sc_hd__nand2_1 _17046_ (.A(_05383_),
    .B(_08346_),
    .Y(_03773_));
 sky130_fd_sc_hd__nor2_1 _17048_ (.A(_07572_),
    .B(_03773_),
    .Y(_02193_));
 sky130_fd_sc_hd__nor2_1 _17049_ (.A(_07660_),
    .B(_03773_),
    .Y(_02194_));
 sky130_fd_sc_hd__nor2_1 _17050_ (.A(_07669_),
    .B(_03773_),
    .Y(_02195_));
 sky130_fd_sc_hd__nor2_1 _17051_ (.A(_07677_),
    .B(_03773_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _17052_ (.A(_07689_),
    .B(_03773_),
    .Y(_02197_));
 sky130_fd_sc_hd__nor2_1 _17053_ (.A(_07703_),
    .B(_03773_),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _17054_ (.A(_07709_),
    .B(_03773_),
    .Y(_02199_));
 sky130_fd_sc_hd__nor2_1 _17055_ (.A(_07715_),
    .B(_03773_),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_1 _17056_ (.A(_07731_),
    .B(_03773_),
    .Y(_02201_));
 sky130_fd_sc_hd__nor2_1 _17057_ (.A(_07745_),
    .B(_03773_),
    .Y(_02202_));
 sky130_fd_sc_hd__nor2_1 _17059_ (.A(_07752_),
    .B(_03773_),
    .Y(_02203_));
 sky130_fd_sc_hd__nor2_1 _17060_ (.A(_07577_),
    .B(_03773_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _17061_ (.A(_07766_),
    .B(_03773_),
    .Y(_02205_));
 sky130_fd_sc_hd__nor2_1 _17062_ (.A(_07777_),
    .B(_03773_),
    .Y(_02206_));
 sky130_fd_sc_hd__nor2_1 _17063_ (.A(_07786_),
    .B(_03773_),
    .Y(_02207_));
 sky130_fd_sc_hd__nor2_1 _17064_ (.A(_07800_),
    .B(_03773_),
    .Y(_02208_));
 sky130_fd_sc_hd__nor2_1 _17065_ (.A(_07809_),
    .B(_03773_),
    .Y(_02209_));
 sky130_fd_sc_hd__nor2_1 _17066_ (.A(_07818_),
    .B(_03773_),
    .Y(_02210_));
 sky130_fd_sc_hd__nor2_1 _17067_ (.A(_07831_),
    .B(_03773_),
    .Y(_02211_));
 sky130_fd_sc_hd__nor2_1 _17068_ (.A(_07843_),
    .B(_03773_),
    .Y(_02212_));
 sky130_fd_sc_hd__nor2_1 _17070_ (.A(_07850_),
    .B(_03773_),
    .Y(_02213_));
 sky130_fd_sc_hd__nor2_1 _17071_ (.A(_03491_),
    .B(_03773_),
    .Y(_02214_));
 sky130_fd_sc_hd__nor2_1 _17072_ (.A(_07581_),
    .B(_03773_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _17073_ (.A(_07873_),
    .B(_03773_),
    .Y(_02216_));
 sky130_fd_sc_hd__nor2_1 _17074_ (.A(_07925_),
    .B(_03773_),
    .Y(_02217_));
 sky130_fd_sc_hd__nor2_1 _17075_ (.A(_07588_),
    .B(_03773_),
    .Y(_02218_));
 sky130_fd_sc_hd__nor2_1 _17076_ (.A(_07601_),
    .B(_03773_),
    .Y(_02219_));
 sky130_fd_sc_hd__nor2_1 _17077_ (.A(_07610_),
    .B(_03773_),
    .Y(_02220_));
 sky130_fd_sc_hd__nor2_1 _17078_ (.A(_07620_),
    .B(_03773_),
    .Y(_02221_));
 sky130_fd_sc_hd__nor2_1 _17079_ (.A(_07628_),
    .B(_03773_),
    .Y(_02222_));
 sky130_fd_sc_hd__nor2_1 _17080_ (.A(_07635_),
    .B(_03773_),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _17081_ (.A(_07646_),
    .B(_03773_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_1 _17082_ (.A(_05436_),
    .B(_08390_),
    .Y(_03777_));
 sky130_fd_sc_hd__nor2_1 _17084_ (.A(_07930_),
    .B(_03777_),
    .Y(_02225_));
 sky130_fd_sc_hd__nor2_1 _17085_ (.A(_08006_),
    .B(_03777_),
    .Y(_02226_));
 sky130_fd_sc_hd__nor2_1 _17086_ (.A(_08018_),
    .B(_03777_),
    .Y(_02227_));
 sky130_fd_sc_hd__nor2_1 _17087_ (.A(_08025_),
    .B(_03777_),
    .Y(_02228_));
 sky130_fd_sc_hd__nor2_1 _17088_ (.A(_08031_),
    .B(_03777_),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _17089_ (.A(_08039_),
    .B(_03777_),
    .Y(_02230_));
 sky130_fd_sc_hd__nor2_1 _17090_ (.A(_08051_),
    .B(_03777_),
    .Y(_02231_));
 sky130_fd_sc_hd__nor2_1 _17091_ (.A(_08064_),
    .B(_03777_),
    .Y(_02232_));
 sky130_fd_sc_hd__nor2_1 _17092_ (.A(_08071_),
    .B(_03777_),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_1 _17093_ (.A(_08082_),
    .B(_03777_),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _17095_ (.A(_08091_),
    .B(_03777_),
    .Y(_02235_));
 sky130_fd_sc_hd__nor2_1 _17096_ (.A(_07934_),
    .B(_03777_),
    .Y(_02236_));
 sky130_fd_sc_hd__nor2_1 _17097_ (.A(_08102_),
    .B(_03777_),
    .Y(_02237_));
 sky130_fd_sc_hd__nor2_1 _17098_ (.A(_08114_),
    .B(_03777_),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_1 _17099_ (.A(_08125_),
    .B(_03777_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _17100_ (.A(_08142_),
    .B(_03777_),
    .Y(_02240_));
 sky130_fd_sc_hd__nor2_1 _17101_ (.A(_08152_),
    .B(_03777_),
    .Y(_02241_));
 sky130_fd_sc_hd__nor2_1 _17102_ (.A(_08160_),
    .B(_03777_),
    .Y(_02242_));
 sky130_fd_sc_hd__nor2_1 _17103_ (.A(_08171_),
    .B(_03777_),
    .Y(_02243_));
 sky130_fd_sc_hd__nor2_1 _17104_ (.A(_08184_),
    .B(_03777_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_1 _17106_ (.A(_08204_),
    .B(_03777_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _17107_ (.A(_08209_),
    .B(_03777_),
    .Y(_02246_));
 sky130_fd_sc_hd__nor2_1 _17108_ (.A(_07937_),
    .B(_03777_),
    .Y(_02247_));
 sky130_fd_sc_hd__nor2_1 _17109_ (.A(_08221_),
    .B(_03777_),
    .Y(_02248_));
 sky130_fd_sc_hd__nor2_1 _17110_ (.A(_08254_),
    .B(_03777_),
    .Y(_02249_));
 sky130_fd_sc_hd__nor2_1 _17111_ (.A(_07942_),
    .B(_03777_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _17112_ (.A(_07949_),
    .B(_03777_),
    .Y(_02251_));
 sky130_fd_sc_hd__nor2_1 _17113_ (.A(_07956_),
    .B(_03777_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor2_1 _17114_ (.A(_07965_),
    .B(_03777_),
    .Y(_02253_));
 sky130_fd_sc_hd__nor2_1 _17115_ (.A(_07974_),
    .B(_03777_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor2_1 _17116_ (.A(_07981_),
    .B(_03777_),
    .Y(_02255_));
 sky130_fd_sc_hd__nor2_1 _17117_ (.A(_07989_),
    .B(_03777_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand2_1 _17118_ (.A(_05383_),
    .B(_08431_),
    .Y(_03781_));
 sky130_fd_sc_hd__nor2_1 _17120_ (.A(_07572_),
    .B(_03781_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _17121_ (.A(_07660_),
    .B(_03781_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _17122_ (.A(_07669_),
    .B(_03781_),
    .Y(_02259_));
 sky130_fd_sc_hd__nor2_1 _17123_ (.A(_07677_),
    .B(_03781_),
    .Y(_02260_));
 sky130_fd_sc_hd__nor2_1 _17124_ (.A(_07689_),
    .B(_03781_),
    .Y(_02261_));
 sky130_fd_sc_hd__nor2_1 _17125_ (.A(_07703_),
    .B(_03781_),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_1 _17126_ (.A(_07709_),
    .B(_03781_),
    .Y(_02263_));
 sky130_fd_sc_hd__nor2_1 _17127_ (.A(_07715_),
    .B(_03781_),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _17128_ (.A(_07731_),
    .B(_03781_),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _17129_ (.A(_07745_),
    .B(_03781_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_1 _17131_ (.A(_07752_),
    .B(_03781_),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _17132_ (.A(_07577_),
    .B(_03781_),
    .Y(_02268_));
 sky130_fd_sc_hd__nor2_1 _17133_ (.A(_07766_),
    .B(_03781_),
    .Y(_02269_));
 sky130_fd_sc_hd__nor2_1 _17134_ (.A(_07777_),
    .B(_03781_),
    .Y(_02270_));
 sky130_fd_sc_hd__nor2_1 _17135_ (.A(_07786_),
    .B(_03781_),
    .Y(_02271_));
 sky130_fd_sc_hd__nor2_1 _17136_ (.A(_07800_),
    .B(_03781_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _17137_ (.A(_07809_),
    .B(_03781_),
    .Y(_02273_));
 sky130_fd_sc_hd__nor2_1 _17138_ (.A(_07818_),
    .B(_03781_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _17139_ (.A(_07831_),
    .B(_03781_),
    .Y(_02275_));
 sky130_fd_sc_hd__nor2_1 _17140_ (.A(_07843_),
    .B(_03781_),
    .Y(_02276_));
 sky130_fd_sc_hd__nor2_1 _17142_ (.A(_07850_),
    .B(_03781_),
    .Y(_02277_));
 sky130_fd_sc_hd__nor2_1 _17143_ (.A(_03491_),
    .B(_03781_),
    .Y(_02278_));
 sky130_fd_sc_hd__nor2_1 _17144_ (.A(_07581_),
    .B(_03781_),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_1 _17145_ (.A(_07873_),
    .B(_03781_),
    .Y(_02280_));
 sky130_fd_sc_hd__nor2_1 _17146_ (.A(_07925_),
    .B(_03781_),
    .Y(_02281_));
 sky130_fd_sc_hd__nor2_1 _17147_ (.A(_07588_),
    .B(_03781_),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2_1 _17148_ (.A(_07601_),
    .B(_03781_),
    .Y(_02283_));
 sky130_fd_sc_hd__nor2_1 _17149_ (.A(_07610_),
    .B(_03781_),
    .Y(_02284_));
 sky130_fd_sc_hd__nor2_1 _17150_ (.A(_07620_),
    .B(_03781_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _17151_ (.A(_07628_),
    .B(_03781_),
    .Y(_02286_));
 sky130_fd_sc_hd__nor2_1 _17152_ (.A(_07635_),
    .B(_03781_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_1 _17153_ (.A(_07646_),
    .B(_03781_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2b_1 _17154_ (.A_N(_05330_),
    .B(_05334_),
    .Y(_03785_));
 sky130_fd_sc_hd__nor2_1 _17156_ (.A(_07930_),
    .B(_03785_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _17157_ (.A(_08006_),
    .B(_03785_),
    .Y(_02290_));
 sky130_fd_sc_hd__nor2_1 _17158_ (.A(_08018_),
    .B(_03785_),
    .Y(_02291_));
 sky130_fd_sc_hd__nor2_1 _17159_ (.A(_08025_),
    .B(_03785_),
    .Y(_02292_));
 sky130_fd_sc_hd__nor2_1 _17160_ (.A(_08031_),
    .B(_03785_),
    .Y(_02293_));
 sky130_fd_sc_hd__nor2_1 _17161_ (.A(_08039_),
    .B(_03785_),
    .Y(_02294_));
 sky130_fd_sc_hd__nor2_1 _17162_ (.A(_08051_),
    .B(_03785_),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_1 _17163_ (.A(_08064_),
    .B(_03785_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor2_1 _17164_ (.A(_08071_),
    .B(_03785_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _17165_ (.A(_08082_),
    .B(_03785_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _17167_ (.A(_08091_),
    .B(_03785_),
    .Y(_02299_));
 sky130_fd_sc_hd__nor2_1 _17168_ (.A(_07934_),
    .B(_03785_),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _17169_ (.A(_08102_),
    .B(_03785_),
    .Y(_02301_));
 sky130_fd_sc_hd__nor2_1 _17170_ (.A(_08114_),
    .B(_03785_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _17171_ (.A(_08125_),
    .B(_03785_),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _17172_ (.A(_08142_),
    .B(_03785_),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _17173_ (.A(_08152_),
    .B(_03785_),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _17174_ (.A(_08160_),
    .B(_03785_),
    .Y(_02306_));
 sky130_fd_sc_hd__nor2_1 _17175_ (.A(_08171_),
    .B(_03785_),
    .Y(_02307_));
 sky130_fd_sc_hd__nor2_1 _17176_ (.A(_08184_),
    .B(_03785_),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2_1 _17178_ (.A(_08204_),
    .B(_03785_),
    .Y(_02309_));
 sky130_fd_sc_hd__nor2_1 _17179_ (.A(_08209_),
    .B(_03785_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor2_1 _17180_ (.A(_07937_),
    .B(_03785_),
    .Y(_02311_));
 sky130_fd_sc_hd__nor2_1 _17181_ (.A(_08221_),
    .B(_03785_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _17182_ (.A(_08254_),
    .B(_03785_),
    .Y(_02313_));
 sky130_fd_sc_hd__nor2_1 _17183_ (.A(_07942_),
    .B(_03785_),
    .Y(_02314_));
 sky130_fd_sc_hd__nor2_1 _17184_ (.A(_07949_),
    .B(_03785_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _17185_ (.A(_07956_),
    .B(_03785_),
    .Y(_02316_));
 sky130_fd_sc_hd__nor2_1 _17186_ (.A(_07965_),
    .B(_03785_),
    .Y(_02317_));
 sky130_fd_sc_hd__nor2_1 _17187_ (.A(_07974_),
    .B(_03785_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_1 _17188_ (.A(_07981_),
    .B(_03785_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _17189_ (.A(_07989_),
    .B(_03785_),
    .Y(_02320_));
 sky130_fd_sc_hd__inv_8 _17190_ (.A(ready),
    .Y(select));
 sky130_fd_sc_hd__mux4_2 _17195_ (.A0(\w[1][0] ),
    .A1(\w[3][0] ),
    .A2(\w[5][0] ),
    .A3(\w[7][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03793_));
 sky130_fd_sc_hd__mux4_2 _17199_ (.A0(\w[9][0] ),
    .A1(\w[11][0] ),
    .A2(\w[13][0] ),
    .A3(\w[15][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03797_));
 sky130_fd_sc_hd__mux4_2 _17203_ (.A0(\w[33][0] ),
    .A1(\w[35][0] ),
    .A2(\w[37][0] ),
    .A3(\w[39][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03801_));
 sky130_fd_sc_hd__mux4_2 _17206_ (.A0(\w[41][0] ),
    .A1(\w[43][0] ),
    .A2(\w[45][0] ),
    .A3(\w[47][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03804_));
 sky130_fd_sc_hd__mux4_2 _17210_ (.A0(_03793_),
    .A1(_03797_),
    .A2(_03801_),
    .A3(_03804_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03808_));
 sky130_fd_sc_hd__mux4_2 _17213_ (.A0(\w[17][0] ),
    .A1(\w[19][0] ),
    .A2(\w[21][0] ),
    .A3(\w[23][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03811_));
 sky130_fd_sc_hd__mux4_2 _17216_ (.A0(\w[25][0] ),
    .A1(\w[27][0] ),
    .A2(\w[29][0] ),
    .A3(\w[31][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03814_));
 sky130_fd_sc_hd__mux4_2 _17219_ (.A0(\w[49][0] ),
    .A1(\w[51][0] ),
    .A2(\w[53][0] ),
    .A3(\w[55][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03817_));
 sky130_fd_sc_hd__mux4_2 _17220_ (.A0(\w[57][0] ),
    .A1(\w[59][0] ),
    .A2(\w[61][0] ),
    .A3(\w[63][0] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03818_));
 sky130_fd_sc_hd__mux4_2 _17221_ (.A0(_03811_),
    .A1(_03814_),
    .A2(_03817_),
    .A3(_03818_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03819_));
 sky130_fd_sc_hd__mux2_2 _17222_ (.A0(_03808_),
    .A1(_03819_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[0] ));
 sky130_fd_sc_hd__mux4_2 _17223_ (.A0(\w[1][10] ),
    .A1(\w[3][10] ),
    .A2(\w[5][10] ),
    .A3(\w[7][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03820_));
 sky130_fd_sc_hd__mux4_2 _17224_ (.A0(\w[9][10] ),
    .A1(\w[11][10] ),
    .A2(\w[13][10] ),
    .A3(\w[15][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03821_));
 sky130_fd_sc_hd__mux4_2 _17225_ (.A0(\w[33][10] ),
    .A1(\w[35][10] ),
    .A2(\w[37][10] ),
    .A3(\w[39][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03822_));
 sky130_fd_sc_hd__mux4_2 _17226_ (.A0(\w[41][10] ),
    .A1(\w[43][10] ),
    .A2(\w[45][10] ),
    .A3(\w[47][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03823_));
 sky130_fd_sc_hd__mux4_2 _17227_ (.A0(_03820_),
    .A1(_03821_),
    .A2(_03822_),
    .A3(_03823_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03824_));
 sky130_fd_sc_hd__mux4_2 _17228_ (.A0(\w[17][10] ),
    .A1(\w[19][10] ),
    .A2(\w[21][10] ),
    .A3(\w[23][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03825_));
 sky130_fd_sc_hd__mux4_2 _17229_ (.A0(\w[25][10] ),
    .A1(\w[27][10] ),
    .A2(\w[29][10] ),
    .A3(\w[31][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03826_));
 sky130_fd_sc_hd__mux4_2 _17231_ (.A0(\w[49][10] ),
    .A1(\w[51][10] ),
    .A2(\w[53][10] ),
    .A3(\w[55][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03828_));
 sky130_fd_sc_hd__mux4_2 _17232_ (.A0(\w[57][10] ),
    .A1(\w[59][10] ),
    .A2(\w[61][10] ),
    .A3(\w[63][10] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03829_));
 sky130_fd_sc_hd__mux4_2 _17233_ (.A0(_03825_),
    .A1(_03826_),
    .A2(_03828_),
    .A3(_03829_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_2 _17234_ (.A0(_03824_),
    .A1(_03830_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[10] ));
 sky130_fd_sc_hd__mux4_2 _17236_ (.A0(\w[1][11] ),
    .A1(\w[3][11] ),
    .A2(\w[5][11] ),
    .A3(\w[7][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03832_));
 sky130_fd_sc_hd__mux4_2 _17237_ (.A0(\w[9][11] ),
    .A1(\w[11][11] ),
    .A2(\w[13][11] ),
    .A3(\w[15][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03833_));
 sky130_fd_sc_hd__mux4_2 _17238_ (.A0(\w[33][11] ),
    .A1(\w[35][11] ),
    .A2(\w[37][11] ),
    .A3(\w[39][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03834_));
 sky130_fd_sc_hd__mux4_2 _17239_ (.A0(\w[41][11] ),
    .A1(\w[43][11] ),
    .A2(\w[45][11] ),
    .A3(\w[47][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03835_));
 sky130_fd_sc_hd__mux4_2 _17240_ (.A0(_03832_),
    .A1(_03833_),
    .A2(_03834_),
    .A3(_03835_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03836_));
 sky130_fd_sc_hd__mux4_2 _17241_ (.A0(\w[17][11] ),
    .A1(\w[19][11] ),
    .A2(\w[21][11] ),
    .A3(\w[23][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03837_));
 sky130_fd_sc_hd__mux4_2 _17242_ (.A0(\w[25][11] ),
    .A1(\w[27][11] ),
    .A2(\w[29][11] ),
    .A3(\w[31][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03838_));
 sky130_fd_sc_hd__mux4_2 _17243_ (.A0(\w[49][11] ),
    .A1(\w[51][11] ),
    .A2(\w[53][11] ),
    .A3(\w[55][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03839_));
 sky130_fd_sc_hd__mux4_2 _17244_ (.A0(\w[57][11] ),
    .A1(\w[59][11] ),
    .A2(\w[61][11] ),
    .A3(\w[63][11] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03840_));
 sky130_fd_sc_hd__mux4_2 _17245_ (.A0(_03837_),
    .A1(_03838_),
    .A2(_03839_),
    .A3(_03840_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03841_));
 sky130_fd_sc_hd__mux2_2 _17246_ (.A0(_03836_),
    .A1(_03841_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[11] ));
 sky130_fd_sc_hd__mux4_2 _17248_ (.A0(\w[1][12] ),
    .A1(\w[3][12] ),
    .A2(\w[5][12] ),
    .A3(\w[7][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03843_));
 sky130_fd_sc_hd__mux4_2 _17249_ (.A0(\w[9][12] ),
    .A1(\w[11][12] ),
    .A2(\w[13][12] ),
    .A3(\w[15][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03844_));
 sky130_fd_sc_hd__mux4_2 _17250_ (.A0(\w[33][12] ),
    .A1(\w[35][12] ),
    .A2(\w[37][12] ),
    .A3(\w[39][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03845_));
 sky130_fd_sc_hd__mux4_2 _17251_ (.A0(\w[41][12] ),
    .A1(\w[43][12] ),
    .A2(\w[45][12] ),
    .A3(\w[47][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03846_));
 sky130_fd_sc_hd__mux4_2 _17252_ (.A0(_03843_),
    .A1(_03844_),
    .A2(_03845_),
    .A3(_03846_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03847_));
 sky130_fd_sc_hd__mux4_2 _17253_ (.A0(\w[17][12] ),
    .A1(\w[19][12] ),
    .A2(\w[21][12] ),
    .A3(\w[23][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03848_));
 sky130_fd_sc_hd__mux4_2 _17254_ (.A0(\w[25][12] ),
    .A1(\w[27][12] ),
    .A2(\w[29][12] ),
    .A3(\w[31][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03849_));
 sky130_fd_sc_hd__mux4_2 _17255_ (.A0(\w[49][12] ),
    .A1(\w[51][12] ),
    .A2(\w[53][12] ),
    .A3(\w[55][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03850_));
 sky130_fd_sc_hd__mux4_2 _17256_ (.A0(\w[57][12] ),
    .A1(\w[59][12] ),
    .A2(\w[61][12] ),
    .A3(\w[63][12] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03851_));
 sky130_fd_sc_hd__mux4_2 _17257_ (.A0(_03848_),
    .A1(_03849_),
    .A2(_03850_),
    .A3(_03851_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03852_));
 sky130_fd_sc_hd__mux2_2 _17258_ (.A0(_03847_),
    .A1(_03852_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[12] ));
 sky130_fd_sc_hd__mux4_2 _17259_ (.A0(\w[1][13] ),
    .A1(\w[3][13] ),
    .A2(\w[5][13] ),
    .A3(\w[7][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03853_));
 sky130_fd_sc_hd__mux4_2 _17261_ (.A0(\w[9][13] ),
    .A1(\w[11][13] ),
    .A2(\w[13][13] ),
    .A3(\w[15][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03855_));
 sky130_fd_sc_hd__mux4_2 _17262_ (.A0(\w[33][13] ),
    .A1(\w[35][13] ),
    .A2(\w[37][13] ),
    .A3(\w[39][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03856_));
 sky130_fd_sc_hd__mux4_2 _17263_ (.A0(\w[41][13] ),
    .A1(\w[43][13] ),
    .A2(\w[45][13] ),
    .A3(\w[47][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03857_));
 sky130_fd_sc_hd__mux4_2 _17264_ (.A0(_03853_),
    .A1(_03855_),
    .A2(_03856_),
    .A3(_03857_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03858_));
 sky130_fd_sc_hd__mux4_2 _17266_ (.A0(\w[17][13] ),
    .A1(\w[19][13] ),
    .A2(\w[21][13] ),
    .A3(\w[23][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03860_));
 sky130_fd_sc_hd__mux4_2 _17267_ (.A0(\w[25][13] ),
    .A1(\w[27][13] ),
    .A2(\w[29][13] ),
    .A3(\w[31][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03861_));
 sky130_fd_sc_hd__mux4_2 _17268_ (.A0(\w[49][13] ),
    .A1(\w[51][13] ),
    .A2(\w[53][13] ),
    .A3(\w[55][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03862_));
 sky130_fd_sc_hd__mux4_2 _17269_ (.A0(\w[57][13] ),
    .A1(\w[59][13] ),
    .A2(\w[61][13] ),
    .A3(\w[63][13] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03863_));
 sky130_fd_sc_hd__mux4_2 _17270_ (.A0(_03860_),
    .A1(_03861_),
    .A2(_03862_),
    .A3(_03863_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03864_));
 sky130_fd_sc_hd__mux2_2 _17271_ (.A0(_03858_),
    .A1(_03864_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[13] ));
 sky130_fd_sc_hd__mux4_2 _17272_ (.A0(\w[1][14] ),
    .A1(\w[3][14] ),
    .A2(\w[5][14] ),
    .A3(\w[7][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03865_));
 sky130_fd_sc_hd__mux4_2 _17274_ (.A0(\w[9][14] ),
    .A1(\w[11][14] ),
    .A2(\w[13][14] ),
    .A3(\w[15][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03867_));
 sky130_fd_sc_hd__mux4_2 _17275_ (.A0(\w[33][14] ),
    .A1(\w[35][14] ),
    .A2(\w[37][14] ),
    .A3(\w[39][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03868_));
 sky130_fd_sc_hd__mux4_2 _17276_ (.A0(\w[41][14] ),
    .A1(\w[43][14] ),
    .A2(\w[45][14] ),
    .A3(\w[47][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03869_));
 sky130_fd_sc_hd__mux4_2 _17278_ (.A0(_03865_),
    .A1(_03867_),
    .A2(_03868_),
    .A3(_03869_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03871_));
 sky130_fd_sc_hd__mux4_2 _17280_ (.A0(\w[17][14] ),
    .A1(\w[19][14] ),
    .A2(\w[21][14] ),
    .A3(\w[23][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03873_));
 sky130_fd_sc_hd__mux4_2 _17281_ (.A0(\w[25][14] ),
    .A1(\w[27][14] ),
    .A2(\w[29][14] ),
    .A3(\w[31][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03874_));
 sky130_fd_sc_hd__mux4_2 _17282_ (.A0(\w[49][14] ),
    .A1(\w[51][14] ),
    .A2(\w[53][14] ),
    .A3(\w[55][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03875_));
 sky130_fd_sc_hd__mux4_2 _17283_ (.A0(\w[57][14] ),
    .A1(\w[59][14] ),
    .A2(\w[61][14] ),
    .A3(\w[63][14] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03876_));
 sky130_fd_sc_hd__mux4_2 _17284_ (.A0(_03873_),
    .A1(_03874_),
    .A2(_03875_),
    .A3(_03876_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03877_));
 sky130_fd_sc_hd__mux2_2 _17285_ (.A0(_03871_),
    .A1(_03877_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[14] ));
 sky130_fd_sc_hd__mux4_2 _17286_ (.A0(\w[1][15] ),
    .A1(\w[3][15] ),
    .A2(\w[5][15] ),
    .A3(\w[7][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03878_));
 sky130_fd_sc_hd__mux4_2 _17287_ (.A0(\w[9][15] ),
    .A1(\w[11][15] ),
    .A2(\w[13][15] ),
    .A3(\w[15][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03879_));
 sky130_fd_sc_hd__mux4_2 _17288_ (.A0(\w[33][15] ),
    .A1(\w[35][15] ),
    .A2(\w[37][15] ),
    .A3(\w[39][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03880_));
 sky130_fd_sc_hd__mux4_2 _17290_ (.A0(\w[41][15] ),
    .A1(\w[43][15] ),
    .A2(\w[45][15] ),
    .A3(\w[47][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03882_));
 sky130_fd_sc_hd__mux4_2 _17291_ (.A0(_03878_),
    .A1(_03879_),
    .A2(_03880_),
    .A3(_03882_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03883_));
 sky130_fd_sc_hd__mux4_2 _17292_ (.A0(\w[17][15] ),
    .A1(\w[19][15] ),
    .A2(\w[21][15] ),
    .A3(\w[23][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03884_));
 sky130_fd_sc_hd__mux4_2 _17294_ (.A0(\w[25][15] ),
    .A1(\w[27][15] ),
    .A2(\w[29][15] ),
    .A3(\w[31][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03886_));
 sky130_fd_sc_hd__mux4_2 _17295_ (.A0(\w[49][15] ),
    .A1(\w[51][15] ),
    .A2(\w[53][15] ),
    .A3(\w[55][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03887_));
 sky130_fd_sc_hd__mux4_2 _17296_ (.A0(\w[57][15] ),
    .A1(\w[59][15] ),
    .A2(\w[61][15] ),
    .A3(\w[63][15] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03888_));
 sky130_fd_sc_hd__mux4_2 _17297_ (.A0(_03884_),
    .A1(_03886_),
    .A2(_03887_),
    .A3(_03888_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_2 _17298_ (.A0(_03883_),
    .A1(_03889_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[15] ));
 sky130_fd_sc_hd__mux4_2 _17299_ (.A0(\w[1][16] ),
    .A1(\w[3][16] ),
    .A2(\w[5][16] ),
    .A3(\w[7][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03890_));
 sky130_fd_sc_hd__mux4_2 _17300_ (.A0(\w[9][16] ),
    .A1(\w[11][16] ),
    .A2(\w[13][16] ),
    .A3(\w[15][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03891_));
 sky130_fd_sc_hd__mux4_2 _17301_ (.A0(\w[33][16] ),
    .A1(\w[35][16] ),
    .A2(\w[37][16] ),
    .A3(\w[39][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03892_));
 sky130_fd_sc_hd__mux4_2 _17303_ (.A0(\w[41][16] ),
    .A1(\w[43][16] ),
    .A2(\w[45][16] ),
    .A3(\w[47][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03894_));
 sky130_fd_sc_hd__mux4_2 _17305_ (.A0(_03890_),
    .A1(_03891_),
    .A2(_03892_),
    .A3(_03894_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03896_));
 sky130_fd_sc_hd__mux4_2 _17306_ (.A0(\w[17][16] ),
    .A1(\w[19][16] ),
    .A2(\w[21][16] ),
    .A3(\w[23][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03897_));
 sky130_fd_sc_hd__mux4_2 _17308_ (.A0(\w[25][16] ),
    .A1(\w[27][16] ),
    .A2(\w[29][16] ),
    .A3(\w[31][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03899_));
 sky130_fd_sc_hd__mux4_2 _17309_ (.A0(\w[49][16] ),
    .A1(\w[51][16] ),
    .A2(\w[53][16] ),
    .A3(\w[55][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03900_));
 sky130_fd_sc_hd__mux4_2 _17310_ (.A0(\w[57][16] ),
    .A1(\w[59][16] ),
    .A2(\w[61][16] ),
    .A3(\w[63][16] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03901_));
 sky130_fd_sc_hd__mux4_2 _17312_ (.A0(_03897_),
    .A1(_03899_),
    .A2(_03900_),
    .A3(_03901_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03903_));
 sky130_fd_sc_hd__mux2_2 _17313_ (.A0(_03896_),
    .A1(_03903_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[16] ));
 sky130_fd_sc_hd__mux4_2 _17314_ (.A0(\w[1][17] ),
    .A1(\w[3][17] ),
    .A2(\w[5][17] ),
    .A3(\w[7][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03904_));
 sky130_fd_sc_hd__mux4_2 _17315_ (.A0(\w[9][17] ),
    .A1(\w[11][17] ),
    .A2(\w[13][17] ),
    .A3(\w[15][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03905_));
 sky130_fd_sc_hd__mux4_2 _17317_ (.A0(\w[33][17] ),
    .A1(\w[35][17] ),
    .A2(\w[37][17] ),
    .A3(\w[39][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03907_));
 sky130_fd_sc_hd__mux4_2 _17318_ (.A0(\w[41][17] ),
    .A1(\w[43][17] ),
    .A2(\w[45][17] ),
    .A3(\w[47][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03908_));
 sky130_fd_sc_hd__mux4_2 _17319_ (.A0(_03904_),
    .A1(_03905_),
    .A2(_03907_),
    .A3(_03908_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03909_));
 sky130_fd_sc_hd__mux4_2 _17320_ (.A0(\w[17][17] ),
    .A1(\w[19][17] ),
    .A2(\w[21][17] ),
    .A3(\w[23][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03910_));
 sky130_fd_sc_hd__mux4_2 _17321_ (.A0(\w[25][17] ),
    .A1(\w[27][17] ),
    .A2(\w[29][17] ),
    .A3(\w[31][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03911_));
 sky130_fd_sc_hd__mux4_2 _17322_ (.A0(\w[49][17] ),
    .A1(\w[51][17] ),
    .A2(\w[53][17] ),
    .A3(\w[55][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03912_));
 sky130_fd_sc_hd__mux4_2 _17324_ (.A0(\w[57][17] ),
    .A1(\w[59][17] ),
    .A2(\w[61][17] ),
    .A3(\w[63][17] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03914_));
 sky130_fd_sc_hd__mux4_2 _17325_ (.A0(_03910_),
    .A1(_03911_),
    .A2(_03912_),
    .A3(_03914_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_2 _17326_ (.A0(_03909_),
    .A1(_03915_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[17] ));
 sky130_fd_sc_hd__mux4_2 _17327_ (.A0(\w[1][18] ),
    .A1(\w[3][18] ),
    .A2(\w[5][18] ),
    .A3(\w[7][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03916_));
 sky130_fd_sc_hd__mux4_2 _17328_ (.A0(\w[9][18] ),
    .A1(\w[11][18] ),
    .A2(\w[13][18] ),
    .A3(\w[15][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03917_));
 sky130_fd_sc_hd__mux4_2 _17330_ (.A0(\w[33][18] ),
    .A1(\w[35][18] ),
    .A2(\w[37][18] ),
    .A3(\w[39][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03919_));
 sky130_fd_sc_hd__mux4_2 _17331_ (.A0(\w[41][18] ),
    .A1(\w[43][18] ),
    .A2(\w[45][18] ),
    .A3(\w[47][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03920_));
 sky130_fd_sc_hd__mux4_2 _17332_ (.A0(_03916_),
    .A1(_03917_),
    .A2(_03919_),
    .A3(_03920_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03921_));
 sky130_fd_sc_hd__mux4_2 _17333_ (.A0(\w[17][18] ),
    .A1(\w[19][18] ),
    .A2(\w[21][18] ),
    .A3(\w[23][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03922_));
 sky130_fd_sc_hd__mux4_2 _17334_ (.A0(\w[25][18] ),
    .A1(\w[27][18] ),
    .A2(\w[29][18] ),
    .A3(\w[31][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03923_));
 sky130_fd_sc_hd__mux4_2 _17335_ (.A0(\w[49][18] ),
    .A1(\w[51][18] ),
    .A2(\w[53][18] ),
    .A3(\w[55][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03924_));
 sky130_fd_sc_hd__mux4_2 _17337_ (.A0(\w[57][18] ),
    .A1(\w[59][18] ),
    .A2(\w[61][18] ),
    .A3(\w[63][18] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03926_));
 sky130_fd_sc_hd__mux4_2 _17339_ (.A0(_03922_),
    .A1(_03923_),
    .A2(_03924_),
    .A3(_03926_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03928_));
 sky130_fd_sc_hd__mux2_2 _17341_ (.A0(_03921_),
    .A1(_03928_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[18] ));
 sky130_fd_sc_hd__mux4_2 _17342_ (.A0(\w[1][19] ),
    .A1(\w[3][19] ),
    .A2(\w[5][19] ),
    .A3(\w[7][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03930_));
 sky130_fd_sc_hd__mux4_2 _17343_ (.A0(\w[9][19] ),
    .A1(\w[11][19] ),
    .A2(\w[13][19] ),
    .A3(\w[15][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03931_));
 sky130_fd_sc_hd__mux4_2 _17344_ (.A0(\w[33][19] ),
    .A1(\w[35][19] ),
    .A2(\w[37][19] ),
    .A3(\w[39][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03932_));
 sky130_fd_sc_hd__mux4_2 _17345_ (.A0(\w[41][19] ),
    .A1(\w[43][19] ),
    .A2(\w[45][19] ),
    .A3(\w[47][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03933_));
 sky130_fd_sc_hd__mux4_2 _17346_ (.A0(_03930_),
    .A1(_03931_),
    .A2(_03932_),
    .A3(_03933_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03934_));
 sky130_fd_sc_hd__mux4_2 _17347_ (.A0(\w[17][19] ),
    .A1(\w[19][19] ),
    .A2(\w[21][19] ),
    .A3(\w[23][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03935_));
 sky130_fd_sc_hd__mux4_2 _17348_ (.A0(\w[25][19] ),
    .A1(\w[27][19] ),
    .A2(\w[29][19] ),
    .A3(\w[31][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03936_));
 sky130_fd_sc_hd__mux4_2 _17350_ (.A0(\w[49][19] ),
    .A1(\w[51][19] ),
    .A2(\w[53][19] ),
    .A3(\w[55][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03938_));
 sky130_fd_sc_hd__mux4_2 _17351_ (.A0(\w[57][19] ),
    .A1(\w[59][19] ),
    .A2(\w[61][19] ),
    .A3(\w[63][19] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03939_));
 sky130_fd_sc_hd__mux4_2 _17352_ (.A0(_03935_),
    .A1(_03936_),
    .A2(_03938_),
    .A3(_03939_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03940_));
 sky130_fd_sc_hd__mux2_2 _17353_ (.A0(_03934_),
    .A1(_03940_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[19] ));
 sky130_fd_sc_hd__mux4_2 _17354_ (.A0(\w[1][1] ),
    .A1(\w[3][1] ),
    .A2(\w[5][1] ),
    .A3(\w[7][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03941_));
 sky130_fd_sc_hd__mux4_2 _17355_ (.A0(\w[9][1] ),
    .A1(\w[11][1] ),
    .A2(\w[13][1] ),
    .A3(\w[15][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03942_));
 sky130_fd_sc_hd__mux4_2 _17356_ (.A0(\w[33][1] ),
    .A1(\w[35][1] ),
    .A2(\w[37][1] ),
    .A3(\w[39][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03943_));
 sky130_fd_sc_hd__mux4_2 _17357_ (.A0(\w[41][1] ),
    .A1(\w[43][1] ),
    .A2(\w[45][1] ),
    .A3(\w[47][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03944_));
 sky130_fd_sc_hd__mux4_2 _17358_ (.A0(_03941_),
    .A1(_03942_),
    .A2(_03943_),
    .A3(_03944_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03945_));
 sky130_fd_sc_hd__mux4_2 _17359_ (.A0(\w[17][1] ),
    .A1(\w[19][1] ),
    .A2(\w[21][1] ),
    .A3(\w[23][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03946_));
 sky130_fd_sc_hd__mux4_2 _17360_ (.A0(\w[25][1] ),
    .A1(\w[27][1] ),
    .A2(\w[29][1] ),
    .A3(\w[31][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03947_));
 sky130_fd_sc_hd__mux4_2 _17362_ (.A0(\w[49][1] ),
    .A1(\w[51][1] ),
    .A2(\w[53][1] ),
    .A3(\w[55][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03949_));
 sky130_fd_sc_hd__mux4_2 _17363_ (.A0(\w[57][1] ),
    .A1(\w[59][1] ),
    .A2(\w[61][1] ),
    .A3(\w[63][1] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03950_));
 sky130_fd_sc_hd__mux4_2 _17364_ (.A0(_03946_),
    .A1(_03947_),
    .A2(_03949_),
    .A3(_03950_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03951_));
 sky130_fd_sc_hd__mux2_2 _17365_ (.A0(_03945_),
    .A1(_03951_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[1] ));
 sky130_fd_sc_hd__mux4_2 _17367_ (.A0(\w[1][20] ),
    .A1(\w[3][20] ),
    .A2(\w[5][20] ),
    .A3(\w[7][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03953_));
 sky130_fd_sc_hd__mux4_2 _17368_ (.A0(\w[9][20] ),
    .A1(\w[11][20] ),
    .A2(\w[13][20] ),
    .A3(\w[15][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03954_));
 sky130_fd_sc_hd__mux4_2 _17369_ (.A0(\w[33][20] ),
    .A1(\w[35][20] ),
    .A2(\w[37][20] ),
    .A3(\w[39][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03955_));
 sky130_fd_sc_hd__mux4_2 _17370_ (.A0(\w[41][20] ),
    .A1(\w[43][20] ),
    .A2(\w[45][20] ),
    .A3(\w[47][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03956_));
 sky130_fd_sc_hd__mux4_2 _17371_ (.A0(_03953_),
    .A1(_03954_),
    .A2(_03955_),
    .A3(_03956_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03957_));
 sky130_fd_sc_hd__mux4_2 _17372_ (.A0(\w[17][20] ),
    .A1(\w[19][20] ),
    .A2(\w[21][20] ),
    .A3(\w[23][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03958_));
 sky130_fd_sc_hd__mux4_2 _17373_ (.A0(\w[25][20] ),
    .A1(\w[27][20] ),
    .A2(\w[29][20] ),
    .A3(\w[31][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03959_));
 sky130_fd_sc_hd__mux4_2 _17374_ (.A0(\w[49][20] ),
    .A1(\w[51][20] ),
    .A2(\w[53][20] ),
    .A3(\w[55][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03960_));
 sky130_fd_sc_hd__mux4_2 _17375_ (.A0(\w[57][20] ),
    .A1(\w[59][20] ),
    .A2(\w[61][20] ),
    .A3(\w[63][20] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03961_));
 sky130_fd_sc_hd__mux4_2 _17376_ (.A0(_03958_),
    .A1(_03959_),
    .A2(_03960_),
    .A3(_03961_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03962_));
 sky130_fd_sc_hd__mux2_2 _17377_ (.A0(_03957_),
    .A1(_03962_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[20] ));
 sky130_fd_sc_hd__mux4_2 _17379_ (.A0(\w[1][21] ),
    .A1(\w[3][21] ),
    .A2(\w[5][21] ),
    .A3(\w[7][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03964_));
 sky130_fd_sc_hd__mux4_2 _17380_ (.A0(\w[9][21] ),
    .A1(\w[11][21] ),
    .A2(\w[13][21] ),
    .A3(\w[15][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03965_));
 sky130_fd_sc_hd__mux4_2 _17381_ (.A0(\w[33][21] ),
    .A1(\w[35][21] ),
    .A2(\w[37][21] ),
    .A3(\w[39][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03966_));
 sky130_fd_sc_hd__mux4_2 _17382_ (.A0(\w[41][21] ),
    .A1(\w[43][21] ),
    .A2(\w[45][21] ),
    .A3(\w[47][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03967_));
 sky130_fd_sc_hd__mux4_2 _17383_ (.A0(_03964_),
    .A1(_03965_),
    .A2(_03966_),
    .A3(_03967_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03968_));
 sky130_fd_sc_hd__mux4_2 _17384_ (.A0(\w[17][21] ),
    .A1(\w[19][21] ),
    .A2(\w[21][21] ),
    .A3(\w[23][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03969_));
 sky130_fd_sc_hd__mux4_2 _17385_ (.A0(\w[25][21] ),
    .A1(\w[27][21] ),
    .A2(\w[29][21] ),
    .A3(\w[31][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03970_));
 sky130_fd_sc_hd__mux4_2 _17386_ (.A0(\w[49][21] ),
    .A1(\w[51][21] ),
    .A2(\w[53][21] ),
    .A3(\w[55][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03971_));
 sky130_fd_sc_hd__mux4_2 _17387_ (.A0(\w[57][21] ),
    .A1(\w[59][21] ),
    .A2(\w[61][21] ),
    .A3(\w[63][21] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03972_));
 sky130_fd_sc_hd__mux4_2 _17388_ (.A0(_03969_),
    .A1(_03970_),
    .A2(_03971_),
    .A3(_03972_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03973_));
 sky130_fd_sc_hd__mux2_2 _17389_ (.A0(_03968_),
    .A1(_03973_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[21] ));
 sky130_fd_sc_hd__mux4_2 _17390_ (.A0(\w[1][22] ),
    .A1(\w[3][22] ),
    .A2(\w[5][22] ),
    .A3(\w[7][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03974_));
 sky130_fd_sc_hd__mux4_2 _17392_ (.A0(\w[9][22] ),
    .A1(\w[11][22] ),
    .A2(\w[13][22] ),
    .A3(\w[15][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03976_));
 sky130_fd_sc_hd__mux4_2 _17393_ (.A0(\w[33][22] ),
    .A1(\w[35][22] ),
    .A2(\w[37][22] ),
    .A3(\w[39][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03977_));
 sky130_fd_sc_hd__mux4_2 _17394_ (.A0(\w[41][22] ),
    .A1(\w[43][22] ),
    .A2(\w[45][22] ),
    .A3(\w[47][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03978_));
 sky130_fd_sc_hd__mux4_2 _17395_ (.A0(_03974_),
    .A1(_03976_),
    .A2(_03977_),
    .A3(_03978_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03979_));
 sky130_fd_sc_hd__mux4_2 _17397_ (.A0(\w[17][22] ),
    .A1(\w[19][22] ),
    .A2(\w[21][22] ),
    .A3(\w[23][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03981_));
 sky130_fd_sc_hd__mux4_2 _17398_ (.A0(\w[25][22] ),
    .A1(\w[27][22] ),
    .A2(\w[29][22] ),
    .A3(\w[31][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03982_));
 sky130_fd_sc_hd__mux4_2 _17399_ (.A0(\w[49][22] ),
    .A1(\w[51][22] ),
    .A2(\w[53][22] ),
    .A3(\w[55][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03983_));
 sky130_fd_sc_hd__mux4_2 _17400_ (.A0(\w[57][22] ),
    .A1(\w[59][22] ),
    .A2(\w[61][22] ),
    .A3(\w[63][22] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03984_));
 sky130_fd_sc_hd__mux4_2 _17401_ (.A0(_03981_),
    .A1(_03982_),
    .A2(_03983_),
    .A3(_03984_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03985_));
 sky130_fd_sc_hd__mux2_2 _17402_ (.A0(_03979_),
    .A1(_03985_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[22] ));
 sky130_fd_sc_hd__mux4_2 _17403_ (.A0(\w[1][23] ),
    .A1(\w[3][23] ),
    .A2(\w[5][23] ),
    .A3(\w[7][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03986_));
 sky130_fd_sc_hd__mux4_2 _17405_ (.A0(\w[9][23] ),
    .A1(\w[11][23] ),
    .A2(\w[13][23] ),
    .A3(\w[15][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03988_));
 sky130_fd_sc_hd__mux4_2 _17406_ (.A0(\w[33][23] ),
    .A1(\w[35][23] ),
    .A2(\w[37][23] ),
    .A3(\w[39][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03989_));
 sky130_fd_sc_hd__mux4_2 _17407_ (.A0(\w[41][23] ),
    .A1(\w[43][23] ),
    .A2(\w[45][23] ),
    .A3(\w[47][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03990_));
 sky130_fd_sc_hd__mux4_2 _17409_ (.A0(_03986_),
    .A1(_03988_),
    .A2(_03989_),
    .A3(_03990_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03992_));
 sky130_fd_sc_hd__mux4_2 _17411_ (.A0(\w[17][23] ),
    .A1(\w[19][23] ),
    .A2(\w[21][23] ),
    .A3(\w[23][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03994_));
 sky130_fd_sc_hd__mux4_2 _17412_ (.A0(\w[25][23] ),
    .A1(\w[27][23] ),
    .A2(\w[29][23] ),
    .A3(\w[31][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03995_));
 sky130_fd_sc_hd__mux4_2 _17413_ (.A0(\w[49][23] ),
    .A1(\w[51][23] ),
    .A2(\w[53][23] ),
    .A3(\w[55][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03996_));
 sky130_fd_sc_hd__mux4_2 _17414_ (.A0(\w[57][23] ),
    .A1(\w[59][23] ),
    .A2(\w[61][23] ),
    .A3(\w[63][23] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03997_));
 sky130_fd_sc_hd__mux4_2 _17415_ (.A0(_03994_),
    .A1(_03995_),
    .A2(_03996_),
    .A3(_03997_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_03998_));
 sky130_fd_sc_hd__mux2_2 _17416_ (.A0(_03992_),
    .A1(_03998_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[23] ));
 sky130_fd_sc_hd__mux4_2 _17417_ (.A0(\w[1][24] ),
    .A1(\w[3][24] ),
    .A2(\w[5][24] ),
    .A3(\w[7][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_03999_));
 sky130_fd_sc_hd__mux4_2 _17418_ (.A0(\w[9][24] ),
    .A1(\w[11][24] ),
    .A2(\w[13][24] ),
    .A3(\w[15][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04000_));
 sky130_fd_sc_hd__mux4_2 _17419_ (.A0(\w[33][24] ),
    .A1(\w[35][24] ),
    .A2(\w[37][24] ),
    .A3(\w[39][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04001_));
 sky130_fd_sc_hd__mux4_2 _17421_ (.A0(\w[41][24] ),
    .A1(\w[43][24] ),
    .A2(\w[45][24] ),
    .A3(\w[47][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04003_));
 sky130_fd_sc_hd__mux4_2 _17422_ (.A0(_03999_),
    .A1(_04000_),
    .A2(_04001_),
    .A3(_04003_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04004_));
 sky130_fd_sc_hd__mux4_2 _17423_ (.A0(\w[17][24] ),
    .A1(\w[19][24] ),
    .A2(\w[21][24] ),
    .A3(\w[23][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04005_));
 sky130_fd_sc_hd__mux4_2 _17425_ (.A0(\w[25][24] ),
    .A1(\w[27][24] ),
    .A2(\w[29][24] ),
    .A3(\w[31][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04007_));
 sky130_fd_sc_hd__mux4_2 _17426_ (.A0(\w[49][24] ),
    .A1(\w[51][24] ),
    .A2(\w[53][24] ),
    .A3(\w[55][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04008_));
 sky130_fd_sc_hd__mux4_2 _17427_ (.A0(\w[57][24] ),
    .A1(\w[59][24] ),
    .A2(\w[61][24] ),
    .A3(\w[63][24] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04009_));
 sky130_fd_sc_hd__mux4_2 _17428_ (.A0(_04005_),
    .A1(_04007_),
    .A2(_04008_),
    .A3(_04009_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04010_));
 sky130_fd_sc_hd__mux2_2 _17429_ (.A0(_04004_),
    .A1(_04010_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[24] ));
 sky130_fd_sc_hd__mux4_2 _17430_ (.A0(\w[1][25] ),
    .A1(\w[3][25] ),
    .A2(\w[5][25] ),
    .A3(\w[7][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04011_));
 sky130_fd_sc_hd__mux4_2 _17431_ (.A0(\w[9][25] ),
    .A1(\w[11][25] ),
    .A2(\w[13][25] ),
    .A3(\w[15][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04012_));
 sky130_fd_sc_hd__mux4_2 _17432_ (.A0(\w[33][25] ),
    .A1(\w[35][25] ),
    .A2(\w[37][25] ),
    .A3(\w[39][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04013_));
 sky130_fd_sc_hd__mux4_2 _17434_ (.A0(\w[41][25] ),
    .A1(\w[43][25] ),
    .A2(\w[45][25] ),
    .A3(\w[47][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04015_));
 sky130_fd_sc_hd__mux4_2 _17436_ (.A0(_04011_),
    .A1(_04012_),
    .A2(_04013_),
    .A3(_04015_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04017_));
 sky130_fd_sc_hd__mux4_2 _17437_ (.A0(\w[17][25] ),
    .A1(\w[19][25] ),
    .A2(\w[21][25] ),
    .A3(\w[23][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04018_));
 sky130_fd_sc_hd__mux4_2 _17439_ (.A0(\w[25][25] ),
    .A1(\w[27][25] ),
    .A2(\w[29][25] ),
    .A3(\w[31][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04020_));
 sky130_fd_sc_hd__mux4_2 _17440_ (.A0(\w[49][25] ),
    .A1(\w[51][25] ),
    .A2(\w[53][25] ),
    .A3(\w[55][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04021_));
 sky130_fd_sc_hd__mux4_2 _17441_ (.A0(\w[57][25] ),
    .A1(\w[59][25] ),
    .A2(\w[61][25] ),
    .A3(\w[63][25] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04022_));
 sky130_fd_sc_hd__mux4_2 _17443_ (.A0(_04018_),
    .A1(_04020_),
    .A2(_04021_),
    .A3(_04022_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04024_));
 sky130_fd_sc_hd__mux2_2 _17444_ (.A0(_04017_),
    .A1(_04024_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[25] ));
 sky130_fd_sc_hd__mux4_2 _17445_ (.A0(\w[1][26] ),
    .A1(\w[3][26] ),
    .A2(\w[5][26] ),
    .A3(\w[7][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04025_));
 sky130_fd_sc_hd__mux4_2 _17446_ (.A0(\w[9][26] ),
    .A1(\w[11][26] ),
    .A2(\w[13][26] ),
    .A3(\w[15][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04026_));
 sky130_fd_sc_hd__mux4_2 _17448_ (.A0(\w[33][26] ),
    .A1(\w[35][26] ),
    .A2(\w[37][26] ),
    .A3(\w[39][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04028_));
 sky130_fd_sc_hd__mux4_2 _17449_ (.A0(\w[41][26] ),
    .A1(\w[43][26] ),
    .A2(\w[45][26] ),
    .A3(\w[47][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04029_));
 sky130_fd_sc_hd__mux4_2 _17450_ (.A0(_04025_),
    .A1(_04026_),
    .A2(_04028_),
    .A3(_04029_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04030_));
 sky130_fd_sc_hd__mux4_2 _17451_ (.A0(\w[17][26] ),
    .A1(\w[19][26] ),
    .A2(\w[21][26] ),
    .A3(\w[23][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04031_));
 sky130_fd_sc_hd__mux4_2 _17452_ (.A0(\w[25][26] ),
    .A1(\w[27][26] ),
    .A2(\w[29][26] ),
    .A3(\w[31][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04032_));
 sky130_fd_sc_hd__mux4_2 _17453_ (.A0(\w[49][26] ),
    .A1(\w[51][26] ),
    .A2(\w[53][26] ),
    .A3(\w[55][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04033_));
 sky130_fd_sc_hd__mux4_2 _17455_ (.A0(\w[57][26] ),
    .A1(\w[59][26] ),
    .A2(\w[61][26] ),
    .A3(\w[63][26] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04035_));
 sky130_fd_sc_hd__mux4_2 _17456_ (.A0(_04031_),
    .A1(_04032_),
    .A2(_04033_),
    .A3(_04035_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04036_));
 sky130_fd_sc_hd__mux2_2 _17457_ (.A0(_04030_),
    .A1(_04036_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[26] ));
 sky130_fd_sc_hd__mux4_2 _17458_ (.A0(\w[1][27] ),
    .A1(\w[3][27] ),
    .A2(\w[5][27] ),
    .A3(\w[7][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04037_));
 sky130_fd_sc_hd__mux4_2 _17459_ (.A0(\w[9][27] ),
    .A1(\w[11][27] ),
    .A2(\w[13][27] ),
    .A3(\w[15][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04038_));
 sky130_fd_sc_hd__mux4_2 _17461_ (.A0(\w[33][27] ),
    .A1(\w[35][27] ),
    .A2(\w[37][27] ),
    .A3(\w[39][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04040_));
 sky130_fd_sc_hd__mux4_2 _17462_ (.A0(\w[41][27] ),
    .A1(\w[43][27] ),
    .A2(\w[45][27] ),
    .A3(\w[47][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04041_));
 sky130_fd_sc_hd__mux4_2 _17463_ (.A0(_04037_),
    .A1(_04038_),
    .A2(_04040_),
    .A3(_04041_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04042_));
 sky130_fd_sc_hd__mux4_2 _17464_ (.A0(\w[17][27] ),
    .A1(\w[19][27] ),
    .A2(\w[21][27] ),
    .A3(\w[23][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04043_));
 sky130_fd_sc_hd__mux4_2 _17465_ (.A0(\w[25][27] ),
    .A1(\w[27][27] ),
    .A2(\w[29][27] ),
    .A3(\w[31][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04044_));
 sky130_fd_sc_hd__mux4_2 _17466_ (.A0(\w[49][27] ),
    .A1(\w[51][27] ),
    .A2(\w[53][27] ),
    .A3(\w[55][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04045_));
 sky130_fd_sc_hd__mux4_2 _17468_ (.A0(\w[57][27] ),
    .A1(\w[59][27] ),
    .A2(\w[61][27] ),
    .A3(\w[63][27] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04047_));
 sky130_fd_sc_hd__mux4_2 _17470_ (.A0(_04043_),
    .A1(_04044_),
    .A2(_04045_),
    .A3(_04047_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04049_));
 sky130_fd_sc_hd__mux2_2 _17472_ (.A0(_04042_),
    .A1(_04049_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[27] ));
 sky130_fd_sc_hd__mux4_2 _17473_ (.A0(\w[1][28] ),
    .A1(\w[3][28] ),
    .A2(\w[5][28] ),
    .A3(\w[7][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04051_));
 sky130_fd_sc_hd__mux4_2 _17474_ (.A0(\w[9][28] ),
    .A1(\w[11][28] ),
    .A2(\w[13][28] ),
    .A3(\w[15][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04052_));
 sky130_fd_sc_hd__mux4_2 _17475_ (.A0(\w[33][28] ),
    .A1(\w[35][28] ),
    .A2(\w[37][28] ),
    .A3(\w[39][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04053_));
 sky130_fd_sc_hd__mux4_2 _17476_ (.A0(\w[41][28] ),
    .A1(\w[43][28] ),
    .A2(\w[45][28] ),
    .A3(\w[47][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04054_));
 sky130_fd_sc_hd__mux4_2 _17477_ (.A0(_04051_),
    .A1(_04052_),
    .A2(_04053_),
    .A3(_04054_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04055_));
 sky130_fd_sc_hd__mux4_2 _17478_ (.A0(\w[17][28] ),
    .A1(\w[19][28] ),
    .A2(\w[21][28] ),
    .A3(\w[23][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04056_));
 sky130_fd_sc_hd__mux4_2 _17479_ (.A0(\w[25][28] ),
    .A1(\w[27][28] ),
    .A2(\w[29][28] ),
    .A3(\w[31][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04057_));
 sky130_fd_sc_hd__mux4_2 _17481_ (.A0(\w[49][28] ),
    .A1(\w[51][28] ),
    .A2(\w[53][28] ),
    .A3(\w[55][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04059_));
 sky130_fd_sc_hd__mux4_2 _17482_ (.A0(\w[57][28] ),
    .A1(\w[59][28] ),
    .A2(\w[61][28] ),
    .A3(\w[63][28] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04060_));
 sky130_fd_sc_hd__mux4_2 _17483_ (.A0(_04056_),
    .A1(_04057_),
    .A2(_04059_),
    .A3(_04060_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04061_));
 sky130_fd_sc_hd__mux2_2 _17484_ (.A0(_04055_),
    .A1(_04061_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[28] ));
 sky130_fd_sc_hd__mux4_2 _17485_ (.A0(\w[1][29] ),
    .A1(\w[3][29] ),
    .A2(\w[5][29] ),
    .A3(\w[7][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04062_));
 sky130_fd_sc_hd__mux4_2 _17486_ (.A0(\w[9][29] ),
    .A1(\w[11][29] ),
    .A2(\w[13][29] ),
    .A3(\w[15][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04063_));
 sky130_fd_sc_hd__mux4_2 _17487_ (.A0(\w[33][29] ),
    .A1(\w[35][29] ),
    .A2(\w[37][29] ),
    .A3(\w[39][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04064_));
 sky130_fd_sc_hd__mux4_2 _17488_ (.A0(\w[41][29] ),
    .A1(\w[43][29] ),
    .A2(\w[45][29] ),
    .A3(\w[47][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04065_));
 sky130_fd_sc_hd__mux4_2 _17489_ (.A0(_04062_),
    .A1(_04063_),
    .A2(_04064_),
    .A3(_04065_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04066_));
 sky130_fd_sc_hd__mux4_2 _17490_ (.A0(\w[17][29] ),
    .A1(\w[19][29] ),
    .A2(\w[21][29] ),
    .A3(\w[23][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04067_));
 sky130_fd_sc_hd__mux4_2 _17491_ (.A0(\w[25][29] ),
    .A1(\w[27][29] ),
    .A2(\w[29][29] ),
    .A3(\w[31][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04068_));
 sky130_fd_sc_hd__mux4_2 _17493_ (.A0(\w[49][29] ),
    .A1(\w[51][29] ),
    .A2(\w[53][29] ),
    .A3(\w[55][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04070_));
 sky130_fd_sc_hd__mux4_2 _17494_ (.A0(\w[57][29] ),
    .A1(\w[59][29] ),
    .A2(\w[61][29] ),
    .A3(\w[63][29] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04071_));
 sky130_fd_sc_hd__mux4_2 _17495_ (.A0(_04067_),
    .A1(_04068_),
    .A2(_04070_),
    .A3(_04071_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04072_));
 sky130_fd_sc_hd__mux2_2 _17496_ (.A0(_04066_),
    .A1(_04072_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[29] ));
 sky130_fd_sc_hd__mux4_2 _17498_ (.A0(\w[1][2] ),
    .A1(\w[3][2] ),
    .A2(\w[5][2] ),
    .A3(\w[7][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04074_));
 sky130_fd_sc_hd__mux4_2 _17499_ (.A0(\w[9][2] ),
    .A1(\w[11][2] ),
    .A2(\w[13][2] ),
    .A3(\w[15][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04075_));
 sky130_fd_sc_hd__mux4_2 _17500_ (.A0(\w[33][2] ),
    .A1(\w[35][2] ),
    .A2(\w[37][2] ),
    .A3(\w[39][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04076_));
 sky130_fd_sc_hd__mux4_2 _17501_ (.A0(\w[41][2] ),
    .A1(\w[43][2] ),
    .A2(\w[45][2] ),
    .A3(\w[47][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04077_));
 sky130_fd_sc_hd__mux4_2 _17502_ (.A0(_04074_),
    .A1(_04075_),
    .A2(_04076_),
    .A3(_04077_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04078_));
 sky130_fd_sc_hd__mux4_2 _17503_ (.A0(\w[17][2] ),
    .A1(\w[19][2] ),
    .A2(\w[21][2] ),
    .A3(\w[23][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04079_));
 sky130_fd_sc_hd__mux4_2 _17504_ (.A0(\w[25][2] ),
    .A1(\w[27][2] ),
    .A2(\w[29][2] ),
    .A3(\w[31][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04080_));
 sky130_fd_sc_hd__mux4_2 _17505_ (.A0(\w[49][2] ),
    .A1(\w[51][2] ),
    .A2(\w[53][2] ),
    .A3(\w[55][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04081_));
 sky130_fd_sc_hd__mux4_2 _17506_ (.A0(\w[57][2] ),
    .A1(\w[59][2] ),
    .A2(\w[61][2] ),
    .A3(\w[63][2] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04082_));
 sky130_fd_sc_hd__mux4_2 _17507_ (.A0(_04079_),
    .A1(_04080_),
    .A2(_04081_),
    .A3(_04082_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04083_));
 sky130_fd_sc_hd__mux2_2 _17508_ (.A0(_04078_),
    .A1(_04083_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[2] ));
 sky130_fd_sc_hd__mux4_2 _17509_ (.A0(\w[1][30] ),
    .A1(\w[3][30] ),
    .A2(\w[5][30] ),
    .A3(\w[7][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04084_));
 sky130_fd_sc_hd__mux4_2 _17510_ (.A0(\w[9][30] ),
    .A1(\w[11][30] ),
    .A2(\w[13][30] ),
    .A3(\w[15][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04085_));
 sky130_fd_sc_hd__mux4_2 _17511_ (.A0(\w[33][30] ),
    .A1(\w[35][30] ),
    .A2(\w[37][30] ),
    .A3(\w[39][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04086_));
 sky130_fd_sc_hd__mux4_2 _17512_ (.A0(\w[41][30] ),
    .A1(\w[43][30] ),
    .A2(\w[45][30] ),
    .A3(\w[47][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04087_));
 sky130_fd_sc_hd__mux4_2 _17513_ (.A0(_04084_),
    .A1(_04085_),
    .A2(_04086_),
    .A3(_04087_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04088_));
 sky130_fd_sc_hd__mux4_2 _17514_ (.A0(\w[17][30] ),
    .A1(\w[19][30] ),
    .A2(\w[21][30] ),
    .A3(\w[23][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04089_));
 sky130_fd_sc_hd__mux4_2 _17515_ (.A0(\w[25][30] ),
    .A1(\w[27][30] ),
    .A2(\w[29][30] ),
    .A3(\w[31][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04090_));
 sky130_fd_sc_hd__mux4_2 _17516_ (.A0(\w[49][30] ),
    .A1(\w[51][30] ),
    .A2(\w[53][30] ),
    .A3(\w[55][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04091_));
 sky130_fd_sc_hd__mux4_2 _17517_ (.A0(\w[57][30] ),
    .A1(\w[59][30] ),
    .A2(\w[61][30] ),
    .A3(\w[63][30] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04092_));
 sky130_fd_sc_hd__mux4_2 _17518_ (.A0(_04089_),
    .A1(_04090_),
    .A2(_04091_),
    .A3(_04092_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04093_));
 sky130_fd_sc_hd__mux2_2 _17519_ (.A0(_04088_),
    .A1(_04093_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[30] ));
 sky130_fd_sc_hd__mux4_2 _17520_ (.A0(\w[1][31] ),
    .A1(\w[3][31] ),
    .A2(\w[5][31] ),
    .A3(\w[7][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04094_));
 sky130_fd_sc_hd__mux4_2 _17521_ (.A0(\w[9][31] ),
    .A1(\w[11][31] ),
    .A2(\w[13][31] ),
    .A3(\w[15][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04095_));
 sky130_fd_sc_hd__mux4_2 _17522_ (.A0(\w[33][31] ),
    .A1(\w[35][31] ),
    .A2(\w[37][31] ),
    .A3(\w[39][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04096_));
 sky130_fd_sc_hd__mux4_2 _17523_ (.A0(\w[41][31] ),
    .A1(\w[43][31] ),
    .A2(\w[45][31] ),
    .A3(\w[47][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04097_));
 sky130_fd_sc_hd__mux4_2 _17524_ (.A0(_04094_),
    .A1(_04095_),
    .A2(_04096_),
    .A3(_04097_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04098_));
 sky130_fd_sc_hd__mux4_2 _17525_ (.A0(\w[17][31] ),
    .A1(\w[19][31] ),
    .A2(\w[21][31] ),
    .A3(\w[23][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04099_));
 sky130_fd_sc_hd__mux4_2 _17526_ (.A0(\w[25][31] ),
    .A1(\w[27][31] ),
    .A2(\w[29][31] ),
    .A3(\w[31][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04100_));
 sky130_fd_sc_hd__mux4_2 _17527_ (.A0(\w[49][31] ),
    .A1(\w[51][31] ),
    .A2(\w[53][31] ),
    .A3(\w[55][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04101_));
 sky130_fd_sc_hd__mux4_2 _17528_ (.A0(\w[57][31] ),
    .A1(\w[59][31] ),
    .A2(\w[61][31] ),
    .A3(\w[63][31] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04102_));
 sky130_fd_sc_hd__mux4_2 _17529_ (.A0(_04099_),
    .A1(_04100_),
    .A2(_04101_),
    .A3(_04102_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04103_));
 sky130_fd_sc_hd__mux2_2 _17530_ (.A0(_04098_),
    .A1(_04103_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[31] ));
 sky130_fd_sc_hd__mux4_2 _17531_ (.A0(\w[1][3] ),
    .A1(\w[3][3] ),
    .A2(\w[5][3] ),
    .A3(\w[7][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04104_));
 sky130_fd_sc_hd__mux4_2 _17532_ (.A0(\w[9][3] ),
    .A1(\w[11][3] ),
    .A2(\w[13][3] ),
    .A3(\w[15][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04105_));
 sky130_fd_sc_hd__mux4_2 _17533_ (.A0(\w[33][3] ),
    .A1(\w[35][3] ),
    .A2(\w[37][3] ),
    .A3(\w[39][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04106_));
 sky130_fd_sc_hd__mux4_2 _17534_ (.A0(\w[41][3] ),
    .A1(\w[43][3] ),
    .A2(\w[45][3] ),
    .A3(\w[47][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04107_));
 sky130_fd_sc_hd__mux4_2 _17535_ (.A0(_04104_),
    .A1(_04105_),
    .A2(_04106_),
    .A3(_04107_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04108_));
 sky130_fd_sc_hd__mux4_2 _17536_ (.A0(\w[17][3] ),
    .A1(\w[19][3] ),
    .A2(\w[21][3] ),
    .A3(\w[23][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04109_));
 sky130_fd_sc_hd__mux4_2 _17537_ (.A0(\w[25][3] ),
    .A1(\w[27][3] ),
    .A2(\w[29][3] ),
    .A3(\w[31][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04110_));
 sky130_fd_sc_hd__mux4_2 _17538_ (.A0(\w[49][3] ),
    .A1(\w[51][3] ),
    .A2(\w[53][3] ),
    .A3(\w[55][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04111_));
 sky130_fd_sc_hd__mux4_2 _17539_ (.A0(\w[57][3] ),
    .A1(\w[59][3] ),
    .A2(\w[61][3] ),
    .A3(\w[63][3] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04112_));
 sky130_fd_sc_hd__mux4_2 _17540_ (.A0(_04109_),
    .A1(_04110_),
    .A2(_04111_),
    .A3(_04112_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04113_));
 sky130_fd_sc_hd__mux2_2 _17541_ (.A0(_04108_),
    .A1(_04113_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[3] ));
 sky130_fd_sc_hd__mux4_2 _17542_ (.A0(\w[1][4] ),
    .A1(\w[3][4] ),
    .A2(\w[5][4] ),
    .A3(\w[7][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04114_));
 sky130_fd_sc_hd__mux4_2 _17543_ (.A0(\w[9][4] ),
    .A1(\w[11][4] ),
    .A2(\w[13][4] ),
    .A3(\w[15][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04115_));
 sky130_fd_sc_hd__mux4_2 _17544_ (.A0(\w[33][4] ),
    .A1(\w[35][4] ),
    .A2(\w[37][4] ),
    .A3(\w[39][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04116_));
 sky130_fd_sc_hd__mux4_2 _17545_ (.A0(\w[41][4] ),
    .A1(\w[43][4] ),
    .A2(\w[45][4] ),
    .A3(\w[47][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04117_));
 sky130_fd_sc_hd__mux4_2 _17546_ (.A0(_04114_),
    .A1(_04115_),
    .A2(_04116_),
    .A3(_04117_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04118_));
 sky130_fd_sc_hd__mux4_2 _17547_ (.A0(\w[17][4] ),
    .A1(\w[19][4] ),
    .A2(\w[21][4] ),
    .A3(\w[23][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04119_));
 sky130_fd_sc_hd__mux4_2 _17548_ (.A0(\w[25][4] ),
    .A1(\w[27][4] ),
    .A2(\w[29][4] ),
    .A3(\w[31][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04120_));
 sky130_fd_sc_hd__mux4_2 _17549_ (.A0(\w[49][4] ),
    .A1(\w[51][4] ),
    .A2(\w[53][4] ),
    .A3(\w[55][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04121_));
 sky130_fd_sc_hd__mux4_2 _17550_ (.A0(\w[57][4] ),
    .A1(\w[59][4] ),
    .A2(\w[61][4] ),
    .A3(\w[63][4] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04122_));
 sky130_fd_sc_hd__mux4_2 _17551_ (.A0(_04119_),
    .A1(_04120_),
    .A2(_04121_),
    .A3(_04122_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04123_));
 sky130_fd_sc_hd__mux2_2 _17552_ (.A0(_04118_),
    .A1(_04123_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[4] ));
 sky130_fd_sc_hd__mux4_2 _17553_ (.A0(\w[1][5] ),
    .A1(\w[3][5] ),
    .A2(\w[5][5] ),
    .A3(\w[7][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04124_));
 sky130_fd_sc_hd__mux4_2 _17554_ (.A0(\w[9][5] ),
    .A1(\w[11][5] ),
    .A2(\w[13][5] ),
    .A3(\w[15][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04125_));
 sky130_fd_sc_hd__mux4_2 _17555_ (.A0(\w[33][5] ),
    .A1(\w[35][5] ),
    .A2(\w[37][5] ),
    .A3(\w[39][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04126_));
 sky130_fd_sc_hd__mux4_2 _17556_ (.A0(\w[41][5] ),
    .A1(\w[43][5] ),
    .A2(\w[45][5] ),
    .A3(\w[47][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04127_));
 sky130_fd_sc_hd__mux4_2 _17557_ (.A0(_04124_),
    .A1(_04125_),
    .A2(_04126_),
    .A3(_04127_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04128_));
 sky130_fd_sc_hd__mux4_2 _17558_ (.A0(\w[17][5] ),
    .A1(\w[19][5] ),
    .A2(\w[21][5] ),
    .A3(\w[23][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04129_));
 sky130_fd_sc_hd__mux4_2 _17559_ (.A0(\w[25][5] ),
    .A1(\w[27][5] ),
    .A2(\w[29][5] ),
    .A3(\w[31][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04130_));
 sky130_fd_sc_hd__mux4_2 _17560_ (.A0(\w[49][5] ),
    .A1(\w[51][5] ),
    .A2(\w[53][5] ),
    .A3(\w[55][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04131_));
 sky130_fd_sc_hd__mux4_2 _17561_ (.A0(\w[57][5] ),
    .A1(\w[59][5] ),
    .A2(\w[61][5] ),
    .A3(\w[63][5] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04132_));
 sky130_fd_sc_hd__mux4_2 _17562_ (.A0(_04129_),
    .A1(_04130_),
    .A2(_04131_),
    .A3(_04132_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04133_));
 sky130_fd_sc_hd__mux2_2 _17563_ (.A0(_04128_),
    .A1(_04133_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[5] ));
 sky130_fd_sc_hd__mux4_2 _17564_ (.A0(\w[1][6] ),
    .A1(\w[3][6] ),
    .A2(\w[5][6] ),
    .A3(\w[7][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04134_));
 sky130_fd_sc_hd__mux4_2 _17565_ (.A0(\w[9][6] ),
    .A1(\w[11][6] ),
    .A2(\w[13][6] ),
    .A3(\w[15][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04135_));
 sky130_fd_sc_hd__mux4_2 _17566_ (.A0(\w[33][6] ),
    .A1(\w[35][6] ),
    .A2(\w[37][6] ),
    .A3(\w[39][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04136_));
 sky130_fd_sc_hd__mux4_2 _17567_ (.A0(\w[41][6] ),
    .A1(\w[43][6] ),
    .A2(\w[45][6] ),
    .A3(\w[47][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04137_));
 sky130_fd_sc_hd__mux4_2 _17568_ (.A0(_04134_),
    .A1(_04135_),
    .A2(_04136_),
    .A3(_04137_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04138_));
 sky130_fd_sc_hd__mux4_2 _17569_ (.A0(\w[17][6] ),
    .A1(\w[19][6] ),
    .A2(\w[21][6] ),
    .A3(\w[23][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04139_));
 sky130_fd_sc_hd__mux4_2 _17570_ (.A0(\w[25][6] ),
    .A1(\w[27][6] ),
    .A2(\w[29][6] ),
    .A3(\w[31][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04140_));
 sky130_fd_sc_hd__mux4_2 _17571_ (.A0(\w[49][6] ),
    .A1(\w[51][6] ),
    .A2(\w[53][6] ),
    .A3(\w[55][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04141_));
 sky130_fd_sc_hd__mux4_2 _17572_ (.A0(\w[57][6] ),
    .A1(\w[59][6] ),
    .A2(\w[61][6] ),
    .A3(\w[63][6] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04142_));
 sky130_fd_sc_hd__mux4_2 _17573_ (.A0(_04139_),
    .A1(_04140_),
    .A2(_04141_),
    .A3(_04142_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04143_));
 sky130_fd_sc_hd__mux2_2 _17574_ (.A0(_04138_),
    .A1(_04143_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[6] ));
 sky130_fd_sc_hd__mux4_2 _17575_ (.A0(\w[1][7] ),
    .A1(\w[3][7] ),
    .A2(\w[5][7] ),
    .A3(\w[7][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04144_));
 sky130_fd_sc_hd__mux4_2 _17576_ (.A0(\w[9][7] ),
    .A1(\w[11][7] ),
    .A2(\w[13][7] ),
    .A3(\w[15][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04145_));
 sky130_fd_sc_hd__mux4_2 _17577_ (.A0(\w[33][7] ),
    .A1(\w[35][7] ),
    .A2(\w[37][7] ),
    .A3(\w[39][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04146_));
 sky130_fd_sc_hd__mux4_2 _17578_ (.A0(\w[41][7] ),
    .A1(\w[43][7] ),
    .A2(\w[45][7] ),
    .A3(\w[47][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04147_));
 sky130_fd_sc_hd__mux4_2 _17579_ (.A0(_04144_),
    .A1(_04145_),
    .A2(_04146_),
    .A3(_04147_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04148_));
 sky130_fd_sc_hd__mux4_2 _17580_ (.A0(\w[17][7] ),
    .A1(\w[19][7] ),
    .A2(\w[21][7] ),
    .A3(\w[23][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04149_));
 sky130_fd_sc_hd__mux4_2 _17581_ (.A0(\w[25][7] ),
    .A1(\w[27][7] ),
    .A2(\w[29][7] ),
    .A3(\w[31][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04150_));
 sky130_fd_sc_hd__mux4_2 _17582_ (.A0(\w[49][7] ),
    .A1(\w[51][7] ),
    .A2(\w[53][7] ),
    .A3(\w[55][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04151_));
 sky130_fd_sc_hd__mux4_2 _17583_ (.A0(\w[57][7] ),
    .A1(\w[59][7] ),
    .A2(\w[61][7] ),
    .A3(\w[63][7] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04152_));
 sky130_fd_sc_hd__mux4_2 _17584_ (.A0(_04149_),
    .A1(_04150_),
    .A2(_04151_),
    .A3(_04152_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04153_));
 sky130_fd_sc_hd__mux2_2 _17585_ (.A0(_04148_),
    .A1(_04153_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[7] ));
 sky130_fd_sc_hd__mux4_2 _17586_ (.A0(\w[1][8] ),
    .A1(\w[3][8] ),
    .A2(\w[5][8] ),
    .A3(\w[7][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04154_));
 sky130_fd_sc_hd__mux4_2 _17587_ (.A0(\w[9][8] ),
    .A1(\w[11][8] ),
    .A2(\w[13][8] ),
    .A3(\w[15][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04155_));
 sky130_fd_sc_hd__mux4_2 _17588_ (.A0(\w[33][8] ),
    .A1(\w[35][8] ),
    .A2(\w[37][8] ),
    .A3(\w[39][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04156_));
 sky130_fd_sc_hd__mux4_2 _17589_ (.A0(\w[41][8] ),
    .A1(\w[43][8] ),
    .A2(\w[45][8] ),
    .A3(\w[47][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04157_));
 sky130_fd_sc_hd__mux4_2 _17590_ (.A0(_04154_),
    .A1(_04155_),
    .A2(_04156_),
    .A3(_04157_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04158_));
 sky130_fd_sc_hd__mux4_2 _17591_ (.A0(\w[17][8] ),
    .A1(\w[19][8] ),
    .A2(\w[21][8] ),
    .A3(\w[23][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04159_));
 sky130_fd_sc_hd__mux4_2 _17592_ (.A0(\w[25][8] ),
    .A1(\w[27][8] ),
    .A2(\w[29][8] ),
    .A3(\w[31][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04160_));
 sky130_fd_sc_hd__mux4_2 _17593_ (.A0(\w[49][8] ),
    .A1(\w[51][8] ),
    .A2(\w[53][8] ),
    .A3(\w[55][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04161_));
 sky130_fd_sc_hd__mux4_2 _17594_ (.A0(\w[57][8] ),
    .A1(\w[59][8] ),
    .A2(\w[61][8] ),
    .A3(\w[63][8] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04162_));
 sky130_fd_sc_hd__mux4_2 _17595_ (.A0(_04159_),
    .A1(_04160_),
    .A2(_04161_),
    .A3(_04162_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_2 _17596_ (.A0(_04158_),
    .A1(_04163_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[8] ));
 sky130_fd_sc_hd__mux4_2 _17597_ (.A0(\w[1][9] ),
    .A1(\w[3][9] ),
    .A2(\w[5][9] ),
    .A3(\w[7][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04164_));
 sky130_fd_sc_hd__mux4_2 _17598_ (.A0(\w[9][9] ),
    .A1(\w[11][9] ),
    .A2(\w[13][9] ),
    .A3(\w[15][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04165_));
 sky130_fd_sc_hd__mux4_2 _17599_ (.A0(\w[33][9] ),
    .A1(\w[35][9] ),
    .A2(\w[37][9] ),
    .A3(\w[39][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04166_));
 sky130_fd_sc_hd__mux4_2 _17600_ (.A0(\w[41][9] ),
    .A1(\w[43][9] ),
    .A2(\w[45][9] ),
    .A3(\w[47][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04167_));
 sky130_fd_sc_hd__mux4_2 _17601_ (.A0(_04164_),
    .A1(_04165_),
    .A2(_04166_),
    .A3(_04167_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04168_));
 sky130_fd_sc_hd__mux4_2 _17602_ (.A0(\w[17][9] ),
    .A1(\w[19][9] ),
    .A2(\w[21][9] ),
    .A3(\w[23][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04169_));
 sky130_fd_sc_hd__mux4_2 _17603_ (.A0(\w[25][9] ),
    .A1(\w[27][9] ),
    .A2(\w[29][9] ),
    .A3(\w[31][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04170_));
 sky130_fd_sc_hd__mux4_2 _17604_ (.A0(\w[49][9] ),
    .A1(\w[51][9] ),
    .A2(\w[53][9] ),
    .A3(\w[55][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04171_));
 sky130_fd_sc_hd__mux4_2 _17605_ (.A0(\w[57][9] ),
    .A1(\w[59][9] ),
    .A2(\w[61][9] ),
    .A3(\w[63][9] ),
    .S0(\count15_1[1] ),
    .S1(\count15_1[2] ),
    .X(_04172_));
 sky130_fd_sc_hd__mux4_2 _17606_ (.A0(_04169_),
    .A1(_04170_),
    .A2(_04171_),
    .A3(_04172_),
    .S0(\count15_1[3] ),
    .S1(\count15_1[5] ),
    .X(_04173_));
 sky130_fd_sc_hd__mux2_2 _17607_ (.A0(_04168_),
    .A1(_04173_),
    .S(\count15_1[4] ),
    .X(\w_new_calc1.w_15[9] ));
 sky130_fd_sc_hd__mux4_2 _17612_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04178_));
 sky130_fd_sc_hd__mux4_2 _17616_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04182_));
 sky130_fd_sc_hd__mux4_2 _17620_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04186_));
 sky130_fd_sc_hd__mux4_2 _17623_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04189_));
 sky130_fd_sc_hd__mux4_2 _17627_ (.A0(_04178_),
    .A1(_04182_),
    .A2(_04186_),
    .A3(_04189_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04193_));
 sky130_fd_sc_hd__mux4_2 _17630_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04196_));
 sky130_fd_sc_hd__mux4_2 _17633_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04199_));
 sky130_fd_sc_hd__mux4_2 _17636_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04202_));
 sky130_fd_sc_hd__mux4_2 _17637_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04203_));
 sky130_fd_sc_hd__mux4_2 _17638_ (.A0(_04196_),
    .A1(_04199_),
    .A2(_04202_),
    .A3(_04203_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04204_));
 sky130_fd_sc_hd__mux2_2 _17639_ (.A0(_04193_),
    .A1(_04204_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[0] ));
 sky130_fd_sc_hd__mux4_2 _17640_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04205_));
 sky130_fd_sc_hd__mux4_2 _17641_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04206_));
 sky130_fd_sc_hd__mux4_2 _17642_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04207_));
 sky130_fd_sc_hd__mux4_2 _17643_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04208_));
 sky130_fd_sc_hd__mux4_2 _17644_ (.A0(_04205_),
    .A1(_04206_),
    .A2(_04207_),
    .A3(_04208_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04209_));
 sky130_fd_sc_hd__mux4_2 _17645_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04210_));
 sky130_fd_sc_hd__mux4_2 _17646_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04211_));
 sky130_fd_sc_hd__mux4_2 _17648_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04213_));
 sky130_fd_sc_hd__mux4_2 _17649_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04214_));
 sky130_fd_sc_hd__mux4_2 _17650_ (.A0(_04210_),
    .A1(_04211_),
    .A2(_04213_),
    .A3(_04214_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04215_));
 sky130_fd_sc_hd__mux2_2 _17651_ (.A0(_04209_),
    .A1(_04215_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[10] ));
 sky130_fd_sc_hd__mux4_2 _17653_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04217_));
 sky130_fd_sc_hd__mux4_2 _17654_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04218_));
 sky130_fd_sc_hd__mux4_2 _17655_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04219_));
 sky130_fd_sc_hd__mux4_2 _17656_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04220_));
 sky130_fd_sc_hd__mux4_2 _17657_ (.A0(_04217_),
    .A1(_04218_),
    .A2(_04219_),
    .A3(_04220_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04221_));
 sky130_fd_sc_hd__mux4_2 _17658_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04222_));
 sky130_fd_sc_hd__mux4_2 _17659_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04223_));
 sky130_fd_sc_hd__mux4_2 _17660_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04224_));
 sky130_fd_sc_hd__mux4_2 _17661_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04225_));
 sky130_fd_sc_hd__mux4_2 _17662_ (.A0(_04222_),
    .A1(_04223_),
    .A2(_04224_),
    .A3(_04225_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04226_));
 sky130_fd_sc_hd__mux2_2 _17663_ (.A0(_04221_),
    .A1(_04226_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[11] ));
 sky130_fd_sc_hd__mux4_2 _17665_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04228_));
 sky130_fd_sc_hd__mux4_2 _17666_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04229_));
 sky130_fd_sc_hd__mux4_2 _17667_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04230_));
 sky130_fd_sc_hd__mux4_2 _17668_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04231_));
 sky130_fd_sc_hd__mux4_2 _17669_ (.A0(_04228_),
    .A1(_04229_),
    .A2(_04230_),
    .A3(_04231_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04232_));
 sky130_fd_sc_hd__mux4_2 _17670_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04233_));
 sky130_fd_sc_hd__mux4_2 _17671_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04234_));
 sky130_fd_sc_hd__mux4_2 _17672_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04235_));
 sky130_fd_sc_hd__mux4_2 _17673_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04236_));
 sky130_fd_sc_hd__mux4_2 _17674_ (.A0(_04233_),
    .A1(_04234_),
    .A2(_04235_),
    .A3(_04236_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04237_));
 sky130_fd_sc_hd__mux2_2 _17675_ (.A0(_04232_),
    .A1(_04237_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[12] ));
 sky130_fd_sc_hd__mux4_2 _17676_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04238_));
 sky130_fd_sc_hd__mux4_2 _17678_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04240_));
 sky130_fd_sc_hd__mux4_2 _17679_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04241_));
 sky130_fd_sc_hd__mux4_2 _17680_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04242_));
 sky130_fd_sc_hd__mux4_2 _17681_ (.A0(_04238_),
    .A1(_04240_),
    .A2(_04241_),
    .A3(_04242_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04243_));
 sky130_fd_sc_hd__mux4_2 _17683_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04245_));
 sky130_fd_sc_hd__mux4_2 _17684_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04246_));
 sky130_fd_sc_hd__mux4_2 _17685_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04247_));
 sky130_fd_sc_hd__mux4_2 _17686_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04248_));
 sky130_fd_sc_hd__mux4_2 _17687_ (.A0(_04245_),
    .A1(_04246_),
    .A2(_04247_),
    .A3(_04248_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04249_));
 sky130_fd_sc_hd__mux2_2 _17688_ (.A0(_04243_),
    .A1(_04249_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[13] ));
 sky130_fd_sc_hd__mux4_2 _17689_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04250_));
 sky130_fd_sc_hd__mux4_2 _17691_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04252_));
 sky130_fd_sc_hd__mux4_2 _17692_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04253_));
 sky130_fd_sc_hd__mux4_2 _17693_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04254_));
 sky130_fd_sc_hd__mux4_2 _17695_ (.A0(_04250_),
    .A1(_04252_),
    .A2(_04253_),
    .A3(_04254_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04256_));
 sky130_fd_sc_hd__mux4_2 _17697_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04258_));
 sky130_fd_sc_hd__mux4_2 _17698_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04259_));
 sky130_fd_sc_hd__mux4_2 _17699_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04260_));
 sky130_fd_sc_hd__mux4_2 _17700_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04261_));
 sky130_fd_sc_hd__mux4_2 _17701_ (.A0(_04258_),
    .A1(_04259_),
    .A2(_04260_),
    .A3(_04261_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04262_));
 sky130_fd_sc_hd__mux2_2 _17702_ (.A0(_04256_),
    .A1(_04262_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[14] ));
 sky130_fd_sc_hd__mux4_2 _17703_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04263_));
 sky130_fd_sc_hd__mux4_2 _17704_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04264_));
 sky130_fd_sc_hd__mux4_2 _17705_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04265_));
 sky130_fd_sc_hd__mux4_2 _17707_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04267_));
 sky130_fd_sc_hd__mux4_2 _17708_ (.A0(_04263_),
    .A1(_04264_),
    .A2(_04265_),
    .A3(_04267_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04268_));
 sky130_fd_sc_hd__mux4_2 _17709_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04269_));
 sky130_fd_sc_hd__mux4_2 _17711_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04271_));
 sky130_fd_sc_hd__mux4_2 _17712_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04272_));
 sky130_fd_sc_hd__mux4_2 _17713_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04273_));
 sky130_fd_sc_hd__mux4_2 _17714_ (.A0(_04269_),
    .A1(_04271_),
    .A2(_04272_),
    .A3(_04273_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04274_));
 sky130_fd_sc_hd__mux2_2 _17715_ (.A0(_04268_),
    .A1(_04274_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[15] ));
 sky130_fd_sc_hd__mux4_2 _17716_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04275_));
 sky130_fd_sc_hd__mux4_2 _17717_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04276_));
 sky130_fd_sc_hd__mux4_2 _17718_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04277_));
 sky130_fd_sc_hd__mux4_2 _17720_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04279_));
 sky130_fd_sc_hd__mux4_2 _17722_ (.A0(_04275_),
    .A1(_04276_),
    .A2(_04277_),
    .A3(_04279_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04281_));
 sky130_fd_sc_hd__mux4_2 _17723_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04282_));
 sky130_fd_sc_hd__mux4_2 _17725_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04284_));
 sky130_fd_sc_hd__mux4_2 _17726_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04285_));
 sky130_fd_sc_hd__mux4_2 _17727_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04286_));
 sky130_fd_sc_hd__mux4_2 _17729_ (.A0(_04282_),
    .A1(_04284_),
    .A2(_04285_),
    .A3(_04286_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04288_));
 sky130_fd_sc_hd__mux2_2 _17730_ (.A0(_04281_),
    .A1(_04288_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[16] ));
 sky130_fd_sc_hd__mux4_2 _17731_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04289_));
 sky130_fd_sc_hd__mux4_2 _17732_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04290_));
 sky130_fd_sc_hd__mux4_2 _17734_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04292_));
 sky130_fd_sc_hd__mux4_2 _17735_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04293_));
 sky130_fd_sc_hd__mux4_2 _17736_ (.A0(_04289_),
    .A1(_04290_),
    .A2(_04292_),
    .A3(_04293_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04294_));
 sky130_fd_sc_hd__mux4_2 _17737_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04295_));
 sky130_fd_sc_hd__mux4_2 _17738_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04296_));
 sky130_fd_sc_hd__mux4_2 _17739_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04297_));
 sky130_fd_sc_hd__mux4_2 _17741_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04299_));
 sky130_fd_sc_hd__mux4_2 _17742_ (.A0(_04295_),
    .A1(_04296_),
    .A2(_04297_),
    .A3(_04299_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04300_));
 sky130_fd_sc_hd__mux2_2 _17743_ (.A0(_04294_),
    .A1(_04300_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[17] ));
 sky130_fd_sc_hd__mux4_2 _17744_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04301_));
 sky130_fd_sc_hd__mux4_2 _17745_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04302_));
 sky130_fd_sc_hd__mux4_2 _17747_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04304_));
 sky130_fd_sc_hd__mux4_2 _17748_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04305_));
 sky130_fd_sc_hd__mux4_2 _17749_ (.A0(_04301_),
    .A1(_04302_),
    .A2(_04304_),
    .A3(_04305_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04306_));
 sky130_fd_sc_hd__mux4_2 _17750_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04307_));
 sky130_fd_sc_hd__mux4_2 _17751_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04308_));
 sky130_fd_sc_hd__mux4_2 _17752_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04309_));
 sky130_fd_sc_hd__mux4_2 _17754_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04311_));
 sky130_fd_sc_hd__mux4_2 _17756_ (.A0(_04307_),
    .A1(_04308_),
    .A2(_04309_),
    .A3(_04311_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04313_));
 sky130_fd_sc_hd__mux2_2 _17758_ (.A0(_04306_),
    .A1(_04313_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[18] ));
 sky130_fd_sc_hd__mux4_2 _17759_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04315_));
 sky130_fd_sc_hd__mux4_2 _17760_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04316_));
 sky130_fd_sc_hd__mux4_2 _17761_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04317_));
 sky130_fd_sc_hd__mux4_2 _17762_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04318_));
 sky130_fd_sc_hd__mux4_2 _17763_ (.A0(_04315_),
    .A1(_04316_),
    .A2(_04317_),
    .A3(_04318_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04319_));
 sky130_fd_sc_hd__mux4_2 _17764_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04320_));
 sky130_fd_sc_hd__mux4_2 _17765_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04321_));
 sky130_fd_sc_hd__mux4_2 _17767_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04323_));
 sky130_fd_sc_hd__mux4_2 _17768_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04324_));
 sky130_fd_sc_hd__mux4_2 _17769_ (.A0(_04320_),
    .A1(_04321_),
    .A2(_04323_),
    .A3(_04324_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04325_));
 sky130_fd_sc_hd__mux2_2 _17770_ (.A0(_04319_),
    .A1(_04325_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[19] ));
 sky130_fd_sc_hd__mux4_2 _17771_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04326_));
 sky130_fd_sc_hd__mux4_2 _17772_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04327_));
 sky130_fd_sc_hd__mux4_2 _17773_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04328_));
 sky130_fd_sc_hd__mux4_2 _17774_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04329_));
 sky130_fd_sc_hd__mux4_2 _17775_ (.A0(_04326_),
    .A1(_04327_),
    .A2(_04328_),
    .A3(_04329_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04330_));
 sky130_fd_sc_hd__mux4_2 _17776_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04331_));
 sky130_fd_sc_hd__mux4_2 _17777_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04332_));
 sky130_fd_sc_hd__mux4_2 _17779_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04334_));
 sky130_fd_sc_hd__mux4_2 _17780_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04335_));
 sky130_fd_sc_hd__mux4_2 _17781_ (.A0(_04331_),
    .A1(_04332_),
    .A2(_04334_),
    .A3(_04335_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04336_));
 sky130_fd_sc_hd__mux2_2 _17782_ (.A0(_04330_),
    .A1(_04336_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[1] ));
 sky130_fd_sc_hd__mux4_2 _17784_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04338_));
 sky130_fd_sc_hd__mux4_2 _17785_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04339_));
 sky130_fd_sc_hd__mux4_2 _17786_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04340_));
 sky130_fd_sc_hd__mux4_2 _17787_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04341_));
 sky130_fd_sc_hd__mux4_2 _17788_ (.A0(_04338_),
    .A1(_04339_),
    .A2(_04340_),
    .A3(_04341_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04342_));
 sky130_fd_sc_hd__mux4_2 _17789_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04343_));
 sky130_fd_sc_hd__mux4_2 _17790_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04344_));
 sky130_fd_sc_hd__mux4_2 _17791_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04345_));
 sky130_fd_sc_hd__mux4_2 _17792_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04346_));
 sky130_fd_sc_hd__mux4_2 _17793_ (.A0(_04343_),
    .A1(_04344_),
    .A2(_04345_),
    .A3(_04346_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04347_));
 sky130_fd_sc_hd__mux2_2 _17794_ (.A0(_04342_),
    .A1(_04347_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[20] ));
 sky130_fd_sc_hd__mux4_2 _17796_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04349_));
 sky130_fd_sc_hd__mux4_2 _17797_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04350_));
 sky130_fd_sc_hd__mux4_2 _17798_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04351_));
 sky130_fd_sc_hd__mux4_2 _17799_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04352_));
 sky130_fd_sc_hd__mux4_2 _17800_ (.A0(_04349_),
    .A1(_04350_),
    .A2(_04351_),
    .A3(_04352_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04353_));
 sky130_fd_sc_hd__mux4_2 _17801_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04354_));
 sky130_fd_sc_hd__mux4_2 _17802_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04355_));
 sky130_fd_sc_hd__mux4_2 _17803_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04356_));
 sky130_fd_sc_hd__mux4_2 _17804_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04357_));
 sky130_fd_sc_hd__mux4_2 _17805_ (.A0(_04354_),
    .A1(_04355_),
    .A2(_04356_),
    .A3(_04357_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04358_));
 sky130_fd_sc_hd__mux2_2 _17806_ (.A0(_04353_),
    .A1(_04358_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[21] ));
 sky130_fd_sc_hd__mux4_2 _17807_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04359_));
 sky130_fd_sc_hd__mux4_2 _17809_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04361_));
 sky130_fd_sc_hd__mux4_2 _17810_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04362_));
 sky130_fd_sc_hd__mux4_2 _17811_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04363_));
 sky130_fd_sc_hd__mux4_2 _17812_ (.A0(_04359_),
    .A1(_04361_),
    .A2(_04362_),
    .A3(_04363_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04364_));
 sky130_fd_sc_hd__mux4_2 _17814_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04366_));
 sky130_fd_sc_hd__mux4_2 _17815_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04367_));
 sky130_fd_sc_hd__mux4_2 _17816_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04368_));
 sky130_fd_sc_hd__mux4_2 _17817_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04369_));
 sky130_fd_sc_hd__mux4_2 _17818_ (.A0(_04366_),
    .A1(_04367_),
    .A2(_04368_),
    .A3(_04369_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04370_));
 sky130_fd_sc_hd__mux2_2 _17819_ (.A0(_04364_),
    .A1(_04370_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[22] ));
 sky130_fd_sc_hd__mux4_2 _17820_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04371_));
 sky130_fd_sc_hd__mux4_2 _17822_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04373_));
 sky130_fd_sc_hd__mux4_2 _17823_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04374_));
 sky130_fd_sc_hd__mux4_2 _17824_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04375_));
 sky130_fd_sc_hd__mux4_2 _17826_ (.A0(_04371_),
    .A1(_04373_),
    .A2(_04374_),
    .A3(_04375_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04377_));
 sky130_fd_sc_hd__mux4_2 _17828_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04379_));
 sky130_fd_sc_hd__mux4_2 _17829_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04380_));
 sky130_fd_sc_hd__mux4_2 _17830_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04381_));
 sky130_fd_sc_hd__mux4_2 _17831_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04382_));
 sky130_fd_sc_hd__mux4_2 _17832_ (.A0(_04379_),
    .A1(_04380_),
    .A2(_04381_),
    .A3(_04382_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04383_));
 sky130_fd_sc_hd__mux2_2 _17833_ (.A0(_04377_),
    .A1(_04383_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[23] ));
 sky130_fd_sc_hd__mux4_2 _17834_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04384_));
 sky130_fd_sc_hd__mux4_2 _17835_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04385_));
 sky130_fd_sc_hd__mux4_2 _17836_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04386_));
 sky130_fd_sc_hd__mux4_2 _17838_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04388_));
 sky130_fd_sc_hd__mux4_2 _17839_ (.A0(_04384_),
    .A1(_04385_),
    .A2(_04386_),
    .A3(_04388_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04389_));
 sky130_fd_sc_hd__mux4_2 _17840_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04390_));
 sky130_fd_sc_hd__mux4_2 _17842_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04392_));
 sky130_fd_sc_hd__mux4_2 _17843_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04393_));
 sky130_fd_sc_hd__mux4_2 _17844_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04394_));
 sky130_fd_sc_hd__mux4_2 _17845_ (.A0(_04390_),
    .A1(_04392_),
    .A2(_04393_),
    .A3(_04394_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04395_));
 sky130_fd_sc_hd__mux2_2 _17846_ (.A0(_04389_),
    .A1(_04395_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[24] ));
 sky130_fd_sc_hd__mux4_2 _17847_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04396_));
 sky130_fd_sc_hd__mux4_2 _17848_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04397_));
 sky130_fd_sc_hd__mux4_2 _17849_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04398_));
 sky130_fd_sc_hd__mux4_2 _17851_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04400_));
 sky130_fd_sc_hd__mux4_2 _17853_ (.A0(_04396_),
    .A1(_04397_),
    .A2(_04398_),
    .A3(_04400_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04402_));
 sky130_fd_sc_hd__mux4_2 _17854_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04403_));
 sky130_fd_sc_hd__mux4_2 _17856_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04405_));
 sky130_fd_sc_hd__mux4_2 _17857_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04406_));
 sky130_fd_sc_hd__mux4_2 _17858_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04407_));
 sky130_fd_sc_hd__mux4_2 _17860_ (.A0(_04403_),
    .A1(_04405_),
    .A2(_04406_),
    .A3(_04407_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04409_));
 sky130_fd_sc_hd__mux2_2 _17861_ (.A0(_04402_),
    .A1(_04409_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[25] ));
 sky130_fd_sc_hd__mux4_2 _17862_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04410_));
 sky130_fd_sc_hd__mux4_2 _17863_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04411_));
 sky130_fd_sc_hd__mux4_2 _17865_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04413_));
 sky130_fd_sc_hd__mux4_2 _17866_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04414_));
 sky130_fd_sc_hd__mux4_2 _17867_ (.A0(_04410_),
    .A1(_04411_),
    .A2(_04413_),
    .A3(_04414_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04415_));
 sky130_fd_sc_hd__mux4_2 _17868_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04416_));
 sky130_fd_sc_hd__mux4_2 _17869_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04417_));
 sky130_fd_sc_hd__mux4_2 _17870_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04418_));
 sky130_fd_sc_hd__mux4_2 _17872_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04420_));
 sky130_fd_sc_hd__mux4_2 _17873_ (.A0(_04416_),
    .A1(_04417_),
    .A2(_04418_),
    .A3(_04420_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04421_));
 sky130_fd_sc_hd__mux2_2 _17874_ (.A0(_04415_),
    .A1(_04421_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[26] ));
 sky130_fd_sc_hd__mux4_2 _17875_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04422_));
 sky130_fd_sc_hd__mux4_2 _17876_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04423_));
 sky130_fd_sc_hd__mux4_2 _17878_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04425_));
 sky130_fd_sc_hd__mux4_2 _17879_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04426_));
 sky130_fd_sc_hd__mux4_2 _17880_ (.A0(_04422_),
    .A1(_04423_),
    .A2(_04425_),
    .A3(_04426_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04427_));
 sky130_fd_sc_hd__mux4_2 _17881_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04428_));
 sky130_fd_sc_hd__mux4_2 _17882_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04429_));
 sky130_fd_sc_hd__mux4_2 _17883_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04430_));
 sky130_fd_sc_hd__mux4_2 _17885_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04432_));
 sky130_fd_sc_hd__mux4_2 _17887_ (.A0(_04428_),
    .A1(_04429_),
    .A2(_04430_),
    .A3(_04432_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_2 _17889_ (.A0(_04427_),
    .A1(_04434_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[27] ));
 sky130_fd_sc_hd__mux4_2 _17890_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04436_));
 sky130_fd_sc_hd__mux4_2 _17891_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04437_));
 sky130_fd_sc_hd__mux4_2 _17892_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04438_));
 sky130_fd_sc_hd__mux4_2 _17893_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04439_));
 sky130_fd_sc_hd__mux4_2 _17894_ (.A0(_04436_),
    .A1(_04437_),
    .A2(_04438_),
    .A3(_04439_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04440_));
 sky130_fd_sc_hd__mux4_2 _17895_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04441_));
 sky130_fd_sc_hd__mux4_2 _17896_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04442_));
 sky130_fd_sc_hd__mux4_2 _17898_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04444_));
 sky130_fd_sc_hd__mux4_2 _17899_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04445_));
 sky130_fd_sc_hd__mux4_2 _17900_ (.A0(_04441_),
    .A1(_04442_),
    .A2(_04444_),
    .A3(_04445_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04446_));
 sky130_fd_sc_hd__mux2_2 _17901_ (.A0(_04440_),
    .A1(_04446_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[28] ));
 sky130_fd_sc_hd__mux4_2 _17902_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04447_));
 sky130_fd_sc_hd__mux4_2 _17903_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04448_));
 sky130_fd_sc_hd__mux4_2 _17904_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04449_));
 sky130_fd_sc_hd__mux4_2 _17905_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04450_));
 sky130_fd_sc_hd__mux4_2 _17906_ (.A0(_04447_),
    .A1(_04448_),
    .A2(_04449_),
    .A3(_04450_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04451_));
 sky130_fd_sc_hd__mux4_2 _17907_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04452_));
 sky130_fd_sc_hd__mux4_2 _17908_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04453_));
 sky130_fd_sc_hd__mux4_2 _17910_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04455_));
 sky130_fd_sc_hd__mux4_2 _17911_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04456_));
 sky130_fd_sc_hd__mux4_2 _17912_ (.A0(_04452_),
    .A1(_04453_),
    .A2(_04455_),
    .A3(_04456_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04457_));
 sky130_fd_sc_hd__mux2_2 _17913_ (.A0(_04451_),
    .A1(_04457_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[29] ));
 sky130_fd_sc_hd__mux4_2 _17915_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04459_));
 sky130_fd_sc_hd__mux4_2 _17916_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04460_));
 sky130_fd_sc_hd__mux4_2 _17917_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04461_));
 sky130_fd_sc_hd__mux4_2 _17918_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04462_));
 sky130_fd_sc_hd__mux4_2 _17919_ (.A0(_04459_),
    .A1(_04460_),
    .A2(_04461_),
    .A3(_04462_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04463_));
 sky130_fd_sc_hd__mux4_2 _17920_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04464_));
 sky130_fd_sc_hd__mux4_2 _17921_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04465_));
 sky130_fd_sc_hd__mux4_2 _17922_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04466_));
 sky130_fd_sc_hd__mux4_2 _17923_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04467_));
 sky130_fd_sc_hd__mux4_2 _17924_ (.A0(_04464_),
    .A1(_04465_),
    .A2(_04466_),
    .A3(_04467_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04468_));
 sky130_fd_sc_hd__mux2_2 _17925_ (.A0(_04463_),
    .A1(_04468_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[2] ));
 sky130_fd_sc_hd__mux4_2 _17926_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04469_));
 sky130_fd_sc_hd__mux4_2 _17927_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04470_));
 sky130_fd_sc_hd__mux4_2 _17928_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04471_));
 sky130_fd_sc_hd__mux4_2 _17929_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04472_));
 sky130_fd_sc_hd__mux4_2 _17930_ (.A0(_04469_),
    .A1(_04470_),
    .A2(_04471_),
    .A3(_04472_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04473_));
 sky130_fd_sc_hd__mux4_2 _17931_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04474_));
 sky130_fd_sc_hd__mux4_2 _17932_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04475_));
 sky130_fd_sc_hd__mux4_2 _17933_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04476_));
 sky130_fd_sc_hd__mux4_2 _17934_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04477_));
 sky130_fd_sc_hd__mux4_2 _17935_ (.A0(_04474_),
    .A1(_04475_),
    .A2(_04476_),
    .A3(_04477_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04478_));
 sky130_fd_sc_hd__mux2_2 _17936_ (.A0(_04473_),
    .A1(_04478_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[30] ));
 sky130_fd_sc_hd__mux4_2 _17937_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04479_));
 sky130_fd_sc_hd__mux4_2 _17938_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04480_));
 sky130_fd_sc_hd__mux4_2 _17939_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04481_));
 sky130_fd_sc_hd__mux4_2 _17940_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04482_));
 sky130_fd_sc_hd__mux4_2 _17941_ (.A0(_04479_),
    .A1(_04480_),
    .A2(_04481_),
    .A3(_04482_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04483_));
 sky130_fd_sc_hd__mux4_2 _17942_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04484_));
 sky130_fd_sc_hd__mux4_2 _17943_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04485_));
 sky130_fd_sc_hd__mux4_2 _17944_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04486_));
 sky130_fd_sc_hd__mux4_2 _17945_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04487_));
 sky130_fd_sc_hd__mux4_2 _17946_ (.A0(_04484_),
    .A1(_04485_),
    .A2(_04486_),
    .A3(_04487_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04488_));
 sky130_fd_sc_hd__mux2_2 _17947_ (.A0(_04483_),
    .A1(_04488_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[31] ));
 sky130_fd_sc_hd__mux4_2 _17948_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04489_));
 sky130_fd_sc_hd__mux4_2 _17949_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04490_));
 sky130_fd_sc_hd__mux4_2 _17950_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04491_));
 sky130_fd_sc_hd__mux4_2 _17951_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04492_));
 sky130_fd_sc_hd__mux4_2 _17952_ (.A0(_04489_),
    .A1(_04490_),
    .A2(_04491_),
    .A3(_04492_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04493_));
 sky130_fd_sc_hd__mux4_2 _17953_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04494_));
 sky130_fd_sc_hd__mux4_2 _17954_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04495_));
 sky130_fd_sc_hd__mux4_2 _17955_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04496_));
 sky130_fd_sc_hd__mux4_2 _17956_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04497_));
 sky130_fd_sc_hd__mux4_2 _17957_ (.A0(_04494_),
    .A1(_04495_),
    .A2(_04496_),
    .A3(_04497_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04498_));
 sky130_fd_sc_hd__mux2_2 _17958_ (.A0(_04493_),
    .A1(_04498_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[3] ));
 sky130_fd_sc_hd__mux4_2 _17959_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04499_));
 sky130_fd_sc_hd__mux4_2 _17960_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04500_));
 sky130_fd_sc_hd__mux4_2 _17961_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04501_));
 sky130_fd_sc_hd__mux4_2 _17962_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04502_));
 sky130_fd_sc_hd__mux4_2 _17963_ (.A0(_04499_),
    .A1(_04500_),
    .A2(_04501_),
    .A3(_04502_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04503_));
 sky130_fd_sc_hd__mux4_2 _17964_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04504_));
 sky130_fd_sc_hd__mux4_2 _17965_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04505_));
 sky130_fd_sc_hd__mux4_2 _17966_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04506_));
 sky130_fd_sc_hd__mux4_2 _17967_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04507_));
 sky130_fd_sc_hd__mux4_2 _17968_ (.A0(_04504_),
    .A1(_04505_),
    .A2(_04506_),
    .A3(_04507_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04508_));
 sky130_fd_sc_hd__mux2_2 _17969_ (.A0(_04503_),
    .A1(_04508_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[4] ));
 sky130_fd_sc_hd__mux4_2 _17970_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04509_));
 sky130_fd_sc_hd__mux4_2 _17971_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04510_));
 sky130_fd_sc_hd__mux4_2 _17972_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04511_));
 sky130_fd_sc_hd__mux4_2 _17973_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04512_));
 sky130_fd_sc_hd__mux4_2 _17974_ (.A0(_04509_),
    .A1(_04510_),
    .A2(_04511_),
    .A3(_04512_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04513_));
 sky130_fd_sc_hd__mux4_2 _17975_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04514_));
 sky130_fd_sc_hd__mux4_2 _17976_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04515_));
 sky130_fd_sc_hd__mux4_2 _17977_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04516_));
 sky130_fd_sc_hd__mux4_2 _17978_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04517_));
 sky130_fd_sc_hd__mux4_2 _17979_ (.A0(_04514_),
    .A1(_04515_),
    .A2(_04516_),
    .A3(_04517_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04518_));
 sky130_fd_sc_hd__mux2_2 _17980_ (.A0(_04513_),
    .A1(_04518_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[5] ));
 sky130_fd_sc_hd__mux4_2 _17981_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04519_));
 sky130_fd_sc_hd__mux4_2 _17982_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04520_));
 sky130_fd_sc_hd__mux4_2 _17983_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04521_));
 sky130_fd_sc_hd__mux4_2 _17984_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04522_));
 sky130_fd_sc_hd__mux4_2 _17985_ (.A0(_04519_),
    .A1(_04520_),
    .A2(_04521_),
    .A3(_04522_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04523_));
 sky130_fd_sc_hd__mux4_2 _17986_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04524_));
 sky130_fd_sc_hd__mux4_2 _17987_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04525_));
 sky130_fd_sc_hd__mux4_2 _17988_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04526_));
 sky130_fd_sc_hd__mux4_2 _17989_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04527_));
 sky130_fd_sc_hd__mux4_2 _17990_ (.A0(_04524_),
    .A1(_04525_),
    .A2(_04526_),
    .A3(_04527_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04528_));
 sky130_fd_sc_hd__mux2_2 _17991_ (.A0(_04523_),
    .A1(_04528_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[6] ));
 sky130_fd_sc_hd__mux4_2 _17992_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04529_));
 sky130_fd_sc_hd__mux4_2 _17993_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04530_));
 sky130_fd_sc_hd__mux4_2 _17994_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04531_));
 sky130_fd_sc_hd__mux4_2 _17995_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04532_));
 sky130_fd_sc_hd__mux4_2 _17996_ (.A0(_04529_),
    .A1(_04530_),
    .A2(_04531_),
    .A3(_04532_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04533_));
 sky130_fd_sc_hd__mux4_2 _17997_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04534_));
 sky130_fd_sc_hd__mux4_2 _17998_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04535_));
 sky130_fd_sc_hd__mux4_2 _17999_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04536_));
 sky130_fd_sc_hd__mux4_2 _18000_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04537_));
 sky130_fd_sc_hd__mux4_2 _18001_ (.A0(_04534_),
    .A1(_04535_),
    .A2(_04536_),
    .A3(_04537_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04538_));
 sky130_fd_sc_hd__mux2_2 _18002_ (.A0(_04533_),
    .A1(_04538_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[7] ));
 sky130_fd_sc_hd__mux4_2 _18003_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04539_));
 sky130_fd_sc_hd__mux4_2 _18004_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04540_));
 sky130_fd_sc_hd__mux4_2 _18005_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04541_));
 sky130_fd_sc_hd__mux4_2 _18006_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04542_));
 sky130_fd_sc_hd__mux4_2 _18007_ (.A0(_04539_),
    .A1(_04540_),
    .A2(_04541_),
    .A3(_04542_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04543_));
 sky130_fd_sc_hd__mux4_2 _18008_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04544_));
 sky130_fd_sc_hd__mux4_2 _18009_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04545_));
 sky130_fd_sc_hd__mux4_2 _18010_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04546_));
 sky130_fd_sc_hd__mux4_2 _18011_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04547_));
 sky130_fd_sc_hd__mux4_2 _18012_ (.A0(_04544_),
    .A1(_04545_),
    .A2(_04546_),
    .A3(_04547_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04548_));
 sky130_fd_sc_hd__mux2_2 _18013_ (.A0(_04543_),
    .A1(_04548_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[8] ));
 sky130_fd_sc_hd__mux4_2 _18014_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04549_));
 sky130_fd_sc_hd__mux4_2 _18015_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04550_));
 sky130_fd_sc_hd__mux4_2 _18016_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04551_));
 sky130_fd_sc_hd__mux4_2 _18017_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04552_));
 sky130_fd_sc_hd__mux4_2 _18018_ (.A0(_04549_),
    .A1(_04550_),
    .A2(_04551_),
    .A3(_04552_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04553_));
 sky130_fd_sc_hd__mux4_2 _18019_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04554_));
 sky130_fd_sc_hd__mux4_2 _18020_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04555_));
 sky130_fd_sc_hd__mux4_2 _18021_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04556_));
 sky130_fd_sc_hd__mux4_2 _18022_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_04557_));
 sky130_fd_sc_hd__mux4_2 _18023_ (.A0(_04554_),
    .A1(_04555_),
    .A2(_04556_),
    .A3(_04557_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[5] ),
    .X(_04558_));
 sky130_fd_sc_hd__mux2_2 _18024_ (.A0(_04553_),
    .A1(_04558_),
    .S(\count2_1[4] ),
    .X(\w_new_calc1.w_2[9] ));
 sky130_fd_sc_hd__mux4_2 _18029_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04563_));
 sky130_fd_sc_hd__mux4_2 _18033_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04567_));
 sky130_fd_sc_hd__mux4_2 _18037_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04571_));
 sky130_fd_sc_hd__mux4_2 _18040_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04574_));
 sky130_fd_sc_hd__mux4_2 _18044_ (.A0(_04563_),
    .A1(_04567_),
    .A2(_04571_),
    .A3(_04574_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04578_));
 sky130_fd_sc_hd__mux4_2 _18047_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04581_));
 sky130_fd_sc_hd__mux4_2 _18050_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04584_));
 sky130_fd_sc_hd__mux4_2 _18053_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04587_));
 sky130_fd_sc_hd__mux4_2 _18054_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04588_));
 sky130_fd_sc_hd__mux4_2 _18055_ (.A0(_04581_),
    .A1(_04584_),
    .A2(_04587_),
    .A3(_04588_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04589_));
 sky130_fd_sc_hd__mux2_2 _18056_ (.A0(_04578_),
    .A1(_04589_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[0] ));
 sky130_fd_sc_hd__mux4_2 _18057_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04590_));
 sky130_fd_sc_hd__mux4_2 _18058_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04591_));
 sky130_fd_sc_hd__mux4_2 _18059_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04592_));
 sky130_fd_sc_hd__mux4_2 _18060_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04593_));
 sky130_fd_sc_hd__mux4_2 _18061_ (.A0(_04590_),
    .A1(_04591_),
    .A2(_04592_),
    .A3(_04593_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04594_));
 sky130_fd_sc_hd__mux4_2 _18062_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04595_));
 sky130_fd_sc_hd__mux4_2 _18063_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04596_));
 sky130_fd_sc_hd__mux4_2 _18065_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04598_));
 sky130_fd_sc_hd__mux4_2 _18066_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04599_));
 sky130_fd_sc_hd__mux4_2 _18067_ (.A0(_04595_),
    .A1(_04596_),
    .A2(_04598_),
    .A3(_04599_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04600_));
 sky130_fd_sc_hd__mux2_2 _18068_ (.A0(_04594_),
    .A1(_04600_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[10] ));
 sky130_fd_sc_hd__mux4_2 _18070_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04602_));
 sky130_fd_sc_hd__mux4_2 _18071_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04603_));
 sky130_fd_sc_hd__mux4_2 _18072_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04604_));
 sky130_fd_sc_hd__mux4_2 _18073_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04605_));
 sky130_fd_sc_hd__mux4_2 _18074_ (.A0(_04602_),
    .A1(_04603_),
    .A2(_04604_),
    .A3(_04605_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04606_));
 sky130_fd_sc_hd__mux4_2 _18075_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04607_));
 sky130_fd_sc_hd__mux4_2 _18076_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04608_));
 sky130_fd_sc_hd__mux4_2 _18077_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04609_));
 sky130_fd_sc_hd__mux4_2 _18078_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04610_));
 sky130_fd_sc_hd__mux4_2 _18079_ (.A0(_04607_),
    .A1(_04608_),
    .A2(_04609_),
    .A3(_04610_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04611_));
 sky130_fd_sc_hd__mux2_2 _18080_ (.A0(_04606_),
    .A1(_04611_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[11] ));
 sky130_fd_sc_hd__mux4_2 _18082_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04613_));
 sky130_fd_sc_hd__mux4_2 _18083_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04614_));
 sky130_fd_sc_hd__mux4_2 _18084_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04615_));
 sky130_fd_sc_hd__mux4_2 _18085_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04616_));
 sky130_fd_sc_hd__mux4_2 _18086_ (.A0(_04613_),
    .A1(_04614_),
    .A2(_04615_),
    .A3(_04616_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04617_));
 sky130_fd_sc_hd__mux4_2 _18087_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04618_));
 sky130_fd_sc_hd__mux4_2 _18088_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04619_));
 sky130_fd_sc_hd__mux4_2 _18089_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04620_));
 sky130_fd_sc_hd__mux4_2 _18090_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04621_));
 sky130_fd_sc_hd__mux4_2 _18091_ (.A0(_04618_),
    .A1(_04619_),
    .A2(_04620_),
    .A3(_04621_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04622_));
 sky130_fd_sc_hd__mux2_2 _18092_ (.A0(_04617_),
    .A1(_04622_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[12] ));
 sky130_fd_sc_hd__mux4_2 _18093_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04623_));
 sky130_fd_sc_hd__mux4_2 _18095_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04625_));
 sky130_fd_sc_hd__mux4_2 _18096_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04626_));
 sky130_fd_sc_hd__mux4_2 _18097_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04627_));
 sky130_fd_sc_hd__mux4_2 _18098_ (.A0(_04623_),
    .A1(_04625_),
    .A2(_04626_),
    .A3(_04627_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04628_));
 sky130_fd_sc_hd__mux4_2 _18100_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04630_));
 sky130_fd_sc_hd__mux4_2 _18101_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04631_));
 sky130_fd_sc_hd__mux4_2 _18102_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04632_));
 sky130_fd_sc_hd__mux4_2 _18103_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04633_));
 sky130_fd_sc_hd__mux4_2 _18104_ (.A0(_04630_),
    .A1(_04631_),
    .A2(_04632_),
    .A3(_04633_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04634_));
 sky130_fd_sc_hd__mux2_2 _18105_ (.A0(_04628_),
    .A1(_04634_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[13] ));
 sky130_fd_sc_hd__mux4_2 _18106_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04635_));
 sky130_fd_sc_hd__mux4_2 _18108_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04637_));
 sky130_fd_sc_hd__mux4_2 _18109_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04638_));
 sky130_fd_sc_hd__mux4_2 _18110_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04639_));
 sky130_fd_sc_hd__mux4_2 _18112_ (.A0(_04635_),
    .A1(_04637_),
    .A2(_04638_),
    .A3(_04639_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04641_));
 sky130_fd_sc_hd__mux4_2 _18114_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04643_));
 sky130_fd_sc_hd__mux4_2 _18115_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04644_));
 sky130_fd_sc_hd__mux4_2 _18116_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04645_));
 sky130_fd_sc_hd__mux4_2 _18117_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04646_));
 sky130_fd_sc_hd__mux4_2 _18118_ (.A0(_04643_),
    .A1(_04644_),
    .A2(_04645_),
    .A3(_04646_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04647_));
 sky130_fd_sc_hd__mux2_2 _18119_ (.A0(_04641_),
    .A1(_04647_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[14] ));
 sky130_fd_sc_hd__mux4_2 _18120_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04648_));
 sky130_fd_sc_hd__mux4_2 _18121_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04649_));
 sky130_fd_sc_hd__mux4_2 _18122_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04650_));
 sky130_fd_sc_hd__mux4_2 _18124_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04652_));
 sky130_fd_sc_hd__mux4_2 _18125_ (.A0(_04648_),
    .A1(_04649_),
    .A2(_04650_),
    .A3(_04652_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04653_));
 sky130_fd_sc_hd__mux4_2 _18126_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04654_));
 sky130_fd_sc_hd__mux4_2 _18128_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04656_));
 sky130_fd_sc_hd__mux4_2 _18129_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04657_));
 sky130_fd_sc_hd__mux4_2 _18130_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04658_));
 sky130_fd_sc_hd__mux4_2 _18131_ (.A0(_04654_),
    .A1(_04656_),
    .A2(_04657_),
    .A3(_04658_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04659_));
 sky130_fd_sc_hd__mux2_2 _18132_ (.A0(_04653_),
    .A1(_04659_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[15] ));
 sky130_fd_sc_hd__mux4_2 _18133_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04660_));
 sky130_fd_sc_hd__mux4_2 _18134_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04661_));
 sky130_fd_sc_hd__mux4_2 _18135_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04662_));
 sky130_fd_sc_hd__mux4_2 _18137_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04664_));
 sky130_fd_sc_hd__mux4_2 _18139_ (.A0(_04660_),
    .A1(_04661_),
    .A2(_04662_),
    .A3(_04664_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04666_));
 sky130_fd_sc_hd__mux4_2 _18140_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04667_));
 sky130_fd_sc_hd__mux4_2 _18142_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04669_));
 sky130_fd_sc_hd__mux4_2 _18143_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04670_));
 sky130_fd_sc_hd__mux4_2 _18144_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04671_));
 sky130_fd_sc_hd__mux4_2 _18146_ (.A0(_04667_),
    .A1(_04669_),
    .A2(_04670_),
    .A3(_04671_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04673_));
 sky130_fd_sc_hd__mux2_2 _18147_ (.A0(_04666_),
    .A1(_04673_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[16] ));
 sky130_fd_sc_hd__mux4_2 _18148_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04674_));
 sky130_fd_sc_hd__mux4_2 _18149_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04675_));
 sky130_fd_sc_hd__mux4_2 _18151_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04677_));
 sky130_fd_sc_hd__mux4_2 _18152_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04678_));
 sky130_fd_sc_hd__mux4_2 _18153_ (.A0(_04674_),
    .A1(_04675_),
    .A2(_04677_),
    .A3(_04678_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04679_));
 sky130_fd_sc_hd__mux4_2 _18154_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04680_));
 sky130_fd_sc_hd__mux4_2 _18155_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04681_));
 sky130_fd_sc_hd__mux4_2 _18156_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04682_));
 sky130_fd_sc_hd__mux4_2 _18158_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04684_));
 sky130_fd_sc_hd__mux4_2 _18159_ (.A0(_04680_),
    .A1(_04681_),
    .A2(_04682_),
    .A3(_04684_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04685_));
 sky130_fd_sc_hd__mux2_2 _18160_ (.A0(_04679_),
    .A1(_04685_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[17] ));
 sky130_fd_sc_hd__mux4_2 _18161_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04686_));
 sky130_fd_sc_hd__mux4_2 _18162_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04687_));
 sky130_fd_sc_hd__mux4_2 _18164_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04689_));
 sky130_fd_sc_hd__mux4_2 _18165_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04690_));
 sky130_fd_sc_hd__mux4_2 _18166_ (.A0(_04686_),
    .A1(_04687_),
    .A2(_04689_),
    .A3(_04690_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04691_));
 sky130_fd_sc_hd__mux4_2 _18167_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04692_));
 sky130_fd_sc_hd__mux4_2 _18168_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04693_));
 sky130_fd_sc_hd__mux4_2 _18169_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04694_));
 sky130_fd_sc_hd__mux4_2 _18171_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04696_));
 sky130_fd_sc_hd__mux4_2 _18173_ (.A0(_04692_),
    .A1(_04693_),
    .A2(_04694_),
    .A3(_04696_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_2 _18175_ (.A0(_04691_),
    .A1(_04698_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[18] ));
 sky130_fd_sc_hd__mux4_2 _18176_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04700_));
 sky130_fd_sc_hd__mux4_2 _18177_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04701_));
 sky130_fd_sc_hd__mux4_2 _18178_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04702_));
 sky130_fd_sc_hd__mux4_2 _18179_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04703_));
 sky130_fd_sc_hd__mux4_2 _18180_ (.A0(_04700_),
    .A1(_04701_),
    .A2(_04702_),
    .A3(_04703_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04704_));
 sky130_fd_sc_hd__mux4_2 _18181_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04705_));
 sky130_fd_sc_hd__mux4_2 _18182_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04706_));
 sky130_fd_sc_hd__mux4_2 _18184_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04708_));
 sky130_fd_sc_hd__mux4_2 _18185_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04709_));
 sky130_fd_sc_hd__mux4_2 _18186_ (.A0(_04705_),
    .A1(_04706_),
    .A2(_04708_),
    .A3(_04709_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04710_));
 sky130_fd_sc_hd__mux2_2 _18187_ (.A0(_04704_),
    .A1(_04710_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[19] ));
 sky130_fd_sc_hd__mux4_2 _18188_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04711_));
 sky130_fd_sc_hd__mux4_2 _18189_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04712_));
 sky130_fd_sc_hd__mux4_2 _18190_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04713_));
 sky130_fd_sc_hd__mux4_2 _18191_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04714_));
 sky130_fd_sc_hd__mux4_2 _18192_ (.A0(_04711_),
    .A1(_04712_),
    .A2(_04713_),
    .A3(_04714_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04715_));
 sky130_fd_sc_hd__mux4_2 _18193_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04716_));
 sky130_fd_sc_hd__mux4_2 _18194_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04717_));
 sky130_fd_sc_hd__mux4_2 _18196_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04719_));
 sky130_fd_sc_hd__mux4_2 _18197_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04720_));
 sky130_fd_sc_hd__mux4_2 _18198_ (.A0(_04716_),
    .A1(_04717_),
    .A2(_04719_),
    .A3(_04720_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04721_));
 sky130_fd_sc_hd__mux2_2 _18199_ (.A0(_04715_),
    .A1(_04721_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[1] ));
 sky130_fd_sc_hd__mux4_2 _18201_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04723_));
 sky130_fd_sc_hd__mux4_2 _18202_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04724_));
 sky130_fd_sc_hd__mux4_2 _18203_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04725_));
 sky130_fd_sc_hd__mux4_2 _18204_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04726_));
 sky130_fd_sc_hd__mux4_2 _18205_ (.A0(_04723_),
    .A1(_04724_),
    .A2(_04725_),
    .A3(_04726_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04727_));
 sky130_fd_sc_hd__mux4_2 _18206_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04728_));
 sky130_fd_sc_hd__mux4_2 _18207_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04729_));
 sky130_fd_sc_hd__mux4_2 _18208_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04730_));
 sky130_fd_sc_hd__mux4_2 _18209_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04731_));
 sky130_fd_sc_hd__mux4_2 _18210_ (.A0(_04728_),
    .A1(_04729_),
    .A2(_04730_),
    .A3(_04731_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04732_));
 sky130_fd_sc_hd__mux2_2 _18211_ (.A0(_04727_),
    .A1(_04732_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[20] ));
 sky130_fd_sc_hd__mux4_2 _18213_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04734_));
 sky130_fd_sc_hd__mux4_2 _18214_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04735_));
 sky130_fd_sc_hd__mux4_2 _18215_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04736_));
 sky130_fd_sc_hd__mux4_2 _18216_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04737_));
 sky130_fd_sc_hd__mux4_2 _18217_ (.A0(_04734_),
    .A1(_04735_),
    .A2(_04736_),
    .A3(_04737_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04738_));
 sky130_fd_sc_hd__mux4_2 _18218_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04739_));
 sky130_fd_sc_hd__mux4_2 _18219_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04740_));
 sky130_fd_sc_hd__mux4_2 _18220_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04741_));
 sky130_fd_sc_hd__mux4_2 _18221_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04742_));
 sky130_fd_sc_hd__mux4_2 _18222_ (.A0(_04739_),
    .A1(_04740_),
    .A2(_04741_),
    .A3(_04742_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04743_));
 sky130_fd_sc_hd__mux2_2 _18223_ (.A0(_04738_),
    .A1(_04743_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[21] ));
 sky130_fd_sc_hd__mux4_2 _18224_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04744_));
 sky130_fd_sc_hd__mux4_2 _18226_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04746_));
 sky130_fd_sc_hd__mux4_2 _18227_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04747_));
 sky130_fd_sc_hd__mux4_2 _18228_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04748_));
 sky130_fd_sc_hd__mux4_2 _18229_ (.A0(_04744_),
    .A1(_04746_),
    .A2(_04747_),
    .A3(_04748_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04749_));
 sky130_fd_sc_hd__mux4_2 _18231_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04751_));
 sky130_fd_sc_hd__mux4_2 _18232_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04752_));
 sky130_fd_sc_hd__mux4_2 _18233_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04753_));
 sky130_fd_sc_hd__mux4_2 _18234_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04754_));
 sky130_fd_sc_hd__mux4_2 _18235_ (.A0(_04751_),
    .A1(_04752_),
    .A2(_04753_),
    .A3(_04754_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04755_));
 sky130_fd_sc_hd__mux2_2 _18236_ (.A0(_04749_),
    .A1(_04755_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[22] ));
 sky130_fd_sc_hd__mux4_2 _18237_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04756_));
 sky130_fd_sc_hd__mux4_2 _18239_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04758_));
 sky130_fd_sc_hd__mux4_2 _18240_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04759_));
 sky130_fd_sc_hd__mux4_2 _18241_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04760_));
 sky130_fd_sc_hd__mux4_2 _18243_ (.A0(_04756_),
    .A1(_04758_),
    .A2(_04759_),
    .A3(_04760_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04762_));
 sky130_fd_sc_hd__mux4_2 _18245_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04764_));
 sky130_fd_sc_hd__mux4_2 _18246_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04765_));
 sky130_fd_sc_hd__mux4_2 _18247_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04766_));
 sky130_fd_sc_hd__mux4_2 _18248_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04767_));
 sky130_fd_sc_hd__mux4_2 _18249_ (.A0(_04764_),
    .A1(_04765_),
    .A2(_04766_),
    .A3(_04767_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04768_));
 sky130_fd_sc_hd__mux2_2 _18250_ (.A0(_04762_),
    .A1(_04768_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[23] ));
 sky130_fd_sc_hd__mux4_2 _18251_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04769_));
 sky130_fd_sc_hd__mux4_2 _18252_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04770_));
 sky130_fd_sc_hd__mux4_2 _18253_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04771_));
 sky130_fd_sc_hd__mux4_2 _18255_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04773_));
 sky130_fd_sc_hd__mux4_2 _18256_ (.A0(_04769_),
    .A1(_04770_),
    .A2(_04771_),
    .A3(_04773_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04774_));
 sky130_fd_sc_hd__mux4_2 _18257_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04775_));
 sky130_fd_sc_hd__mux4_2 _18259_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04777_));
 sky130_fd_sc_hd__mux4_2 _18260_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04778_));
 sky130_fd_sc_hd__mux4_2 _18261_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04779_));
 sky130_fd_sc_hd__mux4_2 _18262_ (.A0(_04775_),
    .A1(_04777_),
    .A2(_04778_),
    .A3(_04779_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_2 _18263_ (.A0(_04774_),
    .A1(_04780_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[24] ));
 sky130_fd_sc_hd__mux4_2 _18264_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04781_));
 sky130_fd_sc_hd__mux4_2 _18265_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04782_));
 sky130_fd_sc_hd__mux4_2 _18266_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04783_));
 sky130_fd_sc_hd__mux4_2 _18268_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04785_));
 sky130_fd_sc_hd__mux4_2 _18270_ (.A0(_04781_),
    .A1(_04782_),
    .A2(_04783_),
    .A3(_04785_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04787_));
 sky130_fd_sc_hd__mux4_2 _18271_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04788_));
 sky130_fd_sc_hd__mux4_2 _18273_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04790_));
 sky130_fd_sc_hd__mux4_2 _18274_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04791_));
 sky130_fd_sc_hd__mux4_2 _18275_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04792_));
 sky130_fd_sc_hd__mux4_2 _18277_ (.A0(_04788_),
    .A1(_04790_),
    .A2(_04791_),
    .A3(_04792_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04794_));
 sky130_fd_sc_hd__mux2_2 _18278_ (.A0(_04787_),
    .A1(_04794_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[25] ));
 sky130_fd_sc_hd__mux4_2 _18279_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04795_));
 sky130_fd_sc_hd__mux4_2 _18280_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04796_));
 sky130_fd_sc_hd__mux4_2 _18282_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04798_));
 sky130_fd_sc_hd__mux4_2 _18283_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04799_));
 sky130_fd_sc_hd__mux4_2 _18284_ (.A0(_04795_),
    .A1(_04796_),
    .A2(_04798_),
    .A3(_04799_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04800_));
 sky130_fd_sc_hd__mux4_2 _18285_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04801_));
 sky130_fd_sc_hd__mux4_2 _18286_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04802_));
 sky130_fd_sc_hd__mux4_2 _18287_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04803_));
 sky130_fd_sc_hd__mux4_2 _18289_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04805_));
 sky130_fd_sc_hd__mux4_2 _18290_ (.A0(_04801_),
    .A1(_04802_),
    .A2(_04803_),
    .A3(_04805_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04806_));
 sky130_fd_sc_hd__mux2_2 _18291_ (.A0(_04800_),
    .A1(_04806_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[26] ));
 sky130_fd_sc_hd__mux4_2 _18292_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04807_));
 sky130_fd_sc_hd__mux4_2 _18293_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04808_));
 sky130_fd_sc_hd__mux4_2 _18295_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04810_));
 sky130_fd_sc_hd__mux4_2 _18296_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04811_));
 sky130_fd_sc_hd__mux4_2 _18297_ (.A0(_04807_),
    .A1(_04808_),
    .A2(_04810_),
    .A3(_04811_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04812_));
 sky130_fd_sc_hd__mux4_2 _18298_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04813_));
 sky130_fd_sc_hd__mux4_2 _18299_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04814_));
 sky130_fd_sc_hd__mux4_2 _18300_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04815_));
 sky130_fd_sc_hd__mux4_2 _18302_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04817_));
 sky130_fd_sc_hd__mux4_2 _18304_ (.A0(_04813_),
    .A1(_04814_),
    .A2(_04815_),
    .A3(_04817_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04819_));
 sky130_fd_sc_hd__mux2_2 _18306_ (.A0(_04812_),
    .A1(_04819_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[27] ));
 sky130_fd_sc_hd__mux4_2 _18307_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04821_));
 sky130_fd_sc_hd__mux4_2 _18308_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04822_));
 sky130_fd_sc_hd__mux4_2 _18309_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04823_));
 sky130_fd_sc_hd__mux4_2 _18310_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04824_));
 sky130_fd_sc_hd__mux4_2 _18311_ (.A0(_04821_),
    .A1(_04822_),
    .A2(_04823_),
    .A3(_04824_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04825_));
 sky130_fd_sc_hd__mux4_2 _18312_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04826_));
 sky130_fd_sc_hd__mux4_2 _18313_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04827_));
 sky130_fd_sc_hd__mux4_2 _18315_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04829_));
 sky130_fd_sc_hd__mux4_2 _18316_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04830_));
 sky130_fd_sc_hd__mux4_2 _18317_ (.A0(_04826_),
    .A1(_04827_),
    .A2(_04829_),
    .A3(_04830_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04831_));
 sky130_fd_sc_hd__mux2_2 _18318_ (.A0(_04825_),
    .A1(_04831_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[28] ));
 sky130_fd_sc_hd__mux4_2 _18319_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04832_));
 sky130_fd_sc_hd__mux4_2 _18320_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04833_));
 sky130_fd_sc_hd__mux4_2 _18321_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04834_));
 sky130_fd_sc_hd__mux4_2 _18322_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04835_));
 sky130_fd_sc_hd__mux4_2 _18323_ (.A0(_04832_),
    .A1(_04833_),
    .A2(_04834_),
    .A3(_04835_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04836_));
 sky130_fd_sc_hd__mux4_2 _18324_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04837_));
 sky130_fd_sc_hd__mux4_2 _18325_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04838_));
 sky130_fd_sc_hd__mux4_2 _18327_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04840_));
 sky130_fd_sc_hd__mux4_2 _18328_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04841_));
 sky130_fd_sc_hd__mux4_2 _18329_ (.A0(_04837_),
    .A1(_04838_),
    .A2(_04840_),
    .A3(_04841_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04842_));
 sky130_fd_sc_hd__mux2_2 _18330_ (.A0(_04836_),
    .A1(_04842_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[29] ));
 sky130_fd_sc_hd__mux4_2 _18332_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04844_));
 sky130_fd_sc_hd__mux4_2 _18333_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04845_));
 sky130_fd_sc_hd__mux4_2 _18334_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04846_));
 sky130_fd_sc_hd__mux4_2 _18335_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04847_));
 sky130_fd_sc_hd__mux4_2 _18336_ (.A0(_04844_),
    .A1(_04845_),
    .A2(_04846_),
    .A3(_04847_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04848_));
 sky130_fd_sc_hd__mux4_2 _18337_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04849_));
 sky130_fd_sc_hd__mux4_2 _18338_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04850_));
 sky130_fd_sc_hd__mux4_2 _18339_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04851_));
 sky130_fd_sc_hd__mux4_2 _18340_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04852_));
 sky130_fd_sc_hd__mux4_2 _18341_ (.A0(_04849_),
    .A1(_04850_),
    .A2(_04851_),
    .A3(_04852_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04853_));
 sky130_fd_sc_hd__mux2_2 _18342_ (.A0(_04848_),
    .A1(_04853_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[2] ));
 sky130_fd_sc_hd__mux4_2 _18343_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04854_));
 sky130_fd_sc_hd__mux4_2 _18344_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04855_));
 sky130_fd_sc_hd__mux4_2 _18345_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04856_));
 sky130_fd_sc_hd__mux4_2 _18346_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04857_));
 sky130_fd_sc_hd__mux4_2 _18347_ (.A0(_04854_),
    .A1(_04855_),
    .A2(_04856_),
    .A3(_04857_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04858_));
 sky130_fd_sc_hd__mux4_2 _18348_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04859_));
 sky130_fd_sc_hd__mux4_2 _18349_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04860_));
 sky130_fd_sc_hd__mux4_2 _18350_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04861_));
 sky130_fd_sc_hd__mux4_2 _18351_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04862_));
 sky130_fd_sc_hd__mux4_2 _18352_ (.A0(_04859_),
    .A1(_04860_),
    .A2(_04861_),
    .A3(_04862_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04863_));
 sky130_fd_sc_hd__mux2_2 _18353_ (.A0(_04858_),
    .A1(_04863_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[30] ));
 sky130_fd_sc_hd__mux4_2 _18354_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04864_));
 sky130_fd_sc_hd__mux4_2 _18355_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04865_));
 sky130_fd_sc_hd__mux4_2 _18356_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04866_));
 sky130_fd_sc_hd__mux4_2 _18357_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04867_));
 sky130_fd_sc_hd__mux4_2 _18358_ (.A0(_04864_),
    .A1(_04865_),
    .A2(_04866_),
    .A3(_04867_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04868_));
 sky130_fd_sc_hd__mux4_2 _18359_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04869_));
 sky130_fd_sc_hd__mux4_2 _18360_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04870_));
 sky130_fd_sc_hd__mux4_2 _18361_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04871_));
 sky130_fd_sc_hd__mux4_2 _18362_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04872_));
 sky130_fd_sc_hd__mux4_2 _18363_ (.A0(_04869_),
    .A1(_04870_),
    .A2(_04871_),
    .A3(_04872_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04873_));
 sky130_fd_sc_hd__mux2_2 _18364_ (.A0(_04868_),
    .A1(_04873_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[31] ));
 sky130_fd_sc_hd__mux4_2 _18365_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04874_));
 sky130_fd_sc_hd__mux4_2 _18366_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04875_));
 sky130_fd_sc_hd__mux4_2 _18367_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04876_));
 sky130_fd_sc_hd__mux4_2 _18368_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04877_));
 sky130_fd_sc_hd__mux4_2 _18369_ (.A0(_04874_),
    .A1(_04875_),
    .A2(_04876_),
    .A3(_04877_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04878_));
 sky130_fd_sc_hd__mux4_2 _18370_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04879_));
 sky130_fd_sc_hd__mux4_2 _18371_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04880_));
 sky130_fd_sc_hd__mux4_2 _18372_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04881_));
 sky130_fd_sc_hd__mux4_2 _18373_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04882_));
 sky130_fd_sc_hd__mux4_2 _18374_ (.A0(_04879_),
    .A1(_04880_),
    .A2(_04881_),
    .A3(_04882_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04883_));
 sky130_fd_sc_hd__mux2_2 _18375_ (.A0(_04878_),
    .A1(_04883_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[3] ));
 sky130_fd_sc_hd__mux4_2 _18376_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04884_));
 sky130_fd_sc_hd__mux4_2 _18377_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04885_));
 sky130_fd_sc_hd__mux4_2 _18378_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04886_));
 sky130_fd_sc_hd__mux4_2 _18379_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04887_));
 sky130_fd_sc_hd__mux4_2 _18380_ (.A0(_04884_),
    .A1(_04885_),
    .A2(_04886_),
    .A3(_04887_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04888_));
 sky130_fd_sc_hd__mux4_2 _18381_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04889_));
 sky130_fd_sc_hd__mux4_2 _18382_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04890_));
 sky130_fd_sc_hd__mux4_2 _18383_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04891_));
 sky130_fd_sc_hd__mux4_2 _18384_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04892_));
 sky130_fd_sc_hd__mux4_2 _18385_ (.A0(_04889_),
    .A1(_04890_),
    .A2(_04891_),
    .A3(_04892_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04893_));
 sky130_fd_sc_hd__mux2_2 _18386_ (.A0(_04888_),
    .A1(_04893_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[4] ));
 sky130_fd_sc_hd__mux4_2 _18387_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04894_));
 sky130_fd_sc_hd__mux4_2 _18388_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04895_));
 sky130_fd_sc_hd__mux4_2 _18389_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04896_));
 sky130_fd_sc_hd__mux4_2 _18390_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04897_));
 sky130_fd_sc_hd__mux4_2 _18391_ (.A0(_04894_),
    .A1(_04895_),
    .A2(_04896_),
    .A3(_04897_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04898_));
 sky130_fd_sc_hd__mux4_2 _18392_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04899_));
 sky130_fd_sc_hd__mux4_2 _18393_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04900_));
 sky130_fd_sc_hd__mux4_2 _18394_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04901_));
 sky130_fd_sc_hd__mux4_2 _18395_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04902_));
 sky130_fd_sc_hd__mux4_2 _18396_ (.A0(_04899_),
    .A1(_04900_),
    .A2(_04901_),
    .A3(_04902_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04903_));
 sky130_fd_sc_hd__mux2_2 _18397_ (.A0(_04898_),
    .A1(_04903_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[5] ));
 sky130_fd_sc_hd__mux4_2 _18398_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04904_));
 sky130_fd_sc_hd__mux4_2 _18399_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04905_));
 sky130_fd_sc_hd__mux4_2 _18400_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04906_));
 sky130_fd_sc_hd__mux4_2 _18401_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04907_));
 sky130_fd_sc_hd__mux4_2 _18402_ (.A0(_04904_),
    .A1(_04905_),
    .A2(_04906_),
    .A3(_04907_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04908_));
 sky130_fd_sc_hd__mux4_2 _18403_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04909_));
 sky130_fd_sc_hd__mux4_2 _18404_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04910_));
 sky130_fd_sc_hd__mux4_2 _18405_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04911_));
 sky130_fd_sc_hd__mux4_2 _18406_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04912_));
 sky130_fd_sc_hd__mux4_2 _18407_ (.A0(_04909_),
    .A1(_04910_),
    .A2(_04911_),
    .A3(_04912_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04913_));
 sky130_fd_sc_hd__mux2_2 _18408_ (.A0(_04908_),
    .A1(_04913_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[6] ));
 sky130_fd_sc_hd__mux4_2 _18409_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04914_));
 sky130_fd_sc_hd__mux4_2 _18410_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04915_));
 sky130_fd_sc_hd__mux4_2 _18411_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04916_));
 sky130_fd_sc_hd__mux4_2 _18412_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04917_));
 sky130_fd_sc_hd__mux4_2 _18413_ (.A0(_04914_),
    .A1(_04915_),
    .A2(_04916_),
    .A3(_04917_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04918_));
 sky130_fd_sc_hd__mux4_2 _18414_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04919_));
 sky130_fd_sc_hd__mux4_2 _18415_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04920_));
 sky130_fd_sc_hd__mux4_2 _18416_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04921_));
 sky130_fd_sc_hd__mux4_2 _18417_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04922_));
 sky130_fd_sc_hd__mux4_2 _18418_ (.A0(_04919_),
    .A1(_04920_),
    .A2(_04921_),
    .A3(_04922_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04923_));
 sky130_fd_sc_hd__mux2_2 _18419_ (.A0(_04918_),
    .A1(_04923_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[7] ));
 sky130_fd_sc_hd__mux4_2 _18420_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04924_));
 sky130_fd_sc_hd__mux4_2 _18421_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04925_));
 sky130_fd_sc_hd__mux4_2 _18422_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04926_));
 sky130_fd_sc_hd__mux4_2 _18423_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04927_));
 sky130_fd_sc_hd__mux4_2 _18424_ (.A0(_04924_),
    .A1(_04925_),
    .A2(_04926_),
    .A3(_04927_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04928_));
 sky130_fd_sc_hd__mux4_2 _18425_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04929_));
 sky130_fd_sc_hd__mux4_2 _18426_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04930_));
 sky130_fd_sc_hd__mux4_2 _18427_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04931_));
 sky130_fd_sc_hd__mux4_2 _18428_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04932_));
 sky130_fd_sc_hd__mux4_2 _18429_ (.A0(_04929_),
    .A1(_04930_),
    .A2(_04931_),
    .A3(_04932_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04933_));
 sky130_fd_sc_hd__mux2_2 _18430_ (.A0(_04928_),
    .A1(_04933_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[8] ));
 sky130_fd_sc_hd__mux4_2 _18431_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04934_));
 sky130_fd_sc_hd__mux4_2 _18432_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04935_));
 sky130_fd_sc_hd__mux4_2 _18433_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04936_));
 sky130_fd_sc_hd__mux4_2 _18434_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04937_));
 sky130_fd_sc_hd__mux4_2 _18435_ (.A0(_04934_),
    .A1(_04935_),
    .A2(_04936_),
    .A3(_04937_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04938_));
 sky130_fd_sc_hd__mux4_2 _18436_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04939_));
 sky130_fd_sc_hd__mux4_2 _18437_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04940_));
 sky130_fd_sc_hd__mux4_2 _18438_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04941_));
 sky130_fd_sc_hd__mux4_2 _18439_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_04942_));
 sky130_fd_sc_hd__mux4_2 _18440_ (.A0(_04939_),
    .A1(_04940_),
    .A2(_04941_),
    .A3(_04942_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[5] ),
    .X(_04943_));
 sky130_fd_sc_hd__mux2_2 _18441_ (.A0(_04938_),
    .A1(_04943_),
    .S(\count15_2[4] ),
    .X(\w_new_calc2.w_15[9] ));
 sky130_fd_sc_hd__mux4_2 _18446_ (.A0(\w[1][0] ),
    .A1(\w[3][0] ),
    .A2(\w[5][0] ),
    .A3(\w[7][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04948_));
 sky130_fd_sc_hd__mux4_2 _18450_ (.A0(\w[9][0] ),
    .A1(\w[11][0] ),
    .A2(\w[13][0] ),
    .A3(\w[15][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04952_));
 sky130_fd_sc_hd__mux4_2 _18454_ (.A0(\w[33][0] ),
    .A1(\w[35][0] ),
    .A2(\w[37][0] ),
    .A3(\w[39][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04956_));
 sky130_fd_sc_hd__mux4_2 _18457_ (.A0(\w[41][0] ),
    .A1(\w[43][0] ),
    .A2(\w[45][0] ),
    .A3(\w[47][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04959_));
 sky130_fd_sc_hd__mux4_2 _18461_ (.A0(_04948_),
    .A1(_04952_),
    .A2(_04956_),
    .A3(_04959_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_04963_));
 sky130_fd_sc_hd__mux4_2 _18464_ (.A0(\w[17][0] ),
    .A1(\w[19][0] ),
    .A2(\w[21][0] ),
    .A3(\w[23][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04966_));
 sky130_fd_sc_hd__mux4_2 _18467_ (.A0(\w[25][0] ),
    .A1(\w[27][0] ),
    .A2(\w[29][0] ),
    .A3(\w[31][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04969_));
 sky130_fd_sc_hd__mux4_2 _18470_ (.A0(\w[49][0] ),
    .A1(\w[51][0] ),
    .A2(\w[53][0] ),
    .A3(\w[55][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04972_));
 sky130_fd_sc_hd__mux4_2 _18471_ (.A0(\w[57][0] ),
    .A1(\w[59][0] ),
    .A2(\w[61][0] ),
    .A3(\w[63][0] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04973_));
 sky130_fd_sc_hd__mux4_2 _18472_ (.A0(_04966_),
    .A1(_04969_),
    .A2(_04972_),
    .A3(_04973_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_04974_));
 sky130_fd_sc_hd__mux2_2 _18473_ (.A0(_04963_),
    .A1(_04974_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[0] ));
 sky130_fd_sc_hd__mux4_2 _18474_ (.A0(\w[1][10] ),
    .A1(\w[3][10] ),
    .A2(\w[5][10] ),
    .A3(\w[7][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04975_));
 sky130_fd_sc_hd__mux4_2 _18475_ (.A0(\w[9][10] ),
    .A1(\w[11][10] ),
    .A2(\w[13][10] ),
    .A3(\w[15][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04976_));
 sky130_fd_sc_hd__mux4_2 _18476_ (.A0(\w[33][10] ),
    .A1(\w[35][10] ),
    .A2(\w[37][10] ),
    .A3(\w[39][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04977_));
 sky130_fd_sc_hd__mux4_2 _18477_ (.A0(\w[41][10] ),
    .A1(\w[43][10] ),
    .A2(\w[45][10] ),
    .A3(\w[47][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04978_));
 sky130_fd_sc_hd__mux4_2 _18478_ (.A0(_04975_),
    .A1(_04976_),
    .A2(_04977_),
    .A3(_04978_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_04979_));
 sky130_fd_sc_hd__mux4_2 _18479_ (.A0(\w[17][10] ),
    .A1(\w[19][10] ),
    .A2(\w[21][10] ),
    .A3(\w[23][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04980_));
 sky130_fd_sc_hd__mux4_2 _18480_ (.A0(\w[25][10] ),
    .A1(\w[27][10] ),
    .A2(\w[29][10] ),
    .A3(\w[31][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04981_));
 sky130_fd_sc_hd__mux4_2 _18482_ (.A0(\w[49][10] ),
    .A1(\w[51][10] ),
    .A2(\w[53][10] ),
    .A3(\w[55][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04983_));
 sky130_fd_sc_hd__mux4_2 _18483_ (.A0(\w[57][10] ),
    .A1(\w[59][10] ),
    .A2(\w[61][10] ),
    .A3(\w[63][10] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04984_));
 sky130_fd_sc_hd__mux4_2 _18484_ (.A0(_04980_),
    .A1(_04981_),
    .A2(_04983_),
    .A3(_04984_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_04985_));
 sky130_fd_sc_hd__mux2_2 _18485_ (.A0(_04979_),
    .A1(_04985_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[10] ));
 sky130_fd_sc_hd__mux4_2 _18487_ (.A0(\w[1][11] ),
    .A1(\w[3][11] ),
    .A2(\w[5][11] ),
    .A3(\w[7][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04987_));
 sky130_fd_sc_hd__mux4_2 _18488_ (.A0(\w[9][11] ),
    .A1(\w[11][11] ),
    .A2(\w[13][11] ),
    .A3(\w[15][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04988_));
 sky130_fd_sc_hd__mux4_2 _18489_ (.A0(\w[33][11] ),
    .A1(\w[35][11] ),
    .A2(\w[37][11] ),
    .A3(\w[39][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04989_));
 sky130_fd_sc_hd__mux4_2 _18490_ (.A0(\w[41][11] ),
    .A1(\w[43][11] ),
    .A2(\w[45][11] ),
    .A3(\w[47][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04990_));
 sky130_fd_sc_hd__mux4_2 _18491_ (.A0(_04987_),
    .A1(_04988_),
    .A2(_04989_),
    .A3(_04990_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_04991_));
 sky130_fd_sc_hd__mux4_2 _18492_ (.A0(\w[17][11] ),
    .A1(\w[19][11] ),
    .A2(\w[21][11] ),
    .A3(\w[23][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04992_));
 sky130_fd_sc_hd__mux4_2 _18493_ (.A0(\w[25][11] ),
    .A1(\w[27][11] ),
    .A2(\w[29][11] ),
    .A3(\w[31][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04993_));
 sky130_fd_sc_hd__mux4_2 _18494_ (.A0(\w[49][11] ),
    .A1(\w[51][11] ),
    .A2(\w[53][11] ),
    .A3(\w[55][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04994_));
 sky130_fd_sc_hd__mux4_2 _18495_ (.A0(\w[57][11] ),
    .A1(\w[59][11] ),
    .A2(\w[61][11] ),
    .A3(\w[63][11] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04995_));
 sky130_fd_sc_hd__mux4_2 _18496_ (.A0(_04992_),
    .A1(_04993_),
    .A2(_04994_),
    .A3(_04995_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_04996_));
 sky130_fd_sc_hd__mux2_2 _18497_ (.A0(_04991_),
    .A1(_04996_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[11] ));
 sky130_fd_sc_hd__mux4_2 _18499_ (.A0(\w[1][12] ),
    .A1(\w[3][12] ),
    .A2(\w[5][12] ),
    .A3(\w[7][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04998_));
 sky130_fd_sc_hd__mux4_2 _18500_ (.A0(\w[9][12] ),
    .A1(\w[11][12] ),
    .A2(\w[13][12] ),
    .A3(\w[15][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_04999_));
 sky130_fd_sc_hd__mux4_2 _18501_ (.A0(\w[33][12] ),
    .A1(\w[35][12] ),
    .A2(\w[37][12] ),
    .A3(\w[39][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05000_));
 sky130_fd_sc_hd__mux4_2 _18502_ (.A0(\w[41][12] ),
    .A1(\w[43][12] ),
    .A2(\w[45][12] ),
    .A3(\w[47][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05001_));
 sky130_fd_sc_hd__mux4_2 _18503_ (.A0(_04998_),
    .A1(_04999_),
    .A2(_05000_),
    .A3(_05001_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05002_));
 sky130_fd_sc_hd__mux4_2 _18504_ (.A0(\w[17][12] ),
    .A1(\w[19][12] ),
    .A2(\w[21][12] ),
    .A3(\w[23][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05003_));
 sky130_fd_sc_hd__mux4_2 _18505_ (.A0(\w[25][12] ),
    .A1(\w[27][12] ),
    .A2(\w[29][12] ),
    .A3(\w[31][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05004_));
 sky130_fd_sc_hd__mux4_2 _18506_ (.A0(\w[49][12] ),
    .A1(\w[51][12] ),
    .A2(\w[53][12] ),
    .A3(\w[55][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05005_));
 sky130_fd_sc_hd__mux4_2 _18507_ (.A0(\w[57][12] ),
    .A1(\w[59][12] ),
    .A2(\w[61][12] ),
    .A3(\w[63][12] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05006_));
 sky130_fd_sc_hd__mux4_2 _18508_ (.A0(_05003_),
    .A1(_05004_),
    .A2(_05005_),
    .A3(_05006_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_2 _18509_ (.A0(_05002_),
    .A1(_05007_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[12] ));
 sky130_fd_sc_hd__mux4_2 _18510_ (.A0(\w[1][13] ),
    .A1(\w[3][13] ),
    .A2(\w[5][13] ),
    .A3(\w[7][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05008_));
 sky130_fd_sc_hd__mux4_2 _18512_ (.A0(\w[9][13] ),
    .A1(\w[11][13] ),
    .A2(\w[13][13] ),
    .A3(\w[15][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05010_));
 sky130_fd_sc_hd__mux4_2 _18513_ (.A0(\w[33][13] ),
    .A1(\w[35][13] ),
    .A2(\w[37][13] ),
    .A3(\w[39][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05011_));
 sky130_fd_sc_hd__mux4_2 _18514_ (.A0(\w[41][13] ),
    .A1(\w[43][13] ),
    .A2(\w[45][13] ),
    .A3(\w[47][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05012_));
 sky130_fd_sc_hd__mux4_2 _18515_ (.A0(_05008_),
    .A1(_05010_),
    .A2(_05011_),
    .A3(_05012_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05013_));
 sky130_fd_sc_hd__mux4_2 _18517_ (.A0(\w[17][13] ),
    .A1(\w[19][13] ),
    .A2(\w[21][13] ),
    .A3(\w[23][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05015_));
 sky130_fd_sc_hd__mux4_2 _18518_ (.A0(\w[25][13] ),
    .A1(\w[27][13] ),
    .A2(\w[29][13] ),
    .A3(\w[31][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05016_));
 sky130_fd_sc_hd__mux4_2 _18519_ (.A0(\w[49][13] ),
    .A1(\w[51][13] ),
    .A2(\w[53][13] ),
    .A3(\w[55][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05017_));
 sky130_fd_sc_hd__mux4_2 _18520_ (.A0(\w[57][13] ),
    .A1(\w[59][13] ),
    .A2(\w[61][13] ),
    .A3(\w[63][13] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05018_));
 sky130_fd_sc_hd__mux4_2 _18521_ (.A0(_05015_),
    .A1(_05016_),
    .A2(_05017_),
    .A3(_05018_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05019_));
 sky130_fd_sc_hd__mux2_2 _18522_ (.A0(_05013_),
    .A1(_05019_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[13] ));
 sky130_fd_sc_hd__mux4_2 _18523_ (.A0(\w[1][14] ),
    .A1(\w[3][14] ),
    .A2(\w[5][14] ),
    .A3(\w[7][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05020_));
 sky130_fd_sc_hd__mux4_2 _18525_ (.A0(\w[9][14] ),
    .A1(\w[11][14] ),
    .A2(\w[13][14] ),
    .A3(\w[15][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05022_));
 sky130_fd_sc_hd__mux4_2 _18526_ (.A0(\w[33][14] ),
    .A1(\w[35][14] ),
    .A2(\w[37][14] ),
    .A3(\w[39][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05023_));
 sky130_fd_sc_hd__mux4_2 _18527_ (.A0(\w[41][14] ),
    .A1(\w[43][14] ),
    .A2(\w[45][14] ),
    .A3(\w[47][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05024_));
 sky130_fd_sc_hd__mux4_2 _18529_ (.A0(_05020_),
    .A1(_05022_),
    .A2(_05023_),
    .A3(_05024_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05026_));
 sky130_fd_sc_hd__mux4_2 _18531_ (.A0(\w[17][14] ),
    .A1(\w[19][14] ),
    .A2(\w[21][14] ),
    .A3(\w[23][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05028_));
 sky130_fd_sc_hd__mux4_2 _18532_ (.A0(\w[25][14] ),
    .A1(\w[27][14] ),
    .A2(\w[29][14] ),
    .A3(\w[31][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05029_));
 sky130_fd_sc_hd__mux4_2 _18533_ (.A0(\w[49][14] ),
    .A1(\w[51][14] ),
    .A2(\w[53][14] ),
    .A3(\w[55][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05030_));
 sky130_fd_sc_hd__mux4_2 _18534_ (.A0(\w[57][14] ),
    .A1(\w[59][14] ),
    .A2(\w[61][14] ),
    .A3(\w[63][14] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05031_));
 sky130_fd_sc_hd__mux4_2 _18535_ (.A0(_05028_),
    .A1(_05029_),
    .A2(_05030_),
    .A3(_05031_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05032_));
 sky130_fd_sc_hd__mux2_2 _18536_ (.A0(_05026_),
    .A1(_05032_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[14] ));
 sky130_fd_sc_hd__mux4_2 _18537_ (.A0(\w[1][15] ),
    .A1(\w[3][15] ),
    .A2(\w[5][15] ),
    .A3(\w[7][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05033_));
 sky130_fd_sc_hd__mux4_2 _18538_ (.A0(\w[9][15] ),
    .A1(\w[11][15] ),
    .A2(\w[13][15] ),
    .A3(\w[15][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05034_));
 sky130_fd_sc_hd__mux4_2 _18539_ (.A0(\w[33][15] ),
    .A1(\w[35][15] ),
    .A2(\w[37][15] ),
    .A3(\w[39][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05035_));
 sky130_fd_sc_hd__mux4_2 _18541_ (.A0(\w[41][15] ),
    .A1(\w[43][15] ),
    .A2(\w[45][15] ),
    .A3(\w[47][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05037_));
 sky130_fd_sc_hd__mux4_2 _18542_ (.A0(_05033_),
    .A1(_05034_),
    .A2(_05035_),
    .A3(_05037_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05038_));
 sky130_fd_sc_hd__mux4_2 _18543_ (.A0(\w[17][15] ),
    .A1(\w[19][15] ),
    .A2(\w[21][15] ),
    .A3(\w[23][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05039_));
 sky130_fd_sc_hd__mux4_2 _18545_ (.A0(\w[25][15] ),
    .A1(\w[27][15] ),
    .A2(\w[29][15] ),
    .A3(\w[31][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05041_));
 sky130_fd_sc_hd__mux4_2 _18546_ (.A0(\w[49][15] ),
    .A1(\w[51][15] ),
    .A2(\w[53][15] ),
    .A3(\w[55][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05042_));
 sky130_fd_sc_hd__mux4_2 _18547_ (.A0(\w[57][15] ),
    .A1(\w[59][15] ),
    .A2(\w[61][15] ),
    .A3(\w[63][15] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05043_));
 sky130_fd_sc_hd__mux4_2 _18548_ (.A0(_05039_),
    .A1(_05041_),
    .A2(_05042_),
    .A3(_05043_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05044_));
 sky130_fd_sc_hd__mux2_2 _18549_ (.A0(_05038_),
    .A1(_05044_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[15] ));
 sky130_fd_sc_hd__mux4_2 _18550_ (.A0(\w[1][16] ),
    .A1(\w[3][16] ),
    .A2(\w[5][16] ),
    .A3(\w[7][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05045_));
 sky130_fd_sc_hd__mux4_2 _18551_ (.A0(\w[9][16] ),
    .A1(\w[11][16] ),
    .A2(\w[13][16] ),
    .A3(\w[15][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05046_));
 sky130_fd_sc_hd__mux4_2 _18552_ (.A0(\w[33][16] ),
    .A1(\w[35][16] ),
    .A2(\w[37][16] ),
    .A3(\w[39][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05047_));
 sky130_fd_sc_hd__mux4_2 _18554_ (.A0(\w[41][16] ),
    .A1(\w[43][16] ),
    .A2(\w[45][16] ),
    .A3(\w[47][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05049_));
 sky130_fd_sc_hd__mux4_2 _18556_ (.A0(_05045_),
    .A1(_05046_),
    .A2(_05047_),
    .A3(_05049_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05051_));
 sky130_fd_sc_hd__mux4_2 _18557_ (.A0(\w[17][16] ),
    .A1(\w[19][16] ),
    .A2(\w[21][16] ),
    .A3(\w[23][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05052_));
 sky130_fd_sc_hd__mux4_2 _18559_ (.A0(\w[25][16] ),
    .A1(\w[27][16] ),
    .A2(\w[29][16] ),
    .A3(\w[31][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05054_));
 sky130_fd_sc_hd__mux4_2 _18560_ (.A0(\w[49][16] ),
    .A1(\w[51][16] ),
    .A2(\w[53][16] ),
    .A3(\w[55][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05055_));
 sky130_fd_sc_hd__mux4_2 _18561_ (.A0(\w[57][16] ),
    .A1(\w[59][16] ),
    .A2(\w[61][16] ),
    .A3(\w[63][16] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05056_));
 sky130_fd_sc_hd__mux4_2 _18563_ (.A0(_05052_),
    .A1(_05054_),
    .A2(_05055_),
    .A3(_05056_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05058_));
 sky130_fd_sc_hd__mux2_2 _18564_ (.A0(_05051_),
    .A1(_05058_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[16] ));
 sky130_fd_sc_hd__mux4_2 _18565_ (.A0(\w[1][17] ),
    .A1(\w[3][17] ),
    .A2(\w[5][17] ),
    .A3(\w[7][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05059_));
 sky130_fd_sc_hd__mux4_2 _18566_ (.A0(\w[9][17] ),
    .A1(\w[11][17] ),
    .A2(\w[13][17] ),
    .A3(\w[15][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05060_));
 sky130_fd_sc_hd__mux4_2 _18568_ (.A0(\w[33][17] ),
    .A1(\w[35][17] ),
    .A2(\w[37][17] ),
    .A3(\w[39][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05062_));
 sky130_fd_sc_hd__mux4_2 _18569_ (.A0(\w[41][17] ),
    .A1(\w[43][17] ),
    .A2(\w[45][17] ),
    .A3(\w[47][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05063_));
 sky130_fd_sc_hd__mux4_2 _18570_ (.A0(_05059_),
    .A1(_05060_),
    .A2(_05062_),
    .A3(_05063_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05064_));
 sky130_fd_sc_hd__mux4_2 _18571_ (.A0(\w[17][17] ),
    .A1(\w[19][17] ),
    .A2(\w[21][17] ),
    .A3(\w[23][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05065_));
 sky130_fd_sc_hd__mux4_2 _18572_ (.A0(\w[25][17] ),
    .A1(\w[27][17] ),
    .A2(\w[29][17] ),
    .A3(\w[31][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05066_));
 sky130_fd_sc_hd__mux4_2 _18573_ (.A0(\w[49][17] ),
    .A1(\w[51][17] ),
    .A2(\w[53][17] ),
    .A3(\w[55][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05067_));
 sky130_fd_sc_hd__mux4_2 _18575_ (.A0(\w[57][17] ),
    .A1(\w[59][17] ),
    .A2(\w[61][17] ),
    .A3(\w[63][17] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05069_));
 sky130_fd_sc_hd__mux4_2 _18576_ (.A0(_05065_),
    .A1(_05066_),
    .A2(_05067_),
    .A3(_05069_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05070_));
 sky130_fd_sc_hd__mux2_2 _18577_ (.A0(_05064_),
    .A1(_05070_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[17] ));
 sky130_fd_sc_hd__mux4_2 _18578_ (.A0(\w[1][18] ),
    .A1(\w[3][18] ),
    .A2(\w[5][18] ),
    .A3(\w[7][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05071_));
 sky130_fd_sc_hd__mux4_2 _18579_ (.A0(\w[9][18] ),
    .A1(\w[11][18] ),
    .A2(\w[13][18] ),
    .A3(\w[15][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05072_));
 sky130_fd_sc_hd__mux4_2 _18581_ (.A0(\w[33][18] ),
    .A1(\w[35][18] ),
    .A2(\w[37][18] ),
    .A3(\w[39][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05074_));
 sky130_fd_sc_hd__mux4_2 _18582_ (.A0(\w[41][18] ),
    .A1(\w[43][18] ),
    .A2(\w[45][18] ),
    .A3(\w[47][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05075_));
 sky130_fd_sc_hd__mux4_2 _18583_ (.A0(_05071_),
    .A1(_05072_),
    .A2(_05074_),
    .A3(_05075_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05076_));
 sky130_fd_sc_hd__mux4_2 _18584_ (.A0(\w[17][18] ),
    .A1(\w[19][18] ),
    .A2(\w[21][18] ),
    .A3(\w[23][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05077_));
 sky130_fd_sc_hd__mux4_2 _18585_ (.A0(\w[25][18] ),
    .A1(\w[27][18] ),
    .A2(\w[29][18] ),
    .A3(\w[31][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05078_));
 sky130_fd_sc_hd__mux4_2 _18586_ (.A0(\w[49][18] ),
    .A1(\w[51][18] ),
    .A2(\w[53][18] ),
    .A3(\w[55][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05079_));
 sky130_fd_sc_hd__mux4_2 _18588_ (.A0(\w[57][18] ),
    .A1(\w[59][18] ),
    .A2(\w[61][18] ),
    .A3(\w[63][18] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05081_));
 sky130_fd_sc_hd__mux4_2 _18590_ (.A0(_05077_),
    .A1(_05078_),
    .A2(_05079_),
    .A3(_05081_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05083_));
 sky130_fd_sc_hd__mux2_2 _18592_ (.A0(_05076_),
    .A1(_05083_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[18] ));
 sky130_fd_sc_hd__mux4_2 _18593_ (.A0(\w[1][19] ),
    .A1(\w[3][19] ),
    .A2(\w[5][19] ),
    .A3(\w[7][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05085_));
 sky130_fd_sc_hd__mux4_2 _18594_ (.A0(\w[9][19] ),
    .A1(\w[11][19] ),
    .A2(\w[13][19] ),
    .A3(\w[15][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05086_));
 sky130_fd_sc_hd__mux4_2 _18595_ (.A0(\w[33][19] ),
    .A1(\w[35][19] ),
    .A2(\w[37][19] ),
    .A3(\w[39][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05087_));
 sky130_fd_sc_hd__mux4_2 _18596_ (.A0(\w[41][19] ),
    .A1(\w[43][19] ),
    .A2(\w[45][19] ),
    .A3(\w[47][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05088_));
 sky130_fd_sc_hd__mux4_2 _18597_ (.A0(_05085_),
    .A1(_05086_),
    .A2(_05087_),
    .A3(_05088_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05089_));
 sky130_fd_sc_hd__mux4_2 _18598_ (.A0(\w[17][19] ),
    .A1(\w[19][19] ),
    .A2(\w[21][19] ),
    .A3(\w[23][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05090_));
 sky130_fd_sc_hd__mux4_2 _18599_ (.A0(\w[25][19] ),
    .A1(\w[27][19] ),
    .A2(\w[29][19] ),
    .A3(\w[31][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05091_));
 sky130_fd_sc_hd__mux4_2 _18601_ (.A0(\w[49][19] ),
    .A1(\w[51][19] ),
    .A2(\w[53][19] ),
    .A3(\w[55][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05093_));
 sky130_fd_sc_hd__mux4_2 _18602_ (.A0(\w[57][19] ),
    .A1(\w[59][19] ),
    .A2(\w[61][19] ),
    .A3(\w[63][19] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05094_));
 sky130_fd_sc_hd__mux4_2 _18603_ (.A0(_05090_),
    .A1(_05091_),
    .A2(_05093_),
    .A3(_05094_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05095_));
 sky130_fd_sc_hd__mux2_2 _18604_ (.A0(_05089_),
    .A1(_05095_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[19] ));
 sky130_fd_sc_hd__mux4_2 _18605_ (.A0(\w[1][1] ),
    .A1(\w[3][1] ),
    .A2(\w[5][1] ),
    .A3(\w[7][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05096_));
 sky130_fd_sc_hd__mux4_2 _18606_ (.A0(\w[9][1] ),
    .A1(\w[11][1] ),
    .A2(\w[13][1] ),
    .A3(\w[15][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05097_));
 sky130_fd_sc_hd__mux4_2 _18607_ (.A0(\w[33][1] ),
    .A1(\w[35][1] ),
    .A2(\w[37][1] ),
    .A3(\w[39][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05098_));
 sky130_fd_sc_hd__mux4_2 _18608_ (.A0(\w[41][1] ),
    .A1(\w[43][1] ),
    .A2(\w[45][1] ),
    .A3(\w[47][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05099_));
 sky130_fd_sc_hd__mux4_2 _18609_ (.A0(_05096_),
    .A1(_05097_),
    .A2(_05098_),
    .A3(_05099_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05100_));
 sky130_fd_sc_hd__mux4_2 _18610_ (.A0(\w[17][1] ),
    .A1(\w[19][1] ),
    .A2(\w[21][1] ),
    .A3(\w[23][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05101_));
 sky130_fd_sc_hd__mux4_2 _18611_ (.A0(\w[25][1] ),
    .A1(\w[27][1] ),
    .A2(\w[29][1] ),
    .A3(\w[31][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05102_));
 sky130_fd_sc_hd__mux4_2 _18613_ (.A0(\w[49][1] ),
    .A1(\w[51][1] ),
    .A2(\w[53][1] ),
    .A3(\w[55][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05104_));
 sky130_fd_sc_hd__mux4_2 _18614_ (.A0(\w[57][1] ),
    .A1(\w[59][1] ),
    .A2(\w[61][1] ),
    .A3(\w[63][1] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05105_));
 sky130_fd_sc_hd__mux4_2 _18615_ (.A0(_05101_),
    .A1(_05102_),
    .A2(_05104_),
    .A3(_05105_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05106_));
 sky130_fd_sc_hd__mux2_2 _18616_ (.A0(_05100_),
    .A1(_05106_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[1] ));
 sky130_fd_sc_hd__mux4_2 _18618_ (.A0(\w[1][20] ),
    .A1(\w[3][20] ),
    .A2(\w[5][20] ),
    .A3(\w[7][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05108_));
 sky130_fd_sc_hd__mux4_2 _18619_ (.A0(\w[9][20] ),
    .A1(\w[11][20] ),
    .A2(\w[13][20] ),
    .A3(\w[15][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05109_));
 sky130_fd_sc_hd__mux4_2 _18620_ (.A0(\w[33][20] ),
    .A1(\w[35][20] ),
    .A2(\w[37][20] ),
    .A3(\w[39][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05110_));
 sky130_fd_sc_hd__mux4_2 _18621_ (.A0(\w[41][20] ),
    .A1(\w[43][20] ),
    .A2(\w[45][20] ),
    .A3(\w[47][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05111_));
 sky130_fd_sc_hd__mux4_2 _18622_ (.A0(_05108_),
    .A1(_05109_),
    .A2(_05110_),
    .A3(_05111_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05112_));
 sky130_fd_sc_hd__mux4_2 _18623_ (.A0(\w[17][20] ),
    .A1(\w[19][20] ),
    .A2(\w[21][20] ),
    .A3(\w[23][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05113_));
 sky130_fd_sc_hd__mux4_2 _18624_ (.A0(\w[25][20] ),
    .A1(\w[27][20] ),
    .A2(\w[29][20] ),
    .A3(\w[31][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05114_));
 sky130_fd_sc_hd__mux4_2 _18625_ (.A0(\w[49][20] ),
    .A1(\w[51][20] ),
    .A2(\w[53][20] ),
    .A3(\w[55][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05115_));
 sky130_fd_sc_hd__mux4_2 _18626_ (.A0(\w[57][20] ),
    .A1(\w[59][20] ),
    .A2(\w[61][20] ),
    .A3(\w[63][20] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05116_));
 sky130_fd_sc_hd__mux4_2 _18627_ (.A0(_05113_),
    .A1(_05114_),
    .A2(_05115_),
    .A3(_05116_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05117_));
 sky130_fd_sc_hd__mux2_2 _18628_ (.A0(_05112_),
    .A1(_05117_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[20] ));
 sky130_fd_sc_hd__mux4_2 _18630_ (.A0(\w[1][21] ),
    .A1(\w[3][21] ),
    .A2(\w[5][21] ),
    .A3(\w[7][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05119_));
 sky130_fd_sc_hd__mux4_2 _18631_ (.A0(\w[9][21] ),
    .A1(\w[11][21] ),
    .A2(\w[13][21] ),
    .A3(\w[15][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05120_));
 sky130_fd_sc_hd__mux4_2 _18632_ (.A0(\w[33][21] ),
    .A1(\w[35][21] ),
    .A2(\w[37][21] ),
    .A3(\w[39][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05121_));
 sky130_fd_sc_hd__mux4_2 _18633_ (.A0(\w[41][21] ),
    .A1(\w[43][21] ),
    .A2(\w[45][21] ),
    .A3(\w[47][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05122_));
 sky130_fd_sc_hd__mux4_2 _18634_ (.A0(_05119_),
    .A1(_05120_),
    .A2(_05121_),
    .A3(_05122_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05123_));
 sky130_fd_sc_hd__mux4_2 _18635_ (.A0(\w[17][21] ),
    .A1(\w[19][21] ),
    .A2(\w[21][21] ),
    .A3(\w[23][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05124_));
 sky130_fd_sc_hd__mux4_2 _18636_ (.A0(\w[25][21] ),
    .A1(\w[27][21] ),
    .A2(\w[29][21] ),
    .A3(\w[31][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05125_));
 sky130_fd_sc_hd__mux4_2 _18637_ (.A0(\w[49][21] ),
    .A1(\w[51][21] ),
    .A2(\w[53][21] ),
    .A3(\w[55][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05126_));
 sky130_fd_sc_hd__mux4_2 _18638_ (.A0(\w[57][21] ),
    .A1(\w[59][21] ),
    .A2(\w[61][21] ),
    .A3(\w[63][21] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05127_));
 sky130_fd_sc_hd__mux4_2 _18639_ (.A0(_05124_),
    .A1(_05125_),
    .A2(_05126_),
    .A3(_05127_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05128_));
 sky130_fd_sc_hd__mux2_2 _18640_ (.A0(_05123_),
    .A1(_05128_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[21] ));
 sky130_fd_sc_hd__mux4_2 _18641_ (.A0(\w[1][22] ),
    .A1(\w[3][22] ),
    .A2(\w[5][22] ),
    .A3(\w[7][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05129_));
 sky130_fd_sc_hd__mux4_2 _18643_ (.A0(\w[9][22] ),
    .A1(\w[11][22] ),
    .A2(\w[13][22] ),
    .A3(\w[15][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05131_));
 sky130_fd_sc_hd__mux4_2 _18644_ (.A0(\w[33][22] ),
    .A1(\w[35][22] ),
    .A2(\w[37][22] ),
    .A3(\w[39][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05132_));
 sky130_fd_sc_hd__mux4_2 _18645_ (.A0(\w[41][22] ),
    .A1(\w[43][22] ),
    .A2(\w[45][22] ),
    .A3(\w[47][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05133_));
 sky130_fd_sc_hd__mux4_2 _18646_ (.A0(_05129_),
    .A1(_05131_),
    .A2(_05132_),
    .A3(_05133_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05134_));
 sky130_fd_sc_hd__mux4_2 _18648_ (.A0(\w[17][22] ),
    .A1(\w[19][22] ),
    .A2(\w[21][22] ),
    .A3(\w[23][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05136_));
 sky130_fd_sc_hd__mux4_2 _18649_ (.A0(\w[25][22] ),
    .A1(\w[27][22] ),
    .A2(\w[29][22] ),
    .A3(\w[31][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05137_));
 sky130_fd_sc_hd__mux4_2 _18650_ (.A0(\w[49][22] ),
    .A1(\w[51][22] ),
    .A2(\w[53][22] ),
    .A3(\w[55][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05138_));
 sky130_fd_sc_hd__mux4_2 _18651_ (.A0(\w[57][22] ),
    .A1(\w[59][22] ),
    .A2(\w[61][22] ),
    .A3(\w[63][22] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05139_));
 sky130_fd_sc_hd__mux4_2 _18652_ (.A0(_05136_),
    .A1(_05137_),
    .A2(_05138_),
    .A3(_05139_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05140_));
 sky130_fd_sc_hd__mux2_2 _18653_ (.A0(_05134_),
    .A1(_05140_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[22] ));
 sky130_fd_sc_hd__mux4_2 _18654_ (.A0(\w[1][23] ),
    .A1(\w[3][23] ),
    .A2(\w[5][23] ),
    .A3(\w[7][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05141_));
 sky130_fd_sc_hd__mux4_2 _18656_ (.A0(\w[9][23] ),
    .A1(\w[11][23] ),
    .A2(\w[13][23] ),
    .A3(\w[15][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05143_));
 sky130_fd_sc_hd__mux4_2 _18657_ (.A0(\w[33][23] ),
    .A1(\w[35][23] ),
    .A2(\w[37][23] ),
    .A3(\w[39][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05144_));
 sky130_fd_sc_hd__mux4_2 _18658_ (.A0(\w[41][23] ),
    .A1(\w[43][23] ),
    .A2(\w[45][23] ),
    .A3(\w[47][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05145_));
 sky130_fd_sc_hd__mux4_2 _18660_ (.A0(_05141_),
    .A1(_05143_),
    .A2(_05144_),
    .A3(_05145_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05147_));
 sky130_fd_sc_hd__mux4_2 _18662_ (.A0(\w[17][23] ),
    .A1(\w[19][23] ),
    .A2(\w[21][23] ),
    .A3(\w[23][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05149_));
 sky130_fd_sc_hd__mux4_2 _18663_ (.A0(\w[25][23] ),
    .A1(\w[27][23] ),
    .A2(\w[29][23] ),
    .A3(\w[31][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05150_));
 sky130_fd_sc_hd__mux4_2 _18664_ (.A0(\w[49][23] ),
    .A1(\w[51][23] ),
    .A2(\w[53][23] ),
    .A3(\w[55][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05151_));
 sky130_fd_sc_hd__mux4_2 _18665_ (.A0(\w[57][23] ),
    .A1(\w[59][23] ),
    .A2(\w[61][23] ),
    .A3(\w[63][23] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05152_));
 sky130_fd_sc_hd__mux4_2 _18666_ (.A0(_05149_),
    .A1(_05150_),
    .A2(_05151_),
    .A3(_05152_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05153_));
 sky130_fd_sc_hd__mux2_2 _18667_ (.A0(_05147_),
    .A1(_05153_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[23] ));
 sky130_fd_sc_hd__mux4_2 _18668_ (.A0(\w[1][24] ),
    .A1(\w[3][24] ),
    .A2(\w[5][24] ),
    .A3(\w[7][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05154_));
 sky130_fd_sc_hd__mux4_2 _18669_ (.A0(\w[9][24] ),
    .A1(\w[11][24] ),
    .A2(\w[13][24] ),
    .A3(\w[15][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05155_));
 sky130_fd_sc_hd__mux4_2 _18670_ (.A0(\w[33][24] ),
    .A1(\w[35][24] ),
    .A2(\w[37][24] ),
    .A3(\w[39][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05156_));
 sky130_fd_sc_hd__mux4_2 _18672_ (.A0(\w[41][24] ),
    .A1(\w[43][24] ),
    .A2(\w[45][24] ),
    .A3(\w[47][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05158_));
 sky130_fd_sc_hd__mux4_2 _18673_ (.A0(_05154_),
    .A1(_05155_),
    .A2(_05156_),
    .A3(_05158_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05159_));
 sky130_fd_sc_hd__mux4_2 _18674_ (.A0(\w[17][24] ),
    .A1(\w[19][24] ),
    .A2(\w[21][24] ),
    .A3(\w[23][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05160_));
 sky130_fd_sc_hd__mux4_2 _18676_ (.A0(\w[25][24] ),
    .A1(\w[27][24] ),
    .A2(\w[29][24] ),
    .A3(\w[31][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05162_));
 sky130_fd_sc_hd__mux4_2 _18677_ (.A0(\w[49][24] ),
    .A1(\w[51][24] ),
    .A2(\w[53][24] ),
    .A3(\w[55][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05163_));
 sky130_fd_sc_hd__mux4_2 _18678_ (.A0(\w[57][24] ),
    .A1(\w[59][24] ),
    .A2(\w[61][24] ),
    .A3(\w[63][24] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05164_));
 sky130_fd_sc_hd__mux4_2 _18679_ (.A0(_05160_),
    .A1(_05162_),
    .A2(_05163_),
    .A3(_05164_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_2 _18680_ (.A0(_05159_),
    .A1(_05165_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[24] ));
 sky130_fd_sc_hd__mux4_2 _18681_ (.A0(\w[1][25] ),
    .A1(\w[3][25] ),
    .A2(\w[5][25] ),
    .A3(\w[7][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05166_));
 sky130_fd_sc_hd__mux4_2 _18682_ (.A0(\w[9][25] ),
    .A1(\w[11][25] ),
    .A2(\w[13][25] ),
    .A3(\w[15][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05167_));
 sky130_fd_sc_hd__mux4_2 _18683_ (.A0(\w[33][25] ),
    .A1(\w[35][25] ),
    .A2(\w[37][25] ),
    .A3(\w[39][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05168_));
 sky130_fd_sc_hd__mux4_2 _18685_ (.A0(\w[41][25] ),
    .A1(\w[43][25] ),
    .A2(\w[45][25] ),
    .A3(\w[47][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05170_));
 sky130_fd_sc_hd__mux4_2 _18687_ (.A0(_05166_),
    .A1(_05167_),
    .A2(_05168_),
    .A3(_05170_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05172_));
 sky130_fd_sc_hd__mux4_2 _18688_ (.A0(\w[17][25] ),
    .A1(\w[19][25] ),
    .A2(\w[21][25] ),
    .A3(\w[23][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05173_));
 sky130_fd_sc_hd__mux4_2 _18690_ (.A0(\w[25][25] ),
    .A1(\w[27][25] ),
    .A2(\w[29][25] ),
    .A3(\w[31][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05175_));
 sky130_fd_sc_hd__mux4_2 _18691_ (.A0(\w[49][25] ),
    .A1(\w[51][25] ),
    .A2(\w[53][25] ),
    .A3(\w[55][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05176_));
 sky130_fd_sc_hd__mux4_2 _18692_ (.A0(\w[57][25] ),
    .A1(\w[59][25] ),
    .A2(\w[61][25] ),
    .A3(\w[63][25] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05177_));
 sky130_fd_sc_hd__mux4_2 _18694_ (.A0(_05173_),
    .A1(_05175_),
    .A2(_05176_),
    .A3(_05177_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05179_));
 sky130_fd_sc_hd__mux2_2 _18695_ (.A0(_05172_),
    .A1(_05179_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[25] ));
 sky130_fd_sc_hd__mux4_2 _18696_ (.A0(\w[1][26] ),
    .A1(\w[3][26] ),
    .A2(\w[5][26] ),
    .A3(\w[7][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05180_));
 sky130_fd_sc_hd__mux4_2 _18697_ (.A0(\w[9][26] ),
    .A1(\w[11][26] ),
    .A2(\w[13][26] ),
    .A3(\w[15][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05181_));
 sky130_fd_sc_hd__mux4_2 _18699_ (.A0(\w[33][26] ),
    .A1(\w[35][26] ),
    .A2(\w[37][26] ),
    .A3(\w[39][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05183_));
 sky130_fd_sc_hd__mux4_2 _18700_ (.A0(\w[41][26] ),
    .A1(\w[43][26] ),
    .A2(\w[45][26] ),
    .A3(\w[47][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05184_));
 sky130_fd_sc_hd__mux4_2 _18701_ (.A0(_05180_),
    .A1(_05181_),
    .A2(_05183_),
    .A3(_05184_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05185_));
 sky130_fd_sc_hd__mux4_2 _18702_ (.A0(\w[17][26] ),
    .A1(\w[19][26] ),
    .A2(\w[21][26] ),
    .A3(\w[23][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05186_));
 sky130_fd_sc_hd__mux4_2 _18703_ (.A0(\w[25][26] ),
    .A1(\w[27][26] ),
    .A2(\w[29][26] ),
    .A3(\w[31][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05187_));
 sky130_fd_sc_hd__mux4_2 _18704_ (.A0(\w[49][26] ),
    .A1(\w[51][26] ),
    .A2(\w[53][26] ),
    .A3(\w[55][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05188_));
 sky130_fd_sc_hd__mux4_2 _18706_ (.A0(\w[57][26] ),
    .A1(\w[59][26] ),
    .A2(\w[61][26] ),
    .A3(\w[63][26] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05190_));
 sky130_fd_sc_hd__mux4_2 _18707_ (.A0(_05186_),
    .A1(_05187_),
    .A2(_05188_),
    .A3(_05190_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05191_));
 sky130_fd_sc_hd__mux2_2 _18708_ (.A0(_05185_),
    .A1(_05191_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[26] ));
 sky130_fd_sc_hd__mux4_2 _18709_ (.A0(\w[1][27] ),
    .A1(\w[3][27] ),
    .A2(\w[5][27] ),
    .A3(\w[7][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05192_));
 sky130_fd_sc_hd__mux4_2 _18710_ (.A0(\w[9][27] ),
    .A1(\w[11][27] ),
    .A2(\w[13][27] ),
    .A3(\w[15][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05193_));
 sky130_fd_sc_hd__mux4_2 _18712_ (.A0(\w[33][27] ),
    .A1(\w[35][27] ),
    .A2(\w[37][27] ),
    .A3(\w[39][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05195_));
 sky130_fd_sc_hd__mux4_2 _18713_ (.A0(\w[41][27] ),
    .A1(\w[43][27] ),
    .A2(\w[45][27] ),
    .A3(\w[47][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05196_));
 sky130_fd_sc_hd__mux4_2 _18714_ (.A0(_05192_),
    .A1(_05193_),
    .A2(_05195_),
    .A3(_05196_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05197_));
 sky130_fd_sc_hd__mux4_2 _18715_ (.A0(\w[17][27] ),
    .A1(\w[19][27] ),
    .A2(\w[21][27] ),
    .A3(\w[23][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05198_));
 sky130_fd_sc_hd__mux4_2 _18716_ (.A0(\w[25][27] ),
    .A1(\w[27][27] ),
    .A2(\w[29][27] ),
    .A3(\w[31][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05199_));
 sky130_fd_sc_hd__mux4_2 _18717_ (.A0(\w[49][27] ),
    .A1(\w[51][27] ),
    .A2(\w[53][27] ),
    .A3(\w[55][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05200_));
 sky130_fd_sc_hd__mux4_2 _18719_ (.A0(\w[57][27] ),
    .A1(\w[59][27] ),
    .A2(\w[61][27] ),
    .A3(\w[63][27] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05202_));
 sky130_fd_sc_hd__mux4_2 _18721_ (.A0(_05198_),
    .A1(_05199_),
    .A2(_05200_),
    .A3(_05202_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05204_));
 sky130_fd_sc_hd__mux2_2 _18723_ (.A0(_05197_),
    .A1(_05204_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[27] ));
 sky130_fd_sc_hd__mux4_2 _18724_ (.A0(\w[1][28] ),
    .A1(\w[3][28] ),
    .A2(\w[5][28] ),
    .A3(\w[7][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05206_));
 sky130_fd_sc_hd__mux4_2 _18725_ (.A0(\w[9][28] ),
    .A1(\w[11][28] ),
    .A2(\w[13][28] ),
    .A3(\w[15][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05207_));
 sky130_fd_sc_hd__mux4_2 _18726_ (.A0(\w[33][28] ),
    .A1(\w[35][28] ),
    .A2(\w[37][28] ),
    .A3(\w[39][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05208_));
 sky130_fd_sc_hd__mux4_2 _18727_ (.A0(\w[41][28] ),
    .A1(\w[43][28] ),
    .A2(\w[45][28] ),
    .A3(\w[47][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05209_));
 sky130_fd_sc_hd__mux4_2 _18728_ (.A0(_05206_),
    .A1(_05207_),
    .A2(_05208_),
    .A3(_05209_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05210_));
 sky130_fd_sc_hd__mux4_2 _18729_ (.A0(\w[17][28] ),
    .A1(\w[19][28] ),
    .A2(\w[21][28] ),
    .A3(\w[23][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05211_));
 sky130_fd_sc_hd__mux4_2 _18730_ (.A0(\w[25][28] ),
    .A1(\w[27][28] ),
    .A2(\w[29][28] ),
    .A3(\w[31][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05212_));
 sky130_fd_sc_hd__mux4_2 _18732_ (.A0(\w[49][28] ),
    .A1(\w[51][28] ),
    .A2(\w[53][28] ),
    .A3(\w[55][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05214_));
 sky130_fd_sc_hd__mux4_2 _18733_ (.A0(\w[57][28] ),
    .A1(\w[59][28] ),
    .A2(\w[61][28] ),
    .A3(\w[63][28] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05215_));
 sky130_fd_sc_hd__mux4_2 _18734_ (.A0(_05211_),
    .A1(_05212_),
    .A2(_05214_),
    .A3(_05215_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05216_));
 sky130_fd_sc_hd__mux2_2 _18735_ (.A0(_05210_),
    .A1(_05216_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[28] ));
 sky130_fd_sc_hd__mux4_2 _18736_ (.A0(\w[1][29] ),
    .A1(\w[3][29] ),
    .A2(\w[5][29] ),
    .A3(\w[7][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05217_));
 sky130_fd_sc_hd__mux4_2 _18737_ (.A0(\w[9][29] ),
    .A1(\w[11][29] ),
    .A2(\w[13][29] ),
    .A3(\w[15][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05218_));
 sky130_fd_sc_hd__mux4_2 _18738_ (.A0(\w[33][29] ),
    .A1(\w[35][29] ),
    .A2(\w[37][29] ),
    .A3(\w[39][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05219_));
 sky130_fd_sc_hd__mux4_2 _18739_ (.A0(\w[41][29] ),
    .A1(\w[43][29] ),
    .A2(\w[45][29] ),
    .A3(\w[47][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05220_));
 sky130_fd_sc_hd__mux4_2 _18740_ (.A0(_05217_),
    .A1(_05218_),
    .A2(_05219_),
    .A3(_05220_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05221_));
 sky130_fd_sc_hd__mux4_2 _18741_ (.A0(\w[17][29] ),
    .A1(\w[19][29] ),
    .A2(\w[21][29] ),
    .A3(\w[23][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05222_));
 sky130_fd_sc_hd__mux4_2 _18742_ (.A0(\w[25][29] ),
    .A1(\w[27][29] ),
    .A2(\w[29][29] ),
    .A3(\w[31][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05223_));
 sky130_fd_sc_hd__mux4_2 _18744_ (.A0(\w[49][29] ),
    .A1(\w[51][29] ),
    .A2(\w[53][29] ),
    .A3(\w[55][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05225_));
 sky130_fd_sc_hd__mux4_2 _18745_ (.A0(\w[57][29] ),
    .A1(\w[59][29] ),
    .A2(\w[61][29] ),
    .A3(\w[63][29] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05226_));
 sky130_fd_sc_hd__mux4_2 _18746_ (.A0(_05222_),
    .A1(_05223_),
    .A2(_05225_),
    .A3(_05226_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05227_));
 sky130_fd_sc_hd__mux2_2 _18747_ (.A0(_05221_),
    .A1(_05227_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[29] ));
 sky130_fd_sc_hd__mux4_2 _18749_ (.A0(\w[1][2] ),
    .A1(\w[3][2] ),
    .A2(\w[5][2] ),
    .A3(\w[7][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05229_));
 sky130_fd_sc_hd__mux4_2 _18750_ (.A0(\w[9][2] ),
    .A1(\w[11][2] ),
    .A2(\w[13][2] ),
    .A3(\w[15][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05230_));
 sky130_fd_sc_hd__mux4_2 _18751_ (.A0(\w[33][2] ),
    .A1(\w[35][2] ),
    .A2(\w[37][2] ),
    .A3(\w[39][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05231_));
 sky130_fd_sc_hd__mux4_2 _18752_ (.A0(\w[41][2] ),
    .A1(\w[43][2] ),
    .A2(\w[45][2] ),
    .A3(\w[47][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05232_));
 sky130_fd_sc_hd__mux4_2 _18753_ (.A0(_05229_),
    .A1(_05230_),
    .A2(_05231_),
    .A3(_05232_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05233_));
 sky130_fd_sc_hd__mux4_2 _18754_ (.A0(\w[17][2] ),
    .A1(\w[19][2] ),
    .A2(\w[21][2] ),
    .A3(\w[23][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05234_));
 sky130_fd_sc_hd__mux4_2 _18755_ (.A0(\w[25][2] ),
    .A1(\w[27][2] ),
    .A2(\w[29][2] ),
    .A3(\w[31][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05235_));
 sky130_fd_sc_hd__mux4_2 _18756_ (.A0(\w[49][2] ),
    .A1(\w[51][2] ),
    .A2(\w[53][2] ),
    .A3(\w[55][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05236_));
 sky130_fd_sc_hd__mux4_2 _18757_ (.A0(\w[57][2] ),
    .A1(\w[59][2] ),
    .A2(\w[61][2] ),
    .A3(\w[63][2] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05237_));
 sky130_fd_sc_hd__mux4_2 _18758_ (.A0(_05234_),
    .A1(_05235_),
    .A2(_05236_),
    .A3(_05237_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05238_));
 sky130_fd_sc_hd__mux2_2 _18759_ (.A0(_05233_),
    .A1(_05238_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[2] ));
 sky130_fd_sc_hd__mux4_2 _18760_ (.A0(\w[1][30] ),
    .A1(\w[3][30] ),
    .A2(\w[5][30] ),
    .A3(\w[7][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05239_));
 sky130_fd_sc_hd__mux4_2 _18761_ (.A0(\w[9][30] ),
    .A1(\w[11][30] ),
    .A2(\w[13][30] ),
    .A3(\w[15][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05240_));
 sky130_fd_sc_hd__mux4_2 _18762_ (.A0(\w[33][30] ),
    .A1(\w[35][30] ),
    .A2(\w[37][30] ),
    .A3(\w[39][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05241_));
 sky130_fd_sc_hd__mux4_2 _18763_ (.A0(\w[41][30] ),
    .A1(\w[43][30] ),
    .A2(\w[45][30] ),
    .A3(\w[47][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05242_));
 sky130_fd_sc_hd__mux4_2 _18764_ (.A0(_05239_),
    .A1(_05240_),
    .A2(_05241_),
    .A3(_05242_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05243_));
 sky130_fd_sc_hd__mux4_2 _18765_ (.A0(\w[17][30] ),
    .A1(\w[19][30] ),
    .A2(\w[21][30] ),
    .A3(\w[23][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05244_));
 sky130_fd_sc_hd__mux4_2 _18766_ (.A0(\w[25][30] ),
    .A1(\w[27][30] ),
    .A2(\w[29][30] ),
    .A3(\w[31][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05245_));
 sky130_fd_sc_hd__mux4_2 _18767_ (.A0(\w[49][30] ),
    .A1(\w[51][30] ),
    .A2(\w[53][30] ),
    .A3(\w[55][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05246_));
 sky130_fd_sc_hd__mux4_2 _18768_ (.A0(\w[57][30] ),
    .A1(\w[59][30] ),
    .A2(\w[61][30] ),
    .A3(\w[63][30] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05247_));
 sky130_fd_sc_hd__mux4_2 _18769_ (.A0(_05244_),
    .A1(_05245_),
    .A2(_05246_),
    .A3(_05247_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_2 _18770_ (.A0(_05243_),
    .A1(_05248_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[30] ));
 sky130_fd_sc_hd__mux4_2 _18771_ (.A0(\w[1][31] ),
    .A1(\w[3][31] ),
    .A2(\w[5][31] ),
    .A3(\w[7][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05249_));
 sky130_fd_sc_hd__mux4_2 _18772_ (.A0(\w[9][31] ),
    .A1(\w[11][31] ),
    .A2(\w[13][31] ),
    .A3(\w[15][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05250_));
 sky130_fd_sc_hd__mux4_2 _18773_ (.A0(\w[33][31] ),
    .A1(\w[35][31] ),
    .A2(\w[37][31] ),
    .A3(\w[39][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05251_));
 sky130_fd_sc_hd__mux4_2 _18774_ (.A0(\w[41][31] ),
    .A1(\w[43][31] ),
    .A2(\w[45][31] ),
    .A3(\w[47][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05252_));
 sky130_fd_sc_hd__mux4_2 _18775_ (.A0(_05249_),
    .A1(_05250_),
    .A2(_05251_),
    .A3(_05252_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05253_));
 sky130_fd_sc_hd__mux4_2 _18776_ (.A0(\w[17][31] ),
    .A1(\w[19][31] ),
    .A2(\w[21][31] ),
    .A3(\w[23][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05254_));
 sky130_fd_sc_hd__mux4_2 _18777_ (.A0(\w[25][31] ),
    .A1(\w[27][31] ),
    .A2(\w[29][31] ),
    .A3(\w[31][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05255_));
 sky130_fd_sc_hd__mux4_2 _18778_ (.A0(\w[49][31] ),
    .A1(\w[51][31] ),
    .A2(\w[53][31] ),
    .A3(\w[55][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05256_));
 sky130_fd_sc_hd__mux4_2 _18779_ (.A0(\w[57][31] ),
    .A1(\w[59][31] ),
    .A2(\w[61][31] ),
    .A3(\w[63][31] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05257_));
 sky130_fd_sc_hd__mux4_2 _18780_ (.A0(_05254_),
    .A1(_05255_),
    .A2(_05256_),
    .A3(_05257_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05258_));
 sky130_fd_sc_hd__mux2_2 _18781_ (.A0(_05253_),
    .A1(_05258_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[31] ));
 sky130_fd_sc_hd__mux4_2 _18782_ (.A0(\w[1][3] ),
    .A1(\w[3][3] ),
    .A2(\w[5][3] ),
    .A3(\w[7][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05259_));
 sky130_fd_sc_hd__mux4_2 _18783_ (.A0(\w[9][3] ),
    .A1(\w[11][3] ),
    .A2(\w[13][3] ),
    .A3(\w[15][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05260_));
 sky130_fd_sc_hd__mux4_2 _18784_ (.A0(\w[33][3] ),
    .A1(\w[35][3] ),
    .A2(\w[37][3] ),
    .A3(\w[39][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05261_));
 sky130_fd_sc_hd__mux4_2 _18785_ (.A0(\w[41][3] ),
    .A1(\w[43][3] ),
    .A2(\w[45][3] ),
    .A3(\w[47][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05262_));
 sky130_fd_sc_hd__mux4_2 _18786_ (.A0(_05259_),
    .A1(_05260_),
    .A2(_05261_),
    .A3(_05262_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05263_));
 sky130_fd_sc_hd__mux4_2 _18787_ (.A0(\w[17][3] ),
    .A1(\w[19][3] ),
    .A2(\w[21][3] ),
    .A3(\w[23][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05264_));
 sky130_fd_sc_hd__mux4_2 _18788_ (.A0(\w[25][3] ),
    .A1(\w[27][3] ),
    .A2(\w[29][3] ),
    .A3(\w[31][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05265_));
 sky130_fd_sc_hd__mux4_2 _18789_ (.A0(\w[49][3] ),
    .A1(\w[51][3] ),
    .A2(\w[53][3] ),
    .A3(\w[55][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05266_));
 sky130_fd_sc_hd__mux4_2 _18790_ (.A0(\w[57][3] ),
    .A1(\w[59][3] ),
    .A2(\w[61][3] ),
    .A3(\w[63][3] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05267_));
 sky130_fd_sc_hd__mux4_2 _18791_ (.A0(_05264_),
    .A1(_05265_),
    .A2(_05266_),
    .A3(_05267_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_2 _18792_ (.A0(_05263_),
    .A1(_05268_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[3] ));
 sky130_fd_sc_hd__mux4_2 _18793_ (.A0(\w[1][4] ),
    .A1(\w[3][4] ),
    .A2(\w[5][4] ),
    .A3(\w[7][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05269_));
 sky130_fd_sc_hd__mux4_2 _18794_ (.A0(\w[9][4] ),
    .A1(\w[11][4] ),
    .A2(\w[13][4] ),
    .A3(\w[15][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05270_));
 sky130_fd_sc_hd__mux4_2 _18795_ (.A0(\w[33][4] ),
    .A1(\w[35][4] ),
    .A2(\w[37][4] ),
    .A3(\w[39][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05271_));
 sky130_fd_sc_hd__mux4_2 _18796_ (.A0(\w[41][4] ),
    .A1(\w[43][4] ),
    .A2(\w[45][4] ),
    .A3(\w[47][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05272_));
 sky130_fd_sc_hd__mux4_2 _18797_ (.A0(_05269_),
    .A1(_05270_),
    .A2(_05271_),
    .A3(_05272_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05273_));
 sky130_fd_sc_hd__mux4_2 _18798_ (.A0(\w[17][4] ),
    .A1(\w[19][4] ),
    .A2(\w[21][4] ),
    .A3(\w[23][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05274_));
 sky130_fd_sc_hd__mux4_2 _18799_ (.A0(\w[25][4] ),
    .A1(\w[27][4] ),
    .A2(\w[29][4] ),
    .A3(\w[31][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05275_));
 sky130_fd_sc_hd__mux4_2 _18800_ (.A0(\w[49][4] ),
    .A1(\w[51][4] ),
    .A2(\w[53][4] ),
    .A3(\w[55][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05276_));
 sky130_fd_sc_hd__mux4_2 _18801_ (.A0(\w[57][4] ),
    .A1(\w[59][4] ),
    .A2(\w[61][4] ),
    .A3(\w[63][4] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05277_));
 sky130_fd_sc_hd__mux4_2 _18802_ (.A0(_05274_),
    .A1(_05275_),
    .A2(_05276_),
    .A3(_05277_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05278_));
 sky130_fd_sc_hd__mux2_2 _18803_ (.A0(_05273_),
    .A1(_05278_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[4] ));
 sky130_fd_sc_hd__mux4_2 _18804_ (.A0(\w[1][5] ),
    .A1(\w[3][5] ),
    .A2(\w[5][5] ),
    .A3(\w[7][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05279_));
 sky130_fd_sc_hd__mux4_2 _18805_ (.A0(\w[9][5] ),
    .A1(\w[11][5] ),
    .A2(\w[13][5] ),
    .A3(\w[15][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05280_));
 sky130_fd_sc_hd__mux4_2 _18806_ (.A0(\w[33][5] ),
    .A1(\w[35][5] ),
    .A2(\w[37][5] ),
    .A3(\w[39][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05281_));
 sky130_fd_sc_hd__mux4_2 _18807_ (.A0(\w[41][5] ),
    .A1(\w[43][5] ),
    .A2(\w[45][5] ),
    .A3(\w[47][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05282_));
 sky130_fd_sc_hd__mux4_2 _18808_ (.A0(_05279_),
    .A1(_05280_),
    .A2(_05281_),
    .A3(_05282_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05283_));
 sky130_fd_sc_hd__mux4_2 _18809_ (.A0(\w[17][5] ),
    .A1(\w[19][5] ),
    .A2(\w[21][5] ),
    .A3(\w[23][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05284_));
 sky130_fd_sc_hd__mux4_2 _18810_ (.A0(\w[25][5] ),
    .A1(\w[27][5] ),
    .A2(\w[29][5] ),
    .A3(\w[31][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05285_));
 sky130_fd_sc_hd__mux4_2 _18811_ (.A0(\w[49][5] ),
    .A1(\w[51][5] ),
    .A2(\w[53][5] ),
    .A3(\w[55][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05286_));
 sky130_fd_sc_hd__mux4_2 _18812_ (.A0(\w[57][5] ),
    .A1(\w[59][5] ),
    .A2(\w[61][5] ),
    .A3(\w[63][5] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05287_));
 sky130_fd_sc_hd__mux4_2 _18813_ (.A0(_05284_),
    .A1(_05285_),
    .A2(_05286_),
    .A3(_05287_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05288_));
 sky130_fd_sc_hd__mux2_2 _18814_ (.A0(_05283_),
    .A1(_05288_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[5] ));
 sky130_fd_sc_hd__mux4_2 _18815_ (.A0(\w[1][6] ),
    .A1(\w[3][6] ),
    .A2(\w[5][6] ),
    .A3(\w[7][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05289_));
 sky130_fd_sc_hd__mux4_2 _18816_ (.A0(\w[9][6] ),
    .A1(\w[11][6] ),
    .A2(\w[13][6] ),
    .A3(\w[15][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05290_));
 sky130_fd_sc_hd__mux4_2 _18817_ (.A0(\w[33][6] ),
    .A1(\w[35][6] ),
    .A2(\w[37][6] ),
    .A3(\w[39][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05291_));
 sky130_fd_sc_hd__mux4_2 _18818_ (.A0(\w[41][6] ),
    .A1(\w[43][6] ),
    .A2(\w[45][6] ),
    .A3(\w[47][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05292_));
 sky130_fd_sc_hd__mux4_2 _18819_ (.A0(_05289_),
    .A1(_05290_),
    .A2(_05291_),
    .A3(_05292_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05293_));
 sky130_fd_sc_hd__mux4_2 _18820_ (.A0(\w[17][6] ),
    .A1(\w[19][6] ),
    .A2(\w[21][6] ),
    .A3(\w[23][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05294_));
 sky130_fd_sc_hd__mux4_2 _18821_ (.A0(\w[25][6] ),
    .A1(\w[27][6] ),
    .A2(\w[29][6] ),
    .A3(\w[31][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05295_));
 sky130_fd_sc_hd__mux4_2 _18822_ (.A0(\w[49][6] ),
    .A1(\w[51][6] ),
    .A2(\w[53][6] ),
    .A3(\w[55][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05296_));
 sky130_fd_sc_hd__mux4_2 _18823_ (.A0(\w[57][6] ),
    .A1(\w[59][6] ),
    .A2(\w[61][6] ),
    .A3(\w[63][6] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05297_));
 sky130_fd_sc_hd__mux4_2 _18824_ (.A0(_05294_),
    .A1(_05295_),
    .A2(_05296_),
    .A3(_05297_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05298_));
 sky130_fd_sc_hd__mux2_2 _18825_ (.A0(_05293_),
    .A1(_05298_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[6] ));
 sky130_fd_sc_hd__mux4_2 _18826_ (.A0(\w[1][7] ),
    .A1(\w[3][7] ),
    .A2(\w[5][7] ),
    .A3(\w[7][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05299_));
 sky130_fd_sc_hd__mux4_2 _18827_ (.A0(\w[9][7] ),
    .A1(\w[11][7] ),
    .A2(\w[13][7] ),
    .A3(\w[15][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05300_));
 sky130_fd_sc_hd__mux4_2 _18828_ (.A0(\w[33][7] ),
    .A1(\w[35][7] ),
    .A2(\w[37][7] ),
    .A3(\w[39][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05301_));
 sky130_fd_sc_hd__mux4_2 _18829_ (.A0(\w[41][7] ),
    .A1(\w[43][7] ),
    .A2(\w[45][7] ),
    .A3(\w[47][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05302_));
 sky130_fd_sc_hd__mux4_2 _18830_ (.A0(_05299_),
    .A1(_05300_),
    .A2(_05301_),
    .A3(_05302_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05303_));
 sky130_fd_sc_hd__mux4_2 _18831_ (.A0(\w[17][7] ),
    .A1(\w[19][7] ),
    .A2(\w[21][7] ),
    .A3(\w[23][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05304_));
 sky130_fd_sc_hd__mux4_2 _18832_ (.A0(\w[25][7] ),
    .A1(\w[27][7] ),
    .A2(\w[29][7] ),
    .A3(\w[31][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05305_));
 sky130_fd_sc_hd__mux4_2 _18833_ (.A0(\w[49][7] ),
    .A1(\w[51][7] ),
    .A2(\w[53][7] ),
    .A3(\w[55][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05306_));
 sky130_fd_sc_hd__mux4_2 _18834_ (.A0(\w[57][7] ),
    .A1(\w[59][7] ),
    .A2(\w[61][7] ),
    .A3(\w[63][7] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05307_));
 sky130_fd_sc_hd__mux4_2 _18835_ (.A0(_05304_),
    .A1(_05305_),
    .A2(_05306_),
    .A3(_05307_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_2 _18836_ (.A0(_05303_),
    .A1(_05308_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[7] ));
 sky130_fd_sc_hd__mux4_2 _18837_ (.A0(\w[1][8] ),
    .A1(\w[3][8] ),
    .A2(\w[5][8] ),
    .A3(\w[7][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05309_));
 sky130_fd_sc_hd__mux4_2 _18838_ (.A0(\w[9][8] ),
    .A1(\w[11][8] ),
    .A2(\w[13][8] ),
    .A3(\w[15][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05310_));
 sky130_fd_sc_hd__mux4_2 _18839_ (.A0(\w[33][8] ),
    .A1(\w[35][8] ),
    .A2(\w[37][8] ),
    .A3(\w[39][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05311_));
 sky130_fd_sc_hd__mux4_2 _18840_ (.A0(\w[41][8] ),
    .A1(\w[43][8] ),
    .A2(\w[45][8] ),
    .A3(\w[47][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05312_));
 sky130_fd_sc_hd__mux4_2 _18841_ (.A0(_05309_),
    .A1(_05310_),
    .A2(_05311_),
    .A3(_05312_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05313_));
 sky130_fd_sc_hd__mux4_2 _18842_ (.A0(\w[17][8] ),
    .A1(\w[19][8] ),
    .A2(\w[21][8] ),
    .A3(\w[23][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05314_));
 sky130_fd_sc_hd__mux4_2 _18843_ (.A0(\w[25][8] ),
    .A1(\w[27][8] ),
    .A2(\w[29][8] ),
    .A3(\w[31][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05315_));
 sky130_fd_sc_hd__mux4_2 _18844_ (.A0(\w[49][8] ),
    .A1(\w[51][8] ),
    .A2(\w[53][8] ),
    .A3(\w[55][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05316_));
 sky130_fd_sc_hd__mux4_2 _18845_ (.A0(\w[57][8] ),
    .A1(\w[59][8] ),
    .A2(\w[61][8] ),
    .A3(\w[63][8] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05317_));
 sky130_fd_sc_hd__mux4_2 _18846_ (.A0(_05314_),
    .A1(_05315_),
    .A2(_05316_),
    .A3(_05317_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05318_));
 sky130_fd_sc_hd__mux2_2 _18847_ (.A0(_05313_),
    .A1(_05318_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[8] ));
 sky130_fd_sc_hd__mux4_2 _18848_ (.A0(\w[1][9] ),
    .A1(\w[3][9] ),
    .A2(\w[5][9] ),
    .A3(\w[7][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05319_));
 sky130_fd_sc_hd__mux4_2 _18849_ (.A0(\w[9][9] ),
    .A1(\w[11][9] ),
    .A2(\w[13][9] ),
    .A3(\w[15][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05320_));
 sky130_fd_sc_hd__mux4_2 _18850_ (.A0(\w[33][9] ),
    .A1(\w[35][9] ),
    .A2(\w[37][9] ),
    .A3(\w[39][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05321_));
 sky130_fd_sc_hd__mux4_2 _18851_ (.A0(\w[41][9] ),
    .A1(\w[43][9] ),
    .A2(\w[45][9] ),
    .A3(\w[47][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05322_));
 sky130_fd_sc_hd__mux4_2 _18852_ (.A0(_05319_),
    .A1(_05320_),
    .A2(_05321_),
    .A3(_05322_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05323_));
 sky130_fd_sc_hd__mux4_2 _18853_ (.A0(\w[17][9] ),
    .A1(\w[19][9] ),
    .A2(\w[21][9] ),
    .A3(\w[23][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05324_));
 sky130_fd_sc_hd__mux4_2 _18854_ (.A0(\w[25][9] ),
    .A1(\w[27][9] ),
    .A2(\w[29][9] ),
    .A3(\w[31][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05325_));
 sky130_fd_sc_hd__mux4_2 _18855_ (.A0(\w[49][9] ),
    .A1(\w[51][9] ),
    .A2(\w[53][9] ),
    .A3(\w[55][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05326_));
 sky130_fd_sc_hd__mux4_2 _18856_ (.A0(\w[57][9] ),
    .A1(\w[59][9] ),
    .A2(\w[61][9] ),
    .A3(\w[63][9] ),
    .S0(\count2_2[1] ),
    .S1(\count2_2[2] ),
    .X(_05327_));
 sky130_fd_sc_hd__mux4_2 _18857_ (.A0(_05324_),
    .A1(_05325_),
    .A2(_05326_),
    .A3(_05327_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[5] ),
    .X(_05328_));
 sky130_fd_sc_hd__mux2_2 _18858_ (.A0(_05323_),
    .A1(_05328_),
    .S(\count2_2[4] ),
    .X(\w_new_calc2.w_2[9] ));
 sky130_fd_sc_hd__fa_1 _18859_ (.A(\w_new_calc1.temp2[0] ),
    .B(\w_new_calc1.temp1[0] ),
    .CIN(_08822_),
    .COUT(_08823_),
    .SUM(_08824_));
 sky130_fd_sc_hd__fa_1 _18860_ (.A(\w_new_calc1.temp2[1] ),
    .B(\w_new_calc1.temp1[1] ),
    .CIN(_08825_),
    .COUT(_08826_),
    .SUM(_08827_));
 sky130_fd_sc_hd__fa_1 _18861_ (.A(_08828_),
    .B(_08829_),
    .CIN(_08830_),
    .COUT(_08831_),
    .SUM(_08832_));
 sky130_fd_sc_hd__fa_1 _18862_ (.A(\w_new_calc1.temp2[2] ),
    .B(\w_new_calc1.temp1[2] ),
    .CIN(_08833_),
    .COUT(_08834_),
    .SUM(_08835_));
 sky130_fd_sc_hd__fa_1 _18863_ (.A(_08836_),
    .B(_08837_),
    .CIN(_08838_),
    .COUT(_08839_),
    .SUM(_08840_));
 sky130_fd_sc_hd__fa_1 _18864_ (.A(_08841_),
    .B(_08842_),
    .CIN(_08843_),
    .COUT(_08844_),
    .SUM(_08845_));
 sky130_fd_sc_hd__fa_1 _18865_ (.A(\w_new_calc1.temp2[3] ),
    .B(\w_new_calc1.temp1[3] ),
    .CIN(_08846_),
    .COUT(_08847_),
    .SUM(_08848_));
 sky130_fd_sc_hd__fa_1 _18866_ (.A(_08849_),
    .B(_08850_),
    .CIN(_08851_),
    .COUT(_08852_),
    .SUM(_08853_));
 sky130_fd_sc_hd__fa_1 _18867_ (.A(\w_new_calc1.temp2[4] ),
    .B(\w_new_calc1.temp1[4] ),
    .CIN(_08854_),
    .COUT(_08855_),
    .SUM(_08856_));
 sky130_fd_sc_hd__fa_1 _18868_ (.A(_08857_),
    .B(_08858_),
    .CIN(_08859_),
    .COUT(_08860_),
    .SUM(_08861_));
 sky130_fd_sc_hd__fa_1 _18869_ (.A(\w_new_calc1.temp2[5] ),
    .B(\w_new_calc1.temp1[5] ),
    .CIN(_08862_),
    .COUT(_08863_),
    .SUM(_08864_));
 sky130_fd_sc_hd__fa_1 _18870_ (.A(_08865_),
    .B(_08866_),
    .CIN(_08867_),
    .COUT(_08868_),
    .SUM(_08869_));
 sky130_fd_sc_hd__fa_1 _18871_ (.A(\w_new_calc1.temp2[6] ),
    .B(\w_new_calc1.temp1[6] ),
    .CIN(_08870_),
    .COUT(_08871_),
    .SUM(_08872_));
 sky130_fd_sc_hd__fa_1 _18872_ (.A(_08873_),
    .B(_08874_),
    .CIN(_08875_),
    .COUT(_08876_),
    .SUM(_08877_));
 sky130_fd_sc_hd__fa_1 _18873_ (.A(\w_new_calc1.temp2[7] ),
    .B(\w_new_calc1.temp1[7] ),
    .CIN(_08878_),
    .COUT(_08879_),
    .SUM(_08880_));
 sky130_fd_sc_hd__fa_1 _18874_ (.A(_08881_),
    .B(_08882_),
    .CIN(_08883_),
    .COUT(_08884_),
    .SUM(_08885_));
 sky130_fd_sc_hd__fa_1 _18875_ (.A(\w_new_calc1.temp2[8] ),
    .B(\w_new_calc1.temp1[8] ),
    .CIN(_08886_),
    .COUT(_08887_),
    .SUM(_08888_));
 sky130_fd_sc_hd__fa_1 _18876_ (.A(_08889_),
    .B(_08890_),
    .CIN(_08891_),
    .COUT(_08892_),
    .SUM(_08893_));
 sky130_fd_sc_hd__fa_1 _18877_ (.A(\w_new_calc1.temp2[9] ),
    .B(\w_new_calc1.temp1[9] ),
    .CIN(_08894_),
    .COUT(_08895_),
    .SUM(_08896_));
 sky130_fd_sc_hd__fa_1 _18878_ (.A(_08897_),
    .B(_08898_),
    .CIN(_08899_),
    .COUT(_08900_),
    .SUM(_08901_));
 sky130_fd_sc_hd__fa_1 _18879_ (.A(\w_new_calc1.temp2[10] ),
    .B(\w_new_calc1.temp1[10] ),
    .CIN(_08902_),
    .COUT(_08903_),
    .SUM(_08904_));
 sky130_fd_sc_hd__fa_1 _18880_ (.A(_08905_),
    .B(_08906_),
    .CIN(_08907_),
    .COUT(_08908_),
    .SUM(_08909_));
 sky130_fd_sc_hd__fa_1 _18881_ (.A(\w_new_calc1.temp2[11] ),
    .B(\w_new_calc1.temp1[11] ),
    .CIN(_08910_),
    .COUT(_08911_),
    .SUM(_08912_));
 sky130_fd_sc_hd__fa_1 _18882_ (.A(_08913_),
    .B(_08914_),
    .CIN(_08915_),
    .COUT(_08916_),
    .SUM(_08917_));
 sky130_fd_sc_hd__fa_1 _18883_ (.A(\w_new_calc1.temp2[12] ),
    .B(\w_new_calc1.temp1[12] ),
    .CIN(_08918_),
    .COUT(_08919_),
    .SUM(_08920_));
 sky130_fd_sc_hd__fa_1 _18884_ (.A(_08921_),
    .B(_08922_),
    .CIN(_08923_),
    .COUT(_08924_),
    .SUM(_08925_));
 sky130_fd_sc_hd__fa_1 _18885_ (.A(\w_new_calc1.temp2[13] ),
    .B(\w_new_calc1.temp1[13] ),
    .CIN(_08926_),
    .COUT(_08927_),
    .SUM(_08928_));
 sky130_fd_sc_hd__fa_1 _18886_ (.A(_08929_),
    .B(_08930_),
    .CIN(_08931_),
    .COUT(_08932_),
    .SUM(_08933_));
 sky130_fd_sc_hd__fa_1 _18887_ (.A(\w_new_calc1.temp2[14] ),
    .B(\w_new_calc1.temp1[14] ),
    .CIN(_08934_),
    .COUT(_08935_),
    .SUM(_08936_));
 sky130_fd_sc_hd__fa_1 _18888_ (.A(_08937_),
    .B(_08938_),
    .CIN(_08939_),
    .COUT(_08940_),
    .SUM(_08941_));
 sky130_fd_sc_hd__fa_1 _18889_ (.A(\w_new_calc1.temp2[15] ),
    .B(\w_new_calc1.temp1[15] ),
    .CIN(_08942_),
    .COUT(_08943_),
    .SUM(_08944_));
 sky130_fd_sc_hd__fa_1 _18890_ (.A(_08945_),
    .B(_08946_),
    .CIN(_08947_),
    .COUT(_08948_),
    .SUM(_08949_));
 sky130_fd_sc_hd__fa_1 _18891_ (.A(\w_new_calc1.temp2[16] ),
    .B(\w_new_calc1.temp1[16] ),
    .CIN(_08950_),
    .COUT(_08951_),
    .SUM(_08952_));
 sky130_fd_sc_hd__fa_1 _18892_ (.A(_08953_),
    .B(_08954_),
    .CIN(_08955_),
    .COUT(_08956_),
    .SUM(_08957_));
 sky130_fd_sc_hd__fa_1 _18893_ (.A(\w_new_calc1.temp2[17] ),
    .B(\w_new_calc1.temp1[17] ),
    .CIN(_08958_),
    .COUT(_08959_),
    .SUM(_08960_));
 sky130_fd_sc_hd__fa_1 _18894_ (.A(_08961_),
    .B(_08962_),
    .CIN(_08963_),
    .COUT(_08964_),
    .SUM(_08965_));
 sky130_fd_sc_hd__fa_1 _18895_ (.A(\w_new_calc1.temp2[18] ),
    .B(\w_new_calc1.temp1[18] ),
    .CIN(_08966_),
    .COUT(_08967_),
    .SUM(_08968_));
 sky130_fd_sc_hd__fa_1 _18896_ (.A(_08969_),
    .B(_08970_),
    .CIN(_08971_),
    .COUT(_08972_),
    .SUM(_08973_));
 sky130_fd_sc_hd__fa_1 _18897_ (.A(\w_new_calc1.temp2[19] ),
    .B(\w_new_calc1.temp1[19] ),
    .CIN(_08974_),
    .COUT(_08975_),
    .SUM(_08976_));
 sky130_fd_sc_hd__fa_1 _18898_ (.A(_08977_),
    .B(_08978_),
    .CIN(_08979_),
    .COUT(_08980_),
    .SUM(_08981_));
 sky130_fd_sc_hd__fa_1 _18899_ (.A(\w_new_calc1.temp2[20] ),
    .B(\w_new_calc1.temp1[20] ),
    .CIN(_08982_),
    .COUT(_08983_),
    .SUM(_08984_));
 sky130_fd_sc_hd__fa_1 _18900_ (.A(_08985_),
    .B(_08986_),
    .CIN(_08987_),
    .COUT(_08988_),
    .SUM(_08989_));
 sky130_fd_sc_hd__fa_1 _18901_ (.A(\w_new_calc1.temp2[21] ),
    .B(\w_new_calc1.temp1[21] ),
    .CIN(_08990_),
    .COUT(_08991_),
    .SUM(_08992_));
 sky130_fd_sc_hd__fa_1 _18902_ (.A(_08993_),
    .B(_08994_),
    .CIN(_08995_),
    .COUT(_08996_),
    .SUM(_08997_));
 sky130_fd_sc_hd__fa_1 _18903_ (.A(\w_new_calc1.temp2[22] ),
    .B(\w_new_calc1.temp1[22] ),
    .CIN(_08998_),
    .COUT(_08999_),
    .SUM(_09000_));
 sky130_fd_sc_hd__fa_1 _18904_ (.A(_09001_),
    .B(_09002_),
    .CIN(_09003_),
    .COUT(_09004_),
    .SUM(_09005_));
 sky130_fd_sc_hd__fa_1 _18905_ (.A(\w_new_calc1.temp2[23] ),
    .B(\w_new_calc1.temp1[23] ),
    .CIN(_09006_),
    .COUT(_09007_),
    .SUM(_09008_));
 sky130_fd_sc_hd__fa_1 _18906_ (.A(_09009_),
    .B(_09010_),
    .CIN(_09011_),
    .COUT(_09012_),
    .SUM(_09013_));
 sky130_fd_sc_hd__fa_1 _18907_ (.A(\w_new_calc1.temp2[24] ),
    .B(\w_new_calc1.temp1[24] ),
    .CIN(_09014_),
    .COUT(_09015_),
    .SUM(_09016_));
 sky130_fd_sc_hd__fa_1 _18908_ (.A(_09017_),
    .B(_09018_),
    .CIN(_09019_),
    .COUT(_09020_),
    .SUM(_09021_));
 sky130_fd_sc_hd__fa_1 _18909_ (.A(\w_new_calc1.temp2[25] ),
    .B(\w_new_calc1.temp1[25] ),
    .CIN(_09022_),
    .COUT(_09023_),
    .SUM(_09024_));
 sky130_fd_sc_hd__fa_1 _18910_ (.A(_09025_),
    .B(_09026_),
    .CIN(_09027_),
    .COUT(_09028_),
    .SUM(_09029_));
 sky130_fd_sc_hd__fa_1 _18911_ (.A(\w_new_calc1.temp2[26] ),
    .B(\w_new_calc1.temp1[26] ),
    .CIN(_09030_),
    .COUT(_09031_),
    .SUM(_09032_));
 sky130_fd_sc_hd__fa_1 _18912_ (.A(_09033_),
    .B(_09034_),
    .CIN(_09035_),
    .COUT(_09036_),
    .SUM(_09037_));
 sky130_fd_sc_hd__fa_1 _18913_ (.A(\w_new_calc1.temp2[27] ),
    .B(\w_new_calc1.temp1[27] ),
    .CIN(_09038_),
    .COUT(_09039_),
    .SUM(_09040_));
 sky130_fd_sc_hd__fa_1 _18914_ (.A(_09041_),
    .B(_09042_),
    .CIN(_09043_),
    .COUT(_09044_),
    .SUM(_09045_));
 sky130_fd_sc_hd__fa_1 _18915_ (.A(\w_new_calc1.temp2[28] ),
    .B(\w_new_calc1.temp1[28] ),
    .CIN(_09046_),
    .COUT(_09047_),
    .SUM(_09048_));
 sky130_fd_sc_hd__fa_1 _18916_ (.A(_09049_),
    .B(_09050_),
    .CIN(_09051_),
    .COUT(_09052_),
    .SUM(_09053_));
 sky130_fd_sc_hd__fa_1 _18917_ (.A(\w_new_calc1.temp2[29] ),
    .B(\w_new_calc1.temp1[29] ),
    .CIN(_09054_),
    .COUT(_09055_),
    .SUM(_09056_));
 sky130_fd_sc_hd__fa_1 _18918_ (.A(_09057_),
    .B(_09058_),
    .CIN(_09059_),
    .COUT(_09060_),
    .SUM(_09061_));
 sky130_fd_sc_hd__fa_1 _18919_ (.A(\w_new_calc1.temp2[30] ),
    .B(\w_new_calc1.temp1[30] ),
    .CIN(_09062_),
    .COUT(_09063_),
    .SUM(_09064_));
 sky130_fd_sc_hd__fa_1 _18920_ (.A(_09065_),
    .B(_09066_),
    .CIN(_09067_),
    .COUT(_09068_),
    .SUM(_09069_));
 sky130_fd_sc_hd__fa_1 _18921_ (.A(_09070_),
    .B(_09071_),
    .CIN(_09072_),
    .COUT(_09073_),
    .SUM(_09074_));
 sky130_fd_sc_hd__fa_1 _18922_ (.A(_09075_),
    .B(_09076_),
    .CIN(_09077_),
    .COUT(_09078_),
    .SUM(_09079_));
 sky130_fd_sc_hd__fa_1 _18923_ (.A(\w_new_calc2.temp1[1] ),
    .B(_09080_),
    .CIN(_09081_),
    .COUT(_09082_),
    .SUM(_09083_));
 sky130_fd_sc_hd__fa_1 _18924_ (.A(_09084_),
    .B(_09085_),
    .CIN(_09086_),
    .COUT(_09087_),
    .SUM(_09088_));
 sky130_fd_sc_hd__fa_1 _18925_ (.A(\w_new_calc2.temp1[2] ),
    .B(_09089_),
    .CIN(_09090_),
    .COUT(_09091_),
    .SUM(_09092_));
 sky130_fd_sc_hd__fa_1 _18926_ (.A(_09093_),
    .B(_09082_),
    .CIN(_09092_),
    .COUT(_09094_),
    .SUM(_09095_));
 sky130_fd_sc_hd__fa_1 _18927_ (.A(_09096_),
    .B(_09097_),
    .CIN(_09098_),
    .COUT(_09099_),
    .SUM(_09100_));
 sky130_fd_sc_hd__fa_1 _18928_ (.A(\w_new_calc2.temp1[3] ),
    .B(_09101_),
    .CIN(_09102_),
    .COUT(_09103_),
    .SUM(_09104_));
 sky130_fd_sc_hd__fa_1 _18929_ (.A(_09105_),
    .B(_09106_),
    .CIN(_09107_),
    .COUT(_09108_),
    .SUM(_09109_));
 sky130_fd_sc_hd__fa_1 _18930_ (.A(\w_new_calc2.temp1[4] ),
    .B(_09110_),
    .CIN(_09111_),
    .COUT(_09112_),
    .SUM(_09113_));
 sky130_fd_sc_hd__fa_1 _18931_ (.A(_09114_),
    .B(_09115_),
    .CIN(_09116_),
    .COUT(_09117_),
    .SUM(_09118_));
 sky130_fd_sc_hd__fa_1 _18932_ (.A(\w_new_calc2.temp1[5] ),
    .B(_09119_),
    .CIN(_09120_),
    .COUT(_09121_),
    .SUM(_09122_));
 sky130_fd_sc_hd__fa_1 _18933_ (.A(_09123_),
    .B(_09124_),
    .CIN(_09125_),
    .COUT(_09126_),
    .SUM(_09127_));
 sky130_fd_sc_hd__fa_1 _18934_ (.A(\w_new_calc2.temp1[6] ),
    .B(_09128_),
    .CIN(_09129_),
    .COUT(_09130_),
    .SUM(_09131_));
 sky130_fd_sc_hd__fa_1 _18935_ (.A(_09132_),
    .B(_09133_),
    .CIN(_09134_),
    .COUT(_09135_),
    .SUM(_09136_));
 sky130_fd_sc_hd__fa_1 _18936_ (.A(\w_new_calc2.temp1[7] ),
    .B(_09137_),
    .CIN(_09138_),
    .COUT(_09139_),
    .SUM(_09140_));
 sky130_fd_sc_hd__fa_1 _18937_ (.A(_09141_),
    .B(_09142_),
    .CIN(_09143_),
    .COUT(_09144_),
    .SUM(_09145_));
 sky130_fd_sc_hd__fa_1 _18938_ (.A(\w_new_calc2.temp1[8] ),
    .B(_09146_),
    .CIN(_09147_),
    .COUT(_09148_),
    .SUM(_09149_));
 sky130_fd_sc_hd__fa_1 _18939_ (.A(_09150_),
    .B(_09151_),
    .CIN(_09152_),
    .COUT(_09153_),
    .SUM(_09154_));
 sky130_fd_sc_hd__fa_1 _18940_ (.A(\w_new_calc2.temp1[9] ),
    .B(_09155_),
    .CIN(_09156_),
    .COUT(_09157_),
    .SUM(_09158_));
 sky130_fd_sc_hd__fa_1 _18941_ (.A(_09159_),
    .B(_09160_),
    .CIN(_09161_),
    .COUT(_09162_),
    .SUM(_09163_));
 sky130_fd_sc_hd__fa_1 _18942_ (.A(\w_new_calc2.temp1[10] ),
    .B(_09164_),
    .CIN(_09165_),
    .COUT(_09166_),
    .SUM(_09167_));
 sky130_fd_sc_hd__fa_1 _18943_ (.A(_09168_),
    .B(_09169_),
    .CIN(_09170_),
    .COUT(_09171_),
    .SUM(_09172_));
 sky130_fd_sc_hd__fa_1 _18944_ (.A(\w_new_calc2.temp1[11] ),
    .B(_09173_),
    .CIN(_09174_),
    .COUT(_09175_),
    .SUM(_09176_));
 sky130_fd_sc_hd__fa_1 _18945_ (.A(_09177_),
    .B(_09178_),
    .CIN(_09179_),
    .COUT(_09180_),
    .SUM(_09181_));
 sky130_fd_sc_hd__fa_1 _18946_ (.A(\w_new_calc2.temp1[12] ),
    .B(_09182_),
    .CIN(_09183_),
    .COUT(_09184_),
    .SUM(_09185_));
 sky130_fd_sc_hd__fa_1 _18947_ (.A(_09186_),
    .B(_09187_),
    .CIN(_09188_),
    .COUT(_09189_),
    .SUM(_09190_));
 sky130_fd_sc_hd__fa_1 _18948_ (.A(\w_new_calc2.temp1[13] ),
    .B(_09191_),
    .CIN(_09192_),
    .COUT(_09193_),
    .SUM(_09194_));
 sky130_fd_sc_hd__fa_1 _18949_ (.A(_09195_),
    .B(_09196_),
    .CIN(_09197_),
    .COUT(_09198_),
    .SUM(_09199_));
 sky130_fd_sc_hd__fa_1 _18950_ (.A(\w_new_calc2.temp1[14] ),
    .B(_09200_),
    .CIN(_09201_),
    .COUT(_09202_),
    .SUM(_09203_));
 sky130_fd_sc_hd__fa_1 _18951_ (.A(_09204_),
    .B(_09205_),
    .CIN(_09206_),
    .COUT(_09207_),
    .SUM(_09208_));
 sky130_fd_sc_hd__fa_1 _18952_ (.A(\w_new_calc2.temp1[15] ),
    .B(_09209_),
    .CIN(_09210_),
    .COUT(_09211_),
    .SUM(_09212_));
 sky130_fd_sc_hd__fa_1 _18953_ (.A(_09213_),
    .B(_09214_),
    .CIN(_09215_),
    .COUT(_09216_),
    .SUM(_09217_));
 sky130_fd_sc_hd__fa_1 _18954_ (.A(\w_new_calc2.temp1[16] ),
    .B(_09218_),
    .CIN(_09219_),
    .COUT(_09220_),
    .SUM(_09221_));
 sky130_fd_sc_hd__fa_1 _18955_ (.A(_09222_),
    .B(_09223_),
    .CIN(_09224_),
    .COUT(_09225_),
    .SUM(_09226_));
 sky130_fd_sc_hd__fa_1 _18956_ (.A(\w_new_calc2.temp1[17] ),
    .B(_09227_),
    .CIN(_09228_),
    .COUT(_09229_),
    .SUM(_09230_));
 sky130_fd_sc_hd__fa_1 _18957_ (.A(_09231_),
    .B(_09232_),
    .CIN(_09233_),
    .COUT(_09234_),
    .SUM(_09235_));
 sky130_fd_sc_hd__fa_1 _18958_ (.A(\w_new_calc2.temp1[18] ),
    .B(_09236_),
    .CIN(_09237_),
    .COUT(_09238_),
    .SUM(_09239_));
 sky130_fd_sc_hd__fa_1 _18959_ (.A(_09240_),
    .B(_09241_),
    .CIN(_09242_),
    .COUT(_09243_),
    .SUM(_09244_));
 sky130_fd_sc_hd__fa_1 _18960_ (.A(\w_new_calc2.temp1[19] ),
    .B(_09245_),
    .CIN(_09246_),
    .COUT(_09247_),
    .SUM(_09248_));
 sky130_fd_sc_hd__fa_1 _18961_ (.A(_09249_),
    .B(_09250_),
    .CIN(_09251_),
    .COUT(_09252_),
    .SUM(_09253_));
 sky130_fd_sc_hd__fa_1 _18962_ (.A(\w_new_calc2.temp1[20] ),
    .B(_09254_),
    .CIN(_09255_),
    .COUT(_09256_),
    .SUM(_09257_));
 sky130_fd_sc_hd__fa_1 _18963_ (.A(_09258_),
    .B(_09259_),
    .CIN(_09260_),
    .COUT(_09261_),
    .SUM(_09262_));
 sky130_fd_sc_hd__fa_1 _18964_ (.A(\w_new_calc2.temp1[21] ),
    .B(_09263_),
    .CIN(_09264_),
    .COUT(_09265_),
    .SUM(_09266_));
 sky130_fd_sc_hd__fa_1 _18965_ (.A(_09267_),
    .B(_09268_),
    .CIN(_09269_),
    .COUT(_09270_),
    .SUM(_09271_));
 sky130_fd_sc_hd__fa_1 _18966_ (.A(\w_new_calc2.temp1[22] ),
    .B(_09272_),
    .CIN(_09273_),
    .COUT(_09274_),
    .SUM(_09275_));
 sky130_fd_sc_hd__fa_1 _18967_ (.A(_09276_),
    .B(_09277_),
    .CIN(_09278_),
    .COUT(_09279_),
    .SUM(_09280_));
 sky130_fd_sc_hd__fa_1 _18968_ (.A(\w_new_calc2.temp1[23] ),
    .B(_09281_),
    .CIN(_09282_),
    .COUT(_09283_),
    .SUM(_09284_));
 sky130_fd_sc_hd__fa_1 _18969_ (.A(_09285_),
    .B(_09286_),
    .CIN(_09287_),
    .COUT(_09288_),
    .SUM(_09289_));
 sky130_fd_sc_hd__fa_1 _18970_ (.A(\w_new_calc2.temp1[24] ),
    .B(_09290_),
    .CIN(_09291_),
    .COUT(_09292_),
    .SUM(_09293_));
 sky130_fd_sc_hd__fa_1 _18971_ (.A(_09294_),
    .B(_09295_),
    .CIN(_09296_),
    .COUT(_09297_),
    .SUM(_09298_));
 sky130_fd_sc_hd__fa_1 _18972_ (.A(\w_new_calc2.temp1[25] ),
    .B(_09299_),
    .CIN(_09300_),
    .COUT(_09301_),
    .SUM(_09302_));
 sky130_fd_sc_hd__fa_1 _18973_ (.A(_09303_),
    .B(_09304_),
    .CIN(_09305_),
    .COUT(_09306_),
    .SUM(_09307_));
 sky130_fd_sc_hd__fa_1 _18974_ (.A(\w_new_calc2.temp1[26] ),
    .B(_09308_),
    .CIN(_09309_),
    .COUT(_09310_),
    .SUM(_09311_));
 sky130_fd_sc_hd__fa_1 _18975_ (.A(_09312_),
    .B(_09313_),
    .CIN(_09314_),
    .COUT(_09315_),
    .SUM(_09316_));
 sky130_fd_sc_hd__fa_1 _18976_ (.A(\w_new_calc2.temp1[27] ),
    .B(_09317_),
    .CIN(_09318_),
    .COUT(_09319_),
    .SUM(_09320_));
 sky130_fd_sc_hd__fa_1 _18977_ (.A(\w_new_calc2.temp2[28] ),
    .B(_09321_),
    .CIN(_09322_),
    .COUT(_09323_),
    .SUM(_09324_));
 sky130_fd_sc_hd__fa_1 _18978_ (.A(_09325_),
    .B(_09315_),
    .CIN(_09326_),
    .COUT(_09327_),
    .SUM(_09328_));
 sky130_fd_sc_hd__fa_1 _18979_ (.A(\w_new_calc2.temp2[29] ),
    .B(_09329_),
    .CIN(_09330_),
    .COUT(_09331_),
    .SUM(_09332_));
 sky130_fd_sc_hd__fa_1 _18980_ (.A(_09333_),
    .B(_09334_),
    .CIN(_09335_),
    .COUT(_09336_),
    .SUM(_09337_));
 sky130_fd_sc_hd__fa_1 _18981_ (.A(_09338_),
    .B(_09339_),
    .CIN(_09340_),
    .COUT(_09341_),
    .SUM(_09342_));
 sky130_fd_sc_hd__fa_1 _18982_ (.A(\w_new_calc2.temp1[30] ),
    .B(_09331_),
    .CIN(_09343_),
    .COUT(_09344_),
    .SUM(_09345_));
 sky130_fd_sc_hd__ha_4 _18983_ (.A(_00656_),
    .B(_09346_),
    .COUT(_09347_),
    .SUM(_00657_));
 sky130_fd_sc_hd__ha_1 _18984_ (.A(_00656_),
    .B(\count_hash2[2] ),
    .COUT(_09348_),
    .SUM(_09349_));
 sky130_fd_sc_hd__ha_1 _18985_ (.A(\count_hash2[1] ),
    .B(_09346_),
    .COUT(_09350_),
    .SUM(_09351_));
 sky130_fd_sc_hd__ha_1 _18986_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_09352_),
    .SUM(_09353_));
 sky130_fd_sc_hd__ha_1 _18987_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_09354_),
    .SUM(_09355_));
 sky130_fd_sc_hd__ha_4 _18988_ (.A(_00654_),
    .B(_09356_),
    .COUT(_09357_),
    .SUM(_00655_));
 sky130_fd_sc_hd__ha_1 _18989_ (.A(_00654_),
    .B(\count_hash1[2] ),
    .COUT(_09358_),
    .SUM(_09359_));
 sky130_fd_sc_hd__ha_1 _18990_ (.A(_00654_),
    .B(\count_hash1[2] ),
    .COUT(_09360_),
    .SUM(_09361_));
 sky130_fd_sc_hd__ha_1 _18991_ (.A(\count_hash1[1] ),
    .B(_09356_),
    .COUT(_09362_),
    .SUM(_09363_));
 sky130_fd_sc_hd__ha_1 _18992_ (.A(\count_hash1[1] ),
    .B(\count_hash1[2] ),
    .COUT(_09364_),
    .SUM(_09365_));
 sky130_fd_sc_hd__ha_1 _18993_ (.A(\count_hash1[1] ),
    .B(\count_hash1[2] ),
    .COUT(_09366_),
    .SUM(_09367_));
 sky130_fd_sc_hd__ha_1 _18994_ (.A(_09368_),
    .B(_08824_),
    .COUT(_09369_),
    .SUM(_09370_));
 sky130_fd_sc_hd__ha_1 _18995_ (.A(_09369_),
    .B(_09371_),
    .COUT(_08841_),
    .SUM(_09372_));
 sky130_fd_sc_hd__ha_1 _18996_ (.A(_08842_),
    .B(_08843_),
    .COUT(_09373_),
    .SUM(_09374_));
 sky130_fd_sc_hd__ha_1 _18997_ (.A(_09375_),
    .B(_09376_),
    .COUT(_09377_),
    .SUM(_09378_));
 sky130_fd_sc_hd__ha_1 _18998_ (.A(_09379_),
    .B(_09380_),
    .COUT(_09381_),
    .SUM(_09382_));
 sky130_fd_sc_hd__ha_1 _18999_ (.A(_09383_),
    .B(_09384_),
    .COUT(_09385_),
    .SUM(_09386_));
 sky130_fd_sc_hd__ha_1 _19000_ (.A(_09387_),
    .B(_09388_),
    .COUT(_09389_),
    .SUM(_09390_));
 sky130_fd_sc_hd__ha_1 _19001_ (.A(_09391_),
    .B(_09392_),
    .COUT(_09393_),
    .SUM(_09394_));
 sky130_fd_sc_hd__ha_1 _19002_ (.A(_09395_),
    .B(_09396_),
    .COUT(_09397_),
    .SUM(_09398_));
 sky130_fd_sc_hd__ha_1 _19003_ (.A(_09399_),
    .B(_09400_),
    .COUT(_09401_),
    .SUM(_09402_));
 sky130_fd_sc_hd__ha_1 _19004_ (.A(_09403_),
    .B(_09404_),
    .COUT(_09405_),
    .SUM(_09406_));
 sky130_fd_sc_hd__ha_1 _19005_ (.A(_09407_),
    .B(_09408_),
    .COUT(_09409_),
    .SUM(_09410_));
 sky130_fd_sc_hd__ha_1 _19006_ (.A(_09411_),
    .B(_09412_),
    .COUT(_09413_),
    .SUM(_09414_));
 sky130_fd_sc_hd__ha_1 _19007_ (.A(_09415_),
    .B(_09416_),
    .COUT(_09417_),
    .SUM(_09418_));
 sky130_fd_sc_hd__ha_1 _19008_ (.A(_09419_),
    .B(_09420_),
    .COUT(_09421_),
    .SUM(_09422_));
 sky130_fd_sc_hd__ha_1 _19009_ (.A(_09423_),
    .B(_09424_),
    .COUT(_09425_),
    .SUM(_09426_));
 sky130_fd_sc_hd__ha_1 _19010_ (.A(_09427_),
    .B(_09428_),
    .COUT(_09429_),
    .SUM(_09430_));
 sky130_fd_sc_hd__ha_1 _19011_ (.A(_09431_),
    .B(_09432_),
    .COUT(_09433_),
    .SUM(_09434_));
 sky130_fd_sc_hd__ha_1 _19012_ (.A(_09435_),
    .B(_09436_),
    .COUT(_09437_),
    .SUM(_09438_));
 sky130_fd_sc_hd__ha_1 _19013_ (.A(_09439_),
    .B(_09440_),
    .COUT(_09441_),
    .SUM(_09442_));
 sky130_fd_sc_hd__ha_1 _19014_ (.A(_09443_),
    .B(_09444_),
    .COUT(_09445_),
    .SUM(_09446_));
 sky130_fd_sc_hd__ha_1 _19015_ (.A(_09447_),
    .B(_09448_),
    .COUT(_09449_),
    .SUM(_09450_));
 sky130_fd_sc_hd__ha_1 _19016_ (.A(_09451_),
    .B(_09452_),
    .COUT(_09453_),
    .SUM(_09454_));
 sky130_fd_sc_hd__ha_1 _19017_ (.A(_09455_),
    .B(_09456_),
    .COUT(_09457_),
    .SUM(_09458_));
 sky130_fd_sc_hd__ha_1 _19018_ (.A(_09459_),
    .B(_09460_),
    .COUT(_09461_),
    .SUM(_09462_));
 sky130_fd_sc_hd__ha_1 _19019_ (.A(_09463_),
    .B(_09464_),
    .COUT(_09465_),
    .SUM(_09466_));
 sky130_fd_sc_hd__ha_1 _19020_ (.A(_09467_),
    .B(_09468_),
    .COUT(_09469_),
    .SUM(_09470_));
 sky130_fd_sc_hd__ha_1 _19021_ (.A(_09471_),
    .B(_09472_),
    .COUT(_09473_),
    .SUM(_09474_));
 sky130_fd_sc_hd__ha_1 _19022_ (.A(_09475_),
    .B(_09476_),
    .COUT(_09477_),
    .SUM(_09478_));
 sky130_fd_sc_hd__ha_1 _19023_ (.A(_09479_),
    .B(_09480_),
    .COUT(_09481_),
    .SUM(_09482_));
 sky130_fd_sc_hd__ha_1 _19024_ (.A(_09483_),
    .B(_09484_),
    .COUT(_09485_),
    .SUM(_09486_));
 sky130_fd_sc_hd__ha_1 _19025_ (.A(\w_new_calc2.temp1[0] ),
    .B(_09487_),
    .COUT(_09488_),
    .SUM(_09489_));
 sky130_fd_sc_hd__ha_1 _19026_ (.A(_09488_),
    .B(_09083_),
    .COUT(_09093_),
    .SUM(_09490_));
 sky130_fd_sc_hd__ha_1 _19027_ (.A(_09082_),
    .B(_09092_),
    .COUT(_09491_),
    .SUM(_09492_));
 sky130_fd_sc_hd__ha_1 _19028_ (.A(_09091_),
    .B(_09104_),
    .COUT(_09493_),
    .SUM(_09494_));
 sky130_fd_sc_hd__ha_1 _19029_ (.A(_09103_),
    .B(_09113_),
    .COUT(_09495_),
    .SUM(_09496_));
 sky130_fd_sc_hd__ha_1 _19030_ (.A(_09112_),
    .B(_09122_),
    .COUT(_09497_),
    .SUM(_09498_));
 sky130_fd_sc_hd__ha_1 _19031_ (.A(_09121_),
    .B(_09131_),
    .COUT(_09499_),
    .SUM(_09500_));
 sky130_fd_sc_hd__ha_1 _19032_ (.A(_09130_),
    .B(_09140_),
    .COUT(_09501_),
    .SUM(_09502_));
 sky130_fd_sc_hd__ha_1 _19033_ (.A(_09139_),
    .B(_09149_),
    .COUT(_09503_),
    .SUM(_09504_));
 sky130_fd_sc_hd__ha_1 _19034_ (.A(_09148_),
    .B(_09158_),
    .COUT(_09505_),
    .SUM(_09506_));
 sky130_fd_sc_hd__ha_1 _19035_ (.A(_09157_),
    .B(_09167_),
    .COUT(_09507_),
    .SUM(_09508_));
 sky130_fd_sc_hd__ha_1 _19036_ (.A(_09166_),
    .B(_09176_),
    .COUT(_09509_),
    .SUM(_09510_));
 sky130_fd_sc_hd__ha_1 _19037_ (.A(_09175_),
    .B(_09185_),
    .COUT(_09511_),
    .SUM(_09512_));
 sky130_fd_sc_hd__ha_1 _19038_ (.A(_09184_),
    .B(_09194_),
    .COUT(_09513_),
    .SUM(_09514_));
 sky130_fd_sc_hd__ha_1 _19039_ (.A(_09193_),
    .B(_09203_),
    .COUT(_09515_),
    .SUM(_09516_));
 sky130_fd_sc_hd__ha_1 _19040_ (.A(_09202_),
    .B(_09212_),
    .COUT(_09517_),
    .SUM(_09518_));
 sky130_fd_sc_hd__ha_1 _19041_ (.A(_09211_),
    .B(_09221_),
    .COUT(_09519_),
    .SUM(_09520_));
 sky130_fd_sc_hd__ha_1 _19042_ (.A(_09220_),
    .B(_09230_),
    .COUT(_09521_),
    .SUM(_09522_));
 sky130_fd_sc_hd__ha_1 _19043_ (.A(_09229_),
    .B(_09239_),
    .COUT(_09523_),
    .SUM(_09524_));
 sky130_fd_sc_hd__ha_1 _19044_ (.A(_09238_),
    .B(_09248_),
    .COUT(_09525_),
    .SUM(_09526_));
 sky130_fd_sc_hd__ha_1 _19045_ (.A(_09247_),
    .B(_09257_),
    .COUT(_09527_),
    .SUM(_09528_));
 sky130_fd_sc_hd__ha_1 _19046_ (.A(_09256_),
    .B(_09266_),
    .COUT(_09529_),
    .SUM(_09530_));
 sky130_fd_sc_hd__ha_1 _19047_ (.A(_09265_),
    .B(_09275_),
    .COUT(_09531_),
    .SUM(_09532_));
 sky130_fd_sc_hd__ha_1 _19048_ (.A(_09274_),
    .B(_09284_),
    .COUT(_09533_),
    .SUM(_09534_));
 sky130_fd_sc_hd__ha_1 _19049_ (.A(_09283_),
    .B(_09293_),
    .COUT(_09535_),
    .SUM(_09536_));
 sky130_fd_sc_hd__ha_1 _19050_ (.A(_09292_),
    .B(_09302_),
    .COUT(_09537_),
    .SUM(_09538_));
 sky130_fd_sc_hd__ha_1 _19051_ (.A(_09301_),
    .B(_09311_),
    .COUT(_09539_),
    .SUM(_09540_));
 sky130_fd_sc_hd__ha_1 _19052_ (.A(_09310_),
    .B(_09320_),
    .COUT(_09541_),
    .SUM(_09542_));
 sky130_fd_sc_hd__ha_1 _19053_ (.A(_09319_),
    .B(_09543_),
    .COUT(_09544_),
    .SUM(_09545_));
 sky130_fd_sc_hd__ha_1 _19054_ (.A(_09546_),
    .B(_09547_),
    .COUT(_09548_),
    .SUM(_09549_));
 sky130_fd_sc_hd__ha_1 _19055_ (.A(_09550_),
    .B(_09345_),
    .COUT(_09551_),
    .SUM(_09552_));
 sky130_fd_sc_hd__ha_1 _19056_ (.A(_00650_),
    .B(_09553_),
    .COUT(_09554_),
    .SUM(_00651_));
 sky130_fd_sc_hd__ha_1 _19057_ (.A(_00650_),
    .B(\count_1[2] ),
    .COUT(_09555_),
    .SUM(_09556_));
 sky130_fd_sc_hd__ha_1 _19058_ (.A(\count_1[1] ),
    .B(_09553_),
    .COUT(_09557_),
    .SUM(_09558_));
 sky130_fd_sc_hd__ha_1 _19059_ (.A(\count_1[1] ),
    .B(\count_1[2] ),
    .COUT(_09559_),
    .SUM(_09560_));
 sky130_fd_sc_hd__ha_1 _19060_ (.A(_00652_),
    .B(_09561_),
    .COUT(_09562_),
    .SUM(_00653_));
 sky130_fd_sc_hd__ha_1 _19061_ (.A(_00652_),
    .B(\count_2[2] ),
    .COUT(_09563_),
    .SUM(_09564_));
 sky130_fd_sc_hd__ha_1 _19062_ (.A(\count_2[1] ),
    .B(_09561_),
    .COUT(_09565_),
    .SUM(_09566_));
 sky130_fd_sc_hd__ha_1 _19063_ (.A(\count_2[1] ),
    .B(\count_2[2] ),
    .COUT(_09567_),
    .SUM(_09568_));
 sky130_fd_sc_hd__ha_1 _19064_ (.A(\count2_1[1] ),
    .B(\count2_1[2] ),
    .COUT(_09569_),
    .SUM(_00642_));
 sky130_fd_sc_hd__ha_1 _19065_ (.A(\count15_2[1] ),
    .B(\count15_2[2] ),
    .COUT(_09570_),
    .SUM(_00648_));
 sky130_fd_sc_hd__ha_1 _19066_ (.A(\count16_2[1] ),
    .B(\count16_2[2] ),
    .COUT(_09571_),
    .SUM(_00649_));
 sky130_fd_sc_hd__ha_1 _19067_ (.A(\count7_2[1] ),
    .B(\count7_2[2] ),
    .COUT(_09572_),
    .SUM(_00647_));
 sky130_fd_sc_hd__ha_1 _19068_ (.A(\count2_2[1] ),
    .B(\count2_2[2] ),
    .COUT(_09573_),
    .SUM(_00646_));
 sky130_fd_sc_hd__ha_1 _19069_ (.A(\count16_1[1] ),
    .B(\count16_1[2] ),
    .COUT(_09574_),
    .SUM(_00645_));
 sky130_fd_sc_hd__ha_1 _19070_ (.A(\count15_1[1] ),
    .B(\count15_1[2] ),
    .COUT(_09575_),
    .SUM(_00644_));
 sky130_fd_sc_hd__ha_1 _19071_ (.A(\count7_1[1] ),
    .B(\count7_1[2] ),
    .COUT(_09576_),
    .SUM(_00643_));
 sky130_fd_sc_hd__conb_1 _19072_ (.HI(_09577_));
 sky130_fd_sc_hd__conb_1 _19073_ (.LO(_09578_));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[1]$_SDFF_PP0_  (.D(_00658_),
    .Q(\count15_1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[2]$_SDFF_PP0_  (.D(_00659_),
    .Q(\count15_1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[3]$_SDFF_PP0_  (.D(_00660_),
    .Q(\count15_1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[4]$_SDFF_PP0_  (.D(_00661_),
    .Q(\count15_1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count15_1[5]$_SDFF_PP0_  (.D(_00662_),
    .Q(\count15_1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[1]$_SDFF_PP1_  (.D(_00663_),
    .Q(\count15_2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[2]$_SDFF_PP0_  (.D(_00664_),
    .Q(\count15_2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[3]$_SDFF_PP0_  (.D(_00665_),
    .Q(\count15_2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_2[4]$_SDFF_PP0_  (.D(_00666_),
    .Q(\count15_2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count15_2[5]$_SDFF_PP0_  (.D(_00667_),
    .Q(\count15_2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[1]$_SDFF_PP0_  (.D(_00668_),
    .Q(\count16_1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[2]$_SDFF_PP0_  (.D(_00669_),
    .Q(\count16_1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[3]$_SDFF_PP0_  (.D(_00670_),
    .Q(\count16_1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_1[4]$_SDFF_PP0_  (.D(_00671_),
    .Q(\count16_1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[5]$_SDFF_PP0_  (.D(_00672_),
    .Q(\count16_1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[1]$_SDFF_PP0_  (.D(_00673_),
    .Q(\count16_2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[2]$_SDFF_PP0_  (.D(_00674_),
    .Q(\count16_2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[3]$_SDFF_PP0_  (.D(_00675_),
    .Q(\count16_2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_2[4]$_SDFF_PP0_  (.D(_00676_),
    .Q(\count16_2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_2[5]$_SDFF_PP0_  (.D(_00677_),
    .Q(\count16_2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[1]$_SDFF_PP1_  (.D(_00678_),
    .Q(\count2_1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[2]$_SDFF_PP1_  (.D(_00679_),
    .Q(\count2_1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[3]$_SDFF_PP1_  (.D(_00680_),
    .Q(\count2_1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[4]$_SDFF_PP0_  (.D(_00681_),
    .Q(\count2_1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count2_1[5]$_SDFF_PP0_  (.D(_00682_),
    .Q(\count2_1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[1]$_SDFF_PP1_  (.D(_00683_),
    .Q(\count2_2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[2]$_SDFF_PP1_  (.D(_00684_),
    .Q(\count2_2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[3]$_SDFF_PP1_  (.D(_00685_),
    .Q(\count2_2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[4]$_SDFF_PP0_  (.D(_00686_),
    .Q(\count2_2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count2_2[5]$_SDFF_PP0_  (.D(_00687_),
    .Q(\count2_2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[1]$_SDFF_PP0_  (.D(_00688_),
    .Q(\count7_1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[2]$_SDFF_PP0_  (.D(_00689_),
    .Q(\count7_1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[3]$_SDFF_PP1_  (.D(_00690_),
    .Q(\count7_1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count7_1[4]$_SDFF_PP0_  (.D(_00691_),
    .Q(\count7_1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[5]$_SDFF_PP0_  (.D(_00692_),
    .Q(\count7_1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[1]$_SDFF_PP1_  (.D(_00693_),
    .Q(\count7_2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[2]$_SDFF_PP0_  (.D(_00694_),
    .Q(\count7_2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[3]$_SDFF_PP1_  (.D(_00695_),
    .Q(\count7_2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count7_2[4]$_SDFF_PP0_  (.D(_00696_),
    .Q(\count7_2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \count7_2[5]$_SDFF_PP0_  (.D(_00697_),
    .Q(\count7_2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[1]$_SDFFE_PP0N_  (.D(_00698_),
    .Q(\count_1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[2]$_SDFFE_PP0N_  (.D(_00699_),
    .Q(\count_1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[3]$_SDFFE_PP0N_  (.D(_00700_),
    .Q(\count_1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[4]$_SDFFE_PP1N_  (.D(_00701_),
    .Q(\count_1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[5]$_SDFFE_PP0N_  (.D(_00702_),
    .Q(\count_1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[1]$_SDFFE_PP0N_  (.D(_00703_),
    .Q(\count_2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[2]$_SDFFE_PP0N_  (.D(_00704_),
    .Q(\count_2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[3]$_SDFFE_PP0N_  (.D(_00705_),
    .Q(\count_2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[4]$_SDFFE_PP1N_  (.D(_00706_),
    .Q(\count_2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[5]$_SDFFE_PP0N_  (.D(_00707_),
    .Q(\count_2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[6]$_SDFFE_PP0N_  (.D(_00708_),
    .Q(\count_2[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash1[1]$_SDFFE_PP0N_  (.D(_00709_),
    .Q(\count_hash1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[2]$_SDFFE_PP0N_  (.D(_00710_),
    .Q(\count_hash1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[3]$_SDFFE_PP0N_  (.D(_00711_),
    .Q(\count_hash1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[4]$_SDFFE_PP0N_  (.D(_00712_),
    .Q(\count_hash1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[5]$_SDFFE_PP0N_  (.D(_00713_),
    .Q(\count_hash1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[6]$_SDFFE_PP0N_  (.D(_00714_),
    .Q(\count_hash1[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash2[1]$_SDFFE_PP0N_  (.D(_00715_),
    .Q(\count_hash2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[2]$_SDFFE_PP0N_  (.D(_00716_),
    .Q(\count_hash2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[3]$_SDFFE_PP0N_  (.D(_00717_),
    .Q(\count_hash2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[4]$_SDFFE_PP0N_  (.D(_00718_),
    .Q(\count_hash2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[5]$_SDFFE_PP0N_  (.D(_00719_),
    .Q(\count_hash2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \done$_DFFE_PN_  (.D(_00128_),
    .DE(_05334_),
    .Q(done),
    .CLK(clk));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_00_  (.A(\hash/a[13] ),
    .B(\hash/a[2] ),
    .C(\hash/a[22] ),
    .X(\hash/CA1/s0[0] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_01_  (.A(\hash/a[23] ),
    .B(\hash/a[12] ),
    .C(\hash/a[0] ),
    .X(\hash/CA1/s0[10] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_02_  (.A(\hash/a[13] ),
    .B(\hash/a[24] ),
    .C(\hash/a[1] ),
    .X(\hash/CA1/s0[11] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_03_  (.A(\hash/a[2] ),
    .B(\hash/a[14] ),
    .C(\hash/a[25] ),
    .X(\hash/CA1/s0[12] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_04_  (.A(\hash/a[3] ),
    .B(\hash/a[15] ),
    .C(\hash/a[26] ),
    .X(\hash/CA1/s0[13] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_05_  (.A(\hash/a[4] ),
    .B(\hash/a[16] ),
    .C(\hash/a[27] ),
    .X(\hash/CA1/s0[14] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_06_  (.A(\hash/a[5] ),
    .B(\hash/a[17] ),
    .C(\hash/a[28] ),
    .X(\hash/CA1/s0[15] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_07_  (.A(\hash/a[6] ),
    .B(\hash/a[18] ),
    .C(\hash/a[29] ),
    .X(\hash/CA1/s0[16] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_08_  (.A(\hash/a[7] ),
    .B(\hash/a[19] ),
    .C(\hash/a[30] ),
    .X(\hash/CA1/s0[17] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_09_  (.A(\hash/a[8] ),
    .B(\hash/a[20] ),
    .C(\hash/a[31] ),
    .X(\hash/CA1/s0[18] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_10_  (.A(\hash/a[9] ),
    .B(\hash/a[21] ),
    .C(\hash/a[0] ),
    .X(\hash/CA1/s0[19] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_11_  (.A(\hash/a[14] ),
    .B(\hash/a[3] ),
    .C(\hash/a[23] ),
    .X(\hash/CA1/s0[1] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_12_  (.A(\hash/a[10] ),
    .B(\hash/a[22] ),
    .C(\hash/a[1] ),
    .X(\hash/CA1/s0[20] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_13_  (.A(\hash/a[2] ),
    .B(\hash/a[11] ),
    .C(\hash/a[23] ),
    .X(\hash/CA1/s0[21] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_14_  (.A(\hash/a[3] ),
    .B(\hash/a[12] ),
    .C(\hash/a[24] ),
    .X(\hash/CA1/s0[22] ));
 sky130_fd_sc_hd__xor3_4 \hash/CA1/S0/_15_  (.A(\hash/a[13] ),
    .B(\hash/a[4] ),
    .C(\hash/a[25] ),
    .X(\hash/CA1/s0[23] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_16_  (.A(\hash/a[14] ),
    .B(\hash/a[5] ),
    .C(\hash/a[26] ),
    .X(\hash/CA1/s0[24] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_17_  (.A(\hash/a[15] ),
    .B(\hash/a[6] ),
    .C(\hash/a[27] ),
    .X(\hash/CA1/s0[25] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_18_  (.A(\hash/a[16] ),
    .B(\hash/a[7] ),
    .C(\hash/a[28] ),
    .X(\hash/CA1/s0[26] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_19_  (.A(\hash/a[17] ),
    .B(\hash/a[8] ),
    .C(\hash/a[29] ),
    .X(\hash/CA1/s0[27] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_20_  (.A(\hash/a[18] ),
    .B(\hash/a[9] ),
    .C(\hash/a[30] ),
    .X(\hash/CA1/s0[28] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_21_  (.A(\hash/a[19] ),
    .B(\hash/a[10] ),
    .C(\hash/a[31] ),
    .X(\hash/CA1/s0[29] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_22_  (.A(\hash/a[15] ),
    .B(\hash/a[4] ),
    .C(\hash/a[24] ),
    .X(\hash/CA1/s0[2] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_23_  (.A(\hash/a[20] ),
    .B(\hash/a[11] ),
    .C(\hash/a[0] ),
    .X(\hash/CA1/s0[30] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_24_  (.A(\hash/a[21] ),
    .B(\hash/a[12] ),
    .C(\hash/a[1] ),
    .X(\hash/CA1/s0[31] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_25_  (.A(\hash/a[16] ),
    .B(\hash/a[5] ),
    .C(\hash/a[25] ),
    .X(\hash/CA1/s0[3] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_26_  (.A(\hash/a[17] ),
    .B(\hash/a[6] ),
    .C(\hash/a[26] ),
    .X(\hash/CA1/s0[4] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_27_  (.A(\hash/a[18] ),
    .B(\hash/a[7] ),
    .C(\hash/a[27] ),
    .X(\hash/CA1/s0[5] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_28_  (.A(\hash/a[19] ),
    .B(\hash/a[8] ),
    .C(\hash/a[28] ),
    .X(\hash/CA1/s0[6] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_29_  (.A(\hash/a[20] ),
    .B(\hash/a[9] ),
    .C(\hash/a[29] ),
    .X(\hash/CA1/s0[7] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_30_  (.A(\hash/a[21] ),
    .B(\hash/a[10] ),
    .C(\hash/a[30] ),
    .X(\hash/CA1/s0[8] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S0/_31_  (.A(\hash/a[22] ),
    .B(\hash/a[11] ),
    .C(\hash/a[31] ),
    .X(\hash/CA1/s0[9] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_00_  (.A(\hash/e[11] ),
    .B(\hash/e[6] ),
    .C(\hash/e[25] ),
    .X(\hash/CA1/s1[0] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_01_  (.A(\hash/e[16] ),
    .B(\hash/e[21] ),
    .C(\hash/e[3] ),
    .X(\hash/CA1/s1[10] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_02_  (.A(\hash/e[17] ),
    .B(\hash/e[22] ),
    .C(\hash/e[4] ),
    .X(\hash/CA1/s1[11] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_03_  (.A(\hash/e[18] ),
    .B(\hash/e[23] ),
    .C(\hash/e[5] ),
    .X(\hash/CA1/s1[12] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_04_  (.A(\hash/e[6] ),
    .B(\hash/e[19] ),
    .C(\hash/e[24] ),
    .X(\hash/CA1/s1[13] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_05_  (.A(\hash/e[7] ),
    .B(\hash/e[20] ),
    .C(\hash/e[25] ),
    .X(\hash/CA1/s1[14] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_06_  (.A(\hash/e[8] ),
    .B(\hash/e[21] ),
    .C(\hash/e[26] ),
    .X(\hash/CA1/s1[15] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_07_  (.A(\hash/e[9] ),
    .B(\hash/e[22] ),
    .C(\hash/e[27] ),
    .X(\hash/CA1/s1[16] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_08_  (.A(\hash/e[10] ),
    .B(\hash/e[23] ),
    .C(\hash/e[28] ),
    .X(\hash/CA1/s1[17] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_09_  (.A(\hash/e[11] ),
    .B(\hash/e[24] ),
    .C(\hash/e[29] ),
    .X(\hash/CA1/s1[18] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_10_  (.A(\hash/e[12] ),
    .B(\hash/e[25] ),
    .C(\hash/e[30] ),
    .X(\hash/CA1/s1[19] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_11_  (.A(\hash/e[12] ),
    .B(\hash/e[7] ),
    .C(\hash/e[26] ),
    .X(\hash/CA1/s1[1] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_12_  (.A(\hash/e[13] ),
    .B(\hash/e[26] ),
    .C(\hash/e[31] ),
    .X(\hash/CA1/s1[20] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_13_  (.A(\hash/e[14] ),
    .B(\hash/e[27] ),
    .C(\hash/e[0] ),
    .X(\hash/CA1/s1[21] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_14_  (.A(\hash/e[15] ),
    .B(\hash/e[28] ),
    .C(\hash/e[1] ),
    .X(\hash/CA1/s1[22] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_15_  (.A(\hash/e[16] ),
    .B(\hash/e[29] ),
    .C(\hash/e[2] ),
    .X(\hash/CA1/s1[23] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_16_  (.A(\hash/e[17] ),
    .B(\hash/e[30] ),
    .C(\hash/e[3] ),
    .X(\hash/CA1/s1[24] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_17_  (.A(\hash/e[18] ),
    .B(\hash/e[31] ),
    .C(\hash/e[4] ),
    .X(\hash/CA1/s1[25] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_18_  (.A(\hash/e[19] ),
    .B(\hash/e[0] ),
    .C(\hash/e[5] ),
    .X(\hash/CA1/s1[26] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_19_  (.A(\hash/e[6] ),
    .B(\hash/e[20] ),
    .C(\hash/e[1] ),
    .X(\hash/CA1/s1[27] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_20_  (.A(\hash/e[7] ),
    .B(\hash/e[21] ),
    .C(\hash/e[2] ),
    .X(\hash/CA1/s1[28] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_21_  (.A(\hash/e[8] ),
    .B(\hash/e[22] ),
    .C(\hash/e[3] ),
    .X(\hash/CA1/s1[29] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_22_  (.A(\hash/e[13] ),
    .B(\hash/e[8] ),
    .C(\hash/e[27] ),
    .X(\hash/CA1/s1[2] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_23_  (.A(\hash/e[9] ),
    .B(\hash/e[23] ),
    .C(\hash/e[4] ),
    .X(\hash/CA1/s1[30] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_24_  (.A(\hash/e[10] ),
    .B(\hash/e[24] ),
    .C(\hash/e[5] ),
    .X(\hash/CA1/s1[31] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_25_  (.A(\hash/e[14] ),
    .B(\hash/e[9] ),
    .C(\hash/e[28] ),
    .X(\hash/CA1/s1[3] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_26_  (.A(\hash/e[15] ),
    .B(\hash/e[10] ),
    .C(\hash/e[29] ),
    .X(\hash/CA1/s1[4] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_27_  (.A(\hash/e[11] ),
    .B(\hash/e[16] ),
    .C(\hash/e[30] ),
    .X(\hash/CA1/s1[5] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_28_  (.A(\hash/e[12] ),
    .B(\hash/e[17] ),
    .C(\hash/e[31] ),
    .X(\hash/CA1/s1[6] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_29_  (.A(\hash/e[13] ),
    .B(\hash/e[18] ),
    .C(\hash/e[0] ),
    .X(\hash/CA1/s1[7] ));
 sky130_fd_sc_hd__xor3_4 \hash/CA1/S1/_30_  (.A(\hash/e[14] ),
    .B(\hash/e[19] ),
    .C(\hash/e[1] ),
    .X(\hash/CA1/s1[8] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA1/S1/_31_  (.A(\hash/e[15] ),
    .B(\hash/e[20] ),
    .C(\hash/e[2] ),
    .X(\hash/CA1/s1[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_1977_  (.A0(\hash/g[0] ),
    .A1(\hash/f[0] ),
    .S(\hash/e[0] ),
    .X(\hash/CA1/_1640_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA1/_1978_  (.A0(\hash/g[1] ),
    .A1(\hash/f[1] ),
    .S(\hash/e[1] ),
    .Y(\hash/CA1/_1060_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_1979_  (.A(\hash/CA1/_1060_ ),
    .Y(\hash/CA1/_1645_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_1980_  (.A(\hash/CA1/_1057_ ),
    .B(\hash/CA1/_1649_ ),
    .Y(\hash/CA1/_1068_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_1981_  (.A(\hash/CA1/_1068_ ),
    .Y(\hash/CA1/_1226_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_1982_  (.A0(\hash/g[2] ),
    .A1(\hash/f[2] ),
    .S(\hash/e[2] ),
    .X(\hash/CA1/_1650_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_1983_  (.A1(\hash/CA1/_1638_ ),
    .A2(\hash/CA1/_1644_ ),
    .B1(\hash/CA1/_1643_ ),
    .X(\hash/CA1/_0000_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_1984_  (.A1(\hash/CA1/_1649_ ),
    .A2(\hash/CA1/_0000_ ),
    .B1(\hash/CA1/_1648_ ),
    .Y(\hash/CA1/_0001_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_1985_  (.A(\hash/CA1/_1656_ ),
    .B(\hash/CA1/_0001_ ),
    .Y(\hash/CA1/_1073_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_1986_  (.A(\hash/CA1/_1073_ ),
    .Y(\hash/CA1/_1235_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_1987_  (.A0(\hash/g[3] ),
    .A1(\hash/f[3] ),
    .S(\hash/e[3] ),
    .X(\hash/CA1/_1657_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_1988_  (.A(\hash/CA1/_1057_ ),
    .B_N(\hash/CA1/_1649_ ),
    .Y(\hash/CA1/_0002_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_1989_  (.A1(\hash/CA1/_1648_ ),
    .A2(\hash/CA1/_0002_ ),
    .B1(\hash/CA1/_1656_ ),
    .Y(\hash/CA1/_0003_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_1990_  (.A_N(\hash/CA1/_1655_ ),
    .B(\hash/CA1/_0003_ ),
    .Y(\hash/CA1/_0004_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_1991_  (.A(\hash/CA1/_1663_ ),
    .B(\hash/CA1/_0004_ ),
    .Y(\hash/CA1/_1077_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_1992_  (.A(\hash/CA1/_1077_ ),
    .Y(\hash/CA1/_1242_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_1993_  (.A0(\hash/g[4] ),
    .A1(\hash/f[4] ),
    .S(\hash/e[4] ),
    .X(\hash/CA1/_1664_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_1994_  (.A(\hash/CA1/_1062_ ),
    .B_N(\hash/CA1/_1652_ ),
    .Y(\hash/CA1/_0005_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_1995_  (.A1(\hash/CA1/_1651_ ),
    .A2(\hash/CA1/_0005_ ),
    .B1(\hash/CA1/_1659_ ),
    .X(\hash/CA1/_0006_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_1996_  (.A(\hash/CA1/_1658_ ),
    .B(\hash/CA1/_0006_ ),
    .X(\hash/CA1/_0007_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_1997_  (.A(\hash/CA1/_1666_ ),
    .B(\hash/CA1/_0007_ ),
    .X(\hash/CA1/_1245_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_1998_  (.A(\hash/CA1/_1245_ ),
    .Y(\hash/CA1/_1078_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_1999_  (.A0(\hash/g[5] ),
    .A1(\hash/f[5] ),
    .S(\hash/e[5] ),
    .X(\hash/CA1/_1672_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2000_  (.A1(\hash/CA1/_1641_ ),
    .A2(\hash/CA1/_1647_ ),
    .B1(\hash/CA1/_1646_ ),
    .C1(\hash/CA1/_1651_ ),
    .Y(\hash/CA1/_0008_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_2001_  (.A1(\hash/CA1/_1652_ ),
    .A2(\hash/CA1/_1651_ ),
    .B1(\hash/CA1/_1666_ ),
    .C1(\hash/CA1/_1659_ ),
    .Y(\hash/CA1/_0009_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2002_  (.A1(\hash/CA1/_1666_ ),
    .A2(\hash/CA1/_1658_ ),
    .B1(\hash/CA1/_1665_ ),
    .Y(\hash/CA1/_0010_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2003_  (.A1(\hash/CA1/_0008_ ),
    .A2(\hash/CA1/_0009_ ),
    .B1(\hash/CA1/_0010_ ),
    .Y(\hash/CA1/_0011_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2004_  (.A(\hash/CA1/_1674_ ),
    .B(\hash/CA1/_0011_ ),
    .X(\hash/CA1/_1081_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2005_  (.A(\hash/CA1/_1081_ ),
    .Y(\hash/CA1/_1251_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2006_  (.A0(\hash/g[6] ),
    .A1(\hash/f[6] ),
    .S(\hash/e[6] ),
    .X(\hash/CA1/_1680_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_2007_  (.A1(\hash/CA1/_1658_ ),
    .A2(\hash/CA1/_0006_ ),
    .B1(\hash/CA1/_1666_ ),
    .Y(\hash/CA1/_0012_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2008_  (.A_N(\hash/CA1/_1665_ ),
    .B(\hash/CA1/_0012_ ),
    .Y(\hash/CA1/_0013_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2009_  (.A1(\hash/CA1/_1674_ ),
    .A2(\hash/CA1/_0013_ ),
    .B1(\hash/CA1/_1673_ ),
    .Y(\hash/CA1/_0014_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2010_  (.A(\hash/CA1/_1682_ ),
    .B(\hash/CA1/_0014_ ),
    .Y(\hash/CA1/_1085_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2011_  (.A(\hash/CA1/_1085_ ),
    .Y(\hash/CA1/_1258_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2012_  (.A0(\hash/g[7] ),
    .A1(\hash/f[7] ),
    .S(\hash/e[7] ),
    .X(\hash/CA1/_1687_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2013_  (.A(\hash/CA1/_1681_ ),
    .Y(\hash/CA1/_0015_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2014_  (.A1(\hash/CA1/_1674_ ),
    .A2(\hash/CA1/_1673_ ),
    .B1(\hash/CA1/_1682_ ),
    .Y(\hash/CA1/_0016_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2015_  (.A(\hash/CA1/_0015_ ),
    .B(\hash/CA1/_0016_ ),
    .Y(\hash/CA1/_0017_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2016_  (.A(\hash/CA1/_1673_ ),
    .B(\hash/CA1/_1681_ ),
    .Y(\hash/CA1/_0018_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_2017_  (.A1(\hash/CA1/_0008_ ),
    .A2(\hash/CA1/_0009_ ),
    .B1(\hash/CA1/_0010_ ),
    .C1(\hash/CA1/_0018_ ),
    .Y(\hash/CA1/_0019_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2018_  (.A(\hash/CA1/_0017_ ),
    .B(\hash/CA1/_0019_ ),
    .Y(\hash/CA1/_0020_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2019_  (.A(\hash/CA1/_1689_ ),
    .B(\hash/CA1/_0020_ ),
    .Y(\hash/CA1/_1089_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2020_  (.A(\hash/CA1/_1089_ ),
    .Y(\hash/CA1/_1265_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2021_  (.A(\hash/CA1/_1656_ ),
    .B(\hash/CA1/_1663_ ),
    .Y(\hash/CA1/_0021_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2022_  (.A1(\hash/CA1/_1648_ ),
    .A2(\hash/CA1/_0002_ ),
    .B1_N(\hash/CA1/_0021_ ),
    .Y(\hash/CA1/_0022_ ));
 sky130_fd_sc_hd__a2111oi_2 \hash/CA1/_2023_  (.A1(\hash/CA1/_1663_ ),
    .A2(\hash/CA1/_1655_ ),
    .B1(\hash/CA1/_1662_ ),
    .C1(\hash/CA1/_1670_ ),
    .D1(\hash/CA1/_1678_ ),
    .Y(\hash/CA1/_0023_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2024_  (.A1(\hash/CA1/_1671_ ),
    .A2(\hash/CA1/_1670_ ),
    .B1(\hash/CA1/_1679_ ),
    .X(\hash/CA1/_0024_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2025_  (.A1(\hash/CA1/_1678_ ),
    .A2(\hash/CA1/_0024_ ),
    .B1(\hash/CA1/_1686_ ),
    .Y(\hash/CA1/_0025_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2026_  (.A1(\hash/CA1/_0022_ ),
    .A2(\hash/CA1/_0023_ ),
    .B1(\hash/CA1/_0025_ ),
    .Y(\hash/CA1/_0026_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2027_  (.A(\hash/CA1/_1685_ ),
    .B(\hash/CA1/_0026_ ),
    .Y(\hash/CA1/_0027_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2028_  (.A(\hash/CA1/_1693_ ),
    .B(\hash/CA1/_0027_ ),
    .Y(\hash/CA1/_1093_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2029_  (.A(\hash/CA1/_1093_ ),
    .Y(\hash/CA1/_1097_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2030_  (.A0(\hash/g[8] ),
    .A1(\hash/f[8] ),
    .S(\hash/e[8] ),
    .X(\hash/CA1/_1694_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_2031_  (.A(\hash/CA1/_1678_ ),
    .B(\hash/CA1/_0024_ ),
    .X(\hash/CA1/_0028_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2032_  (.A1(\hash/CA1/_1638_ ),
    .A2(\hash/CA1/_1644_ ),
    .B1(\hash/CA1/_1643_ ),
    .C1(\hash/CA1/_1648_ ),
    .Y(\hash/CA1/_0029_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2033_  (.A(\hash/CA1/_1649_ ),
    .B(\hash/CA1/_1648_ ),
    .Y(\hash/CA1/_0030_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2034_  (.A1(\hash/CA1/_0021_ ),
    .A2(\hash/CA1/_0029_ ),
    .A3(\hash/CA1/_0030_ ),
    .B1(\hash/CA1/_0023_ ),
    .Y(\hash/CA1/_0031_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2035_  (.A1(\hash/CA1/_1693_ ),
    .A2(\hash/CA1/_1685_ ),
    .B1(\hash/CA1/_1692_ ),
    .X(\hash/CA1/_0032_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/CA1/_2036_  (.A1(\hash/CA1/_1686_ ),
    .A2(\hash/CA1/_1693_ ),
    .A3(\hash/CA1/_0028_ ),
    .A4(\hash/CA1/_0031_ ),
    .B1(\hash/CA1/_0032_ ),
    .Y(\hash/CA1/_0033_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2037_  (.A(\hash/CA1/_1700_ ),
    .B(\hash/CA1/_0033_ ),
    .X(\hash/CA1/_1100_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2038_  (.A(\hash/CA1/_1100_ ),
    .Y(\hash/CA1/_1276_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2039_  (.A0(\hash/g[9] ),
    .A1(\hash/f[9] ),
    .S(\hash/e[9] ),
    .X(\hash/CA1/_1701_ ));
 sky130_fd_sc_hd__a31o_2 \hash/CA1/_2040_  (.A1(\hash/CA1/_1689_ ),
    .A2(\hash/CA1/_0017_ ),
    .A3(\hash/CA1/_0019_ ),
    .B1(\hash/CA1/_1688_ ),
    .X(\hash/CA1/_0034_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2041_  (.A1(\hash/CA1/_1696_ ),
    .A2(\hash/CA1/_0034_ ),
    .B1(\hash/CA1/_1695_ ),
    .Y(\hash/CA1/_0035_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2042_  (.A(\hash/CA1/_1703_ ),
    .B(\hash/CA1/_0035_ ),
    .X(\hash/CA1/_1101_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2043_  (.A1(\hash/CA1/_1685_ ),
    .A2(\hash/CA1/_0026_ ),
    .B1(\hash/CA1/_1693_ ),
    .Y(\hash/CA1/_0036_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2044_  (.A_N(\hash/CA1/_1692_ ),
    .B(\hash/CA1/_0036_ ),
    .Y(\hash/CA1/_0037_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2045_  (.A1(\hash/CA1/_1700_ ),
    .A2(\hash/CA1/_0037_ ),
    .B1(\hash/CA1/_1699_ ),
    .Y(\hash/CA1/_0038_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2046_  (.A(\hash/CA1/_1708_ ),
    .B(\hash/CA1/_0038_ ),
    .X(\hash/CA1/_1105_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2047_  (.A(\hash/CA1/_1105_ ),
    .Y(\hash/CA1/_1282_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2048_  (.A0(\hash/g[10] ),
    .A1(\hash/f[10] ),
    .S(\hash/e[10] ),
    .X(\hash/CA1/_1709_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2049_  (.A(\hash/CA1/_1711_ ),
    .Y(\hash/CA1/_0039_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2050_  (.A(\hash/CA1/_1688_ ),
    .B(\hash/CA1/_1695_ ),
    .Y(\hash/CA1/_0040_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2051_  (.A(\hash/CA1/_0018_ ),
    .B(\hash/CA1/_0040_ ),
    .Y(\hash/CA1/_0041_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2052_  (.A(\hash/CA1/_1665_ ),
    .B(\hash/CA1/_0041_ ),
    .Y(\hash/CA1/_0042_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2053_  (.A1(\hash/CA1/_1682_ ),
    .A2(\hash/CA1/_1681_ ),
    .B1(\hash/CA1/_1689_ ),
    .X(\hash/CA1/_0043_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2054_  (.A1(\hash/CA1/_1688_ ),
    .A2(\hash/CA1/_0043_ ),
    .B1(\hash/CA1/_1696_ ),
    .X(\hash/CA1/_0044_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA1/_2055_  (.A1(\hash/CA1/_1695_ ),
    .A2(\hash/CA1/_0044_ ),
    .B1(\hash/CA1/_0041_ ),
    .B2(\hash/CA1/_1674_ ),
    .Y(\hash/CA1/_0045_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2056_  (.A1(\hash/CA1/_0012_ ),
    .A2(\hash/CA1/_0042_ ),
    .B1(\hash/CA1/_0045_ ),
    .Y(\hash/CA1/_0046_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2057_  (.A1(\hash/CA1/_1703_ ),
    .A2(\hash/CA1/_0046_ ),
    .B1(\hash/CA1/_1702_ ),
    .Y(\hash/CA1/_0047_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2058_  (.A(\hash/CA1/_0039_ ),
    .B(\hash/CA1/_0047_ ),
    .Y(\hash/CA1/_1106_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2059_  (.A1(\hash/CA1/_1708_ ),
    .A2(\hash/CA1/_1699_ ),
    .B1(\hash/CA1/_1707_ ),
    .X(\hash/CA1/_0048_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2060_  (.A(\hash/CA1/_1700_ ),
    .B(\hash/CA1/_1708_ ),
    .Y(\hash/CA1/_0049_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2061_  (.A(\hash/CA1/_0033_ ),
    .B(\hash/CA1/_0049_ ),
    .Y(\hash/CA1/_0050_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_2062_  (.A(\hash/CA1/_0048_ ),
    .B(\hash/CA1/_0050_ ),
    .X(\hash/CA1/_0051_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2063_  (.A(\hash/CA1/_1717_ ),
    .B(\hash/CA1/_0051_ ),
    .Y(\hash/CA1/_1110_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2064_  (.A(\hash/CA1/_1110_ ),
    .Y(\hash/CA1/_1289_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2065_  (.A0(\hash/g[11] ),
    .A1(\hash/f[11] ),
    .S(\hash/e[11] ),
    .X(\hash/CA1/_1718_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2066_  (.A(\hash/CA1/_1720_ ),
    .Y(\hash/CA1/_0052_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2067_  (.A(\hash/CA1/_1689_ ),
    .B(\hash/CA1/_1696_ ),
    .C(\hash/CA1/_1703_ ),
    .D(\hash/CA1/_1711_ ),
    .Y(\hash/CA1/_0053_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2068_  (.A1(\hash/CA1/_0015_ ),
    .A2(\hash/CA1/_0016_ ),
    .B1(\hash/CA1/_0053_ ),
    .Y(\hash/CA1/_0054_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2069_  (.A(\hash/CA1/_1703_ ),
    .B(\hash/CA1/_1711_ ),
    .Y(\hash/CA1/_0055_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2070_  (.A1(\hash/CA1/_1696_ ),
    .A2(\hash/CA1/_1688_ ),
    .B1(\hash/CA1/_1695_ ),
    .Y(\hash/CA1/_0056_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2071_  (.A1(\hash/CA1/_1711_ ),
    .A2(\hash/CA1/_1702_ ),
    .B1(\hash/CA1/_1710_ ),
    .Y(\hash/CA1/_0057_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2072_  (.A1(\hash/CA1/_0055_ ),
    .A2(\hash/CA1/_0056_ ),
    .B1(\hash/CA1/_0057_ ),
    .Y(\hash/CA1/_0058_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2073_  (.A1(\hash/CA1/_0019_ ),
    .A2(\hash/CA1/_0054_ ),
    .B1(\hash/CA1/_0058_ ),
    .Y(\hash/CA1/_0059_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2074_  (.A(\hash/CA1/_0052_ ),
    .B(\hash/CA1/_0059_ ),
    .Y(\hash/CA1/_1111_ ));
 sky130_fd_sc_hd__o2111ai_1 \hash/CA1/_2075_  (.A1(\hash/CA1/_1685_ ),
    .A2(\hash/CA1/_0026_ ),
    .B1(\hash/CA1/_1693_ ),
    .C1(\hash/CA1/_1700_ ),
    .D1(\hash/CA1/_1708_ ),
    .Y(\hash/CA1/_0060_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2076_  (.A1(\hash/CA1/_1700_ ),
    .A2(\hash/CA1/_1692_ ),
    .B1(\hash/CA1/_1699_ ),
    .X(\hash/CA1/_0061_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2077_  (.A(\hash/CA1/_1708_ ),
    .B(\hash/CA1/_0061_ ),
    .Y(\hash/CA1/_0062_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2078_  (.A(\hash/CA1/_0060_ ),
    .B(\hash/CA1/_0062_ ),
    .Y(\hash/CA1/_0063_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2079_  (.A1(\hash/CA1/_1707_ ),
    .A2(\hash/CA1/_0063_ ),
    .B1(\hash/CA1/_1717_ ),
    .Y(\hash/CA1/_0064_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2080_  (.A(\hash/CA1/_1716_ ),
    .B_N(\hash/CA1/_0064_ ),
    .Y(\hash/CA1/_0065_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2081_  (.A(\hash/CA1/_1726_ ),
    .B(\hash/CA1/_0065_ ),
    .X(\hash/CA1/_1115_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2082_  (.A(\hash/CA1/_1115_ ),
    .Y(\hash/CA1/_1296_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2083_  (.A0(\hash/g[12] ),
    .A1(\hash/f[12] ),
    .S(\hash/e[12] ),
    .X(\hash/CA1/_1727_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2084_  (.A1(\hash/CA1/_0039_ ),
    .A2(\hash/CA1/_0047_ ),
    .B1_N(\hash/CA1/_1710_ ),
    .Y(\hash/CA1/_0066_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2085_  (.A1(\hash/CA1/_1720_ ),
    .A2(\hash/CA1/_0066_ ),
    .B1(\hash/CA1/_1719_ ),
    .Y(\hash/CA1/_0067_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2086_  (.A(\hash/CA1/_1729_ ),
    .B(\hash/CA1/_0067_ ),
    .X(\hash/CA1/_1116_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2087_  (.A1(\hash/CA1/_1717_ ),
    .A2(\hash/CA1/_0051_ ),
    .B1(\hash/CA1/_1716_ ),
    .X(\hash/CA1/_0068_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2088_  (.A1(\hash/CA1/_1726_ ),
    .A2(\hash/CA1/_0068_ ),
    .B1(\hash/CA1/_1725_ ),
    .X(\hash/CA1/_0069_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2089_  (.A(\hash/CA1/_1735_ ),
    .B(\hash/CA1/_0069_ ),
    .Y(\hash/CA1/_1120_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2090_  (.A(\hash/CA1/_1120_ ),
    .Y(\hash/CA1/_1303_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2091_  (.A0(\hash/g[13] ),
    .A1(\hash/f[13] ),
    .S(\hash/e[13] ),
    .X(\hash/CA1/_1736_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2092_  (.A1(\hash/CA1/_0052_ ),
    .A2(\hash/CA1/_0059_ ),
    .B1_N(\hash/CA1/_1719_ ),
    .Y(\hash/CA1/_0070_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2093_  (.A1(\hash/CA1/_1729_ ),
    .A2(\hash/CA1/_0070_ ),
    .B1(\hash/CA1/_1728_ ),
    .Y(\hash/CA1/_0071_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2094_  (.A(\hash/CA1/_1738_ ),
    .B(\hash/CA1/_0071_ ),
    .Y(\hash/CA1/_1306_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2095_  (.A(\hash/CA1/_1306_ ),
    .Y(\hash/CA1/_1121_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2097_  (.A(\hash/CA1/_1717_ ),
    .B(\hash/CA1/_1726_ ),
    .C(\hash/CA1/_1735_ ),
    .X(\hash/CA1/_0073_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2098_  (.A1(\hash/CA1/_1717_ ),
    .A2(\hash/CA1/_1707_ ),
    .B1(\hash/CA1/_1716_ ),
    .X(\hash/CA1/_0074_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2099_  (.A1(\hash/CA1/_1726_ ),
    .A2(\hash/CA1/_0074_ ),
    .B1(\hash/CA1/_1725_ ),
    .Y(\hash/CA1/_0075_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2100_  (.A(\hash/CA1/_0075_ ),
    .B_N(\hash/CA1/_1735_ ),
    .Y(\hash/CA1/_0076_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2101_  (.A1(\hash/CA1/_0063_ ),
    .A2(\hash/CA1/_0073_ ),
    .B1(\hash/CA1/_0076_ ),
    .Y(\hash/CA1/_0077_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2102_  (.A(\hash/CA1/_1734_ ),
    .B_N(\hash/CA1/_0077_ ),
    .Y(\hash/CA1/_0078_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2103_  (.A(\hash/CA1/_1744_ ),
    .B(\hash/CA1/_0078_ ),
    .X(\hash/CA1/_1126_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2104_  (.A(\hash/CA1/_1126_ ),
    .Y(\hash/CA1/_1309_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2105_  (.A0(\hash/g[14] ),
    .A1(\hash/f[14] ),
    .S(\hash/e[14] ),
    .X(\hash/CA1/_1745_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2106_  (.A(\hash/CA1/_1747_ ),
    .Y(\hash/CA1/_0079_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2107_  (.A(\hash/CA1/_1720_ ),
    .B(\hash/CA1/_1729_ ),
    .C(\hash/CA1/_1738_ ),
    .Y(\hash/CA1/_0080_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2108_  (.A(\hash/CA1/_0079_ ),
    .B(\hash/CA1/_0055_ ),
    .C(\hash/CA1/_0080_ ),
    .Y(\hash/CA1/_0081_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2109_  (.A1(\hash/CA1/_0052_ ),
    .A2(\hash/CA1/_0057_ ),
    .B1_N(\hash/CA1/_1719_ ),
    .Y(\hash/CA1/_0082_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2110_  (.A1(\hash/CA1/_1729_ ),
    .A2(\hash/CA1/_0082_ ),
    .B1(\hash/CA1/_1728_ ),
    .X(\hash/CA1/_0083_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2111_  (.A1(\hash/CA1/_1738_ ),
    .A2(\hash/CA1/_0083_ ),
    .B1(\hash/CA1/_1737_ ),
    .Y(\hash/CA1/_0084_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \hash/CA1/_2112_  (.A1_N(\hash/CA1/_0046_ ),
    .A2_N(\hash/CA1/_0081_ ),
    .B1(\hash/CA1/_0084_ ),
    .B2(\hash/CA1/_0079_ ),
    .Y(\hash/CA1/_0085_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2113_  (.A(\hash/CA1/_0055_ ),
    .B(\hash/CA1/_0080_ ),
    .Y(\hash/CA1/_0086_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2114_  (.A(\hash/CA1/_0079_ ),
    .B(\hash/CA1/_0084_ ),
    .Y(\hash/CA1/_0087_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2115_  (.A1(\hash/CA1/_0046_ ),
    .A2(\hash/CA1/_0086_ ),
    .B1(\hash/CA1/_0087_ ),
    .Y(\hash/CA1/_0088_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2116_  (.A(\hash/CA1/_0085_ ),
    .B(\hash/CA1/_0088_ ),
    .Y(\hash/CA1/_1312_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2117_  (.A(\hash/CA1/_1312_ ),
    .Y(\hash/CA1/_1125_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2119_  (.A(\hash/CA1/_1744_ ),
    .B(\hash/CA1/_0073_ ),
    .Y(\hash/CA1/_0090_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2120_  (.A1(\hash/CA1/_1726_ ),
    .A2(\hash/CA1/_1716_ ),
    .B1(\hash/CA1/_1725_ ),
    .X(\hash/CA1/_0091_ ));
 sky130_fd_sc_hd__a221o_1 \hash/CA1/_2121_  (.A1(\hash/CA1/_0048_ ),
    .A2(\hash/CA1/_0073_ ),
    .B1(\hash/CA1/_0091_ ),
    .B2(\hash/CA1/_1735_ ),
    .C1(\hash/CA1/_1734_ ),
    .X(\hash/CA1/_0092_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2122_  (.A1(\hash/CA1/_1744_ ),
    .A2(\hash/CA1/_0092_ ),
    .B1(\hash/CA1/_1743_ ),
    .Y(\hash/CA1/_0093_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2123_  (.A1(\hash/CA1/_0033_ ),
    .A2(\hash/CA1/_0049_ ),
    .A3(\hash/CA1/_0090_ ),
    .B1(\hash/CA1/_0093_ ),
    .Y(\hash/CA1/_0094_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2124_  (.A(\hash/CA1/_1753_ ),
    .B(\hash/CA1/_0094_ ),
    .X(\hash/CA1/_1130_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2125_  (.A(\hash/CA1/_1130_ ),
    .Y(\hash/CA1/_1133_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2126_  (.A0(\hash/g[15] ),
    .A1(\hash/f[15] ),
    .S(\hash/e[15] ),
    .X(\hash/CA1/_1754_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2127_  (.A1(\hash/CA1/_1744_ ),
    .A2(\hash/CA1/_1734_ ),
    .B1(\hash/CA1/_1743_ ),
    .X(\hash/CA1/_0095_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2128_  (.A1(\hash/CA1/_1753_ ),
    .A2(\hash/CA1/_0095_ ),
    .B1(\hash/CA1/_1752_ ),
    .Y(\hash/CA1/_0096_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2129_  (.A(\hash/CA1/_1744_ ),
    .B(\hash/CA1/_1753_ ),
    .C(\hash/CA1/_0076_ ),
    .Y(\hash/CA1/_0097_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA1/_2130_  (.A1(\hash/CA1/_0096_ ),
    .A2(\hash/CA1/_0097_ ),
    .B1_N(\hash/CA1/_1761_ ),
    .Y(\hash/CA1/_0098_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2131_  (.A(\hash/CA1/_1744_ ),
    .B(\hash/CA1/_1753_ ),
    .C(\hash/CA1/_1761_ ),
    .D(\hash/CA1/_0073_ ),
    .Y(\hash/CA1/_0099_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2132_  (.A1(\hash/CA1/_0060_ ),
    .A2(\hash/CA1/_0062_ ),
    .B1(\hash/CA1/_0099_ ),
    .Y(\hash/CA1/_0100_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2133_  (.A(\hash/CA1/_0098_ ),
    .B(\hash/CA1/_0100_ ),
    .Y(\hash/CA1/_0101_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2134_  (.A(\hash/CA1/_1744_ ),
    .B(\hash/CA1/_1753_ ),
    .Y(\hash/CA1/_0102_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2135_  (.A(\hash/CA1/_1761_ ),
    .B_N(\hash/CA1/_0096_ ),
    .Y(\hash/CA1/_0103_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2136_  (.A1(\hash/CA1/_0077_ ),
    .A2(\hash/CA1/_0102_ ),
    .B1(\hash/CA1/_0103_ ),
    .Y(\hash/CA1/_0104_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2137_  (.A(\hash/CA1/_0101_ ),
    .B(\hash/CA1/_0104_ ),
    .Y(\hash/CA1/_1136_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2138_  (.A(\hash/CA1/_1136_ ),
    .Y(\hash/CA1/_1321_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2139_  (.A0(\hash/g[16] ),
    .A1(\hash/f[16] ),
    .S(\hash/e[16] ),
    .X(\hash/CA1/_1762_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2140_  (.A1(\hash/CA1/_1746_ ),
    .A2(\hash/CA1/_0085_ ),
    .B1(\hash/CA1/_1756_ ),
    .X(\hash/CA1/_0105_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2141_  (.A(\hash/CA1/_1755_ ),
    .B(\hash/CA1/_0105_ ),
    .Y(\hash/CA1/_0106_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2142_  (.A(\hash/CA1/_1764_ ),
    .B(\hash/CA1/_0106_ ),
    .X(\hash/CA1/_1137_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2143_  (.A1(\hash/CA1/_1761_ ),
    .A2(\hash/CA1/_1752_ ),
    .B1(\hash/CA1/_1760_ ),
    .Y(\hash/CA1/_0107_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2144_  (.A(\hash/CA1/_1753_ ),
    .B(\hash/CA1/_1761_ ),
    .C(\hash/CA1/_0094_ ),
    .Y(\hash/CA1/_0108_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2145_  (.A(\hash/CA1/_0107_ ),
    .B(\hash/CA1/_0108_ ),
    .Y(\hash/CA1/_0109_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2146_  (.A(\hash/CA1/_1769_ ),
    .B(\hash/CA1/_0109_ ),
    .Y(\hash/CA1/_1142_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2147_  (.A(\hash/CA1/_1142_ ),
    .Y(\hash/CA1/_1327_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2148_  (.A0(\hash/g[17] ),
    .A1(\hash/f[17] ),
    .S(\hash/e[17] ),
    .X(\hash/CA1/_1770_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2149_  (.A(\hash/CA1/_0079_ ),
    .B(\hash/CA1/_0059_ ),
    .C(\hash/CA1/_0080_ ),
    .Y(\hash/CA1/_0110_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2150_  (.A1(\hash/CA1/_1729_ ),
    .A2(\hash/CA1/_1719_ ),
    .B1(\hash/CA1/_1728_ ),
    .Y(\hash/CA1/_0111_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2151_  (.A(\hash/CA1/_1738_ ),
    .B(\hash/CA1/_1747_ ),
    .Y(\hash/CA1/_0112_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2152_  (.A1(\hash/CA1/_1747_ ),
    .A2(\hash/CA1/_1737_ ),
    .B1(\hash/CA1/_1746_ ),
    .Y(\hash/CA1/_0113_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2153_  (.A1(\hash/CA1/_0111_ ),
    .A2(\hash/CA1/_0112_ ),
    .B1(\hash/CA1/_0113_ ),
    .Y(\hash/CA1/_0114_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2154_  (.A(\hash/CA1/_0110_ ),
    .B(\hash/CA1/_0114_ ),
    .Y(\hash/CA1/_0115_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2155_  (.A(\hash/CA1/_1756_ ),
    .B(\hash/CA1/_1764_ ),
    .Y(\hash/CA1/_0116_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2156_  (.A1(\hash/CA1/_1764_ ),
    .A2(\hash/CA1/_1755_ ),
    .B1(\hash/CA1/_1763_ ),
    .X(\hash/CA1/_0117_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2157_  (.A1(\hash/CA1/_0115_ ),
    .A2(\hash/CA1/_0116_ ),
    .B1_N(\hash/CA1/_0117_ ),
    .Y(\hash/CA1/_0118_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2158_  (.A(\hash/CA1/_1772_ ),
    .B(\hash/CA1/_0118_ ),
    .X(\hash/CA1/_1330_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2159_  (.A(\hash/CA1/_1330_ ),
    .Y(\hash/CA1/_1141_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2161_  (.A(\hash/CA1/_1769_ ),
    .Y(\hash/CA1/_0120_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2162_  (.A(\hash/CA1/_1760_ ),
    .B(\hash/CA1/_0098_ ),
    .C(\hash/CA1/_0100_ ),
    .Y(\hash/CA1/_0121_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2163_  (.A1(\hash/CA1/_0120_ ),
    .A2(\hash/CA1/_0121_ ),
    .B1_N(\hash/CA1/_1768_ ),
    .Y(\hash/CA1/_0122_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2164_  (.A(\hash/CA1/_1778_ ),
    .B(\hash/CA1/_0122_ ),
    .Y(\hash/CA1/_1146_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2165_  (.A(\hash/CA1/_1146_ ),
    .Y(\hash/CA1/_1333_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2166_  (.A0(\hash/g[18] ),
    .A1(\hash/f[18] ),
    .S(\hash/e[18] ),
    .X(\hash/CA1/_1779_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2167_  (.A1(\hash/CA1/_1756_ ),
    .A2(\hash/CA1/_1746_ ),
    .B1(\hash/CA1/_1755_ ),
    .X(\hash/CA1/_0123_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2168_  (.A1(\hash/CA1/_1764_ ),
    .A2(\hash/CA1/_0123_ ),
    .B1(\hash/CA1/_1763_ ),
    .Y(\hash/CA1/_0124_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2169_  (.A(\hash/CA1/_1756_ ),
    .B(\hash/CA1/_1764_ ),
    .C(\hash/CA1/_0085_ ),
    .Y(\hash/CA1/_0125_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2170_  (.A(\hash/CA1/_0124_ ),
    .B(\hash/CA1/_0125_ ),
    .Y(\hash/CA1/_0126_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2171_  (.A1(\hash/CA1/_1772_ ),
    .A2(\hash/CA1/_0126_ ),
    .B1(\hash/CA1/_1771_ ),
    .Y(\hash/CA1/_0127_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2172_  (.A(\hash/CA1/_1781_ ),
    .B(\hash/CA1/_0127_ ),
    .Y(\hash/CA1/_1336_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2173_  (.A(\hash/CA1/_1336_ ),
    .Y(\hash/CA1/_1147_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2174_  (.A(\hash/CA1/_1769_ ),
    .B(\hash/CA1/_1778_ ),
    .Y(\hash/CA1/_0128_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2175_  (.A1(\hash/CA1/_0120_ ),
    .A2(\hash/CA1/_0107_ ),
    .B1_N(\hash/CA1/_1768_ ),
    .Y(\hash/CA1/_0129_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2176_  (.A1(\hash/CA1/_1778_ ),
    .A2(\hash/CA1/_0129_ ),
    .B1(\hash/CA1/_1777_ ),
    .Y(\hash/CA1/_0130_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_2177_  (.A1(\hash/CA1/_0108_ ),
    .A2(\hash/CA1/_0128_ ),
    .B1(\hash/CA1/_0130_ ),
    .Y(\hash/CA1/_0131_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2178_  (.A(\hash/CA1/_1787_ ),
    .B(\hash/CA1/_0131_ ),
    .Y(\hash/CA1/_1151_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2179_  (.A(\hash/CA1/_1151_ ),
    .Y(\hash/CA1/_1339_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2180_  (.A0(\hash/g[19] ),
    .A1(\hash/f[19] ),
    .S(\hash/e[19] ),
    .X(\hash/CA1/_1788_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2181_  (.A(\hash/CA1/_1772_ ),
    .B(\hash/CA1/_1781_ ),
    .Y(\hash/CA1/_0132_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2182_  (.A(\hash/CA1/_0116_ ),
    .B(\hash/CA1/_0132_ ),
    .Y(\hash/CA1/_0133_ ));
 sky130_fd_sc_hd__nor4_1 \hash/CA1/_2183_  (.A(\hash/CA1/_0079_ ),
    .B(\hash/CA1/_0080_ ),
    .C(\hash/CA1/_0116_ ),
    .D(\hash/CA1/_0132_ ),
    .Y(\hash/CA1/_0134_ ));
 sky130_fd_sc_hd__a22oi_1 \hash/CA1/_2184_  (.A1(\hash/CA1/_0114_ ),
    .A2(\hash/CA1/_0133_ ),
    .B1(\hash/CA1/_0134_ ),
    .B2(\hash/CA1/_0058_ ),
    .Y(\hash/CA1/_0135_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2185_  (.A(\hash/CA1/_0019_ ),
    .B(\hash/CA1/_0054_ ),
    .C(\hash/CA1/_0134_ ),
    .Y(\hash/CA1/_0136_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2186_  (.A1(\hash/CA1/_1772_ ),
    .A2(\hash/CA1/_0117_ ),
    .B1(\hash/CA1/_1771_ ),
    .X(\hash/CA1/_0137_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2187_  (.A1(\hash/CA1/_1781_ ),
    .A2(\hash/CA1/_0137_ ),
    .B1(\hash/CA1/_1780_ ),
    .Y(\hash/CA1/_0138_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2188_  (.A(\hash/CA1/_0135_ ),
    .B(\hash/CA1/_0136_ ),
    .C(\hash/CA1/_0138_ ),
    .Y(\hash/CA1/_0139_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2189_  (.A(\hash/CA1/_1790_ ),
    .B(\hash/CA1/_0139_ ),
    .X(\hash/CA1/_1342_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2190_  (.A(\hash/CA1/_1342_ ),
    .Y(\hash/CA1/_1152_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2192_  (.A(\hash/CA1/_1768_ ),
    .B(\hash/CA1/_1777_ ),
    .Y(\hash/CA1/_0141_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2193_  (.A1(\hash/CA1/_0120_ ),
    .A2(\hash/CA1/_0121_ ),
    .B1(\hash/CA1/_0141_ ),
    .Y(\hash/CA1/_0142_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2194_  (.A1(\hash/CA1/_1778_ ),
    .A2(\hash/CA1/_1777_ ),
    .B1(\hash/CA1/_1787_ ),
    .X(\hash/CA1/_0143_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2195_  (.A1(\hash/CA1/_0142_ ),
    .A2(\hash/CA1/_0143_ ),
    .B1(\hash/CA1/_1786_ ),
    .Y(\hash/CA1/_0144_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2196_  (.A(\hash/CA1/_1796_ ),
    .B(\hash/CA1/_0144_ ),
    .X(\hash/CA1/_1156_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2197_  (.A(\hash/CA1/_1156_ ),
    .Y(\hash/CA1/_1345_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2198_  (.A0(\hash/g[20] ),
    .A1(\hash/f[20] ),
    .S(\hash/e[20] ),
    .X(\hash/CA1/_1797_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2199_  (.A(\hash/CA1/_1799_ ),
    .Y(\hash/CA1/_0145_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2200_  (.A(\hash/CA1/_1781_ ),
    .B(\hash/CA1/_1771_ ),
    .Y(\hash/CA1/_0146_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2201_  (.A1(\hash/CA1/_0124_ ),
    .A2(\hash/CA1/_0132_ ),
    .B1(\hash/CA1/_0146_ ),
    .Y(\hash/CA1/_0147_ ));
 sky130_fd_sc_hd__a211o_1 \hash/CA1/_2202_  (.A1(\hash/CA1/_0085_ ),
    .A2(\hash/CA1/_0133_ ),
    .B1(\hash/CA1/_0147_ ),
    .C1(\hash/CA1/_1780_ ),
    .X(\hash/CA1/_0148_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2203_  (.A1(\hash/CA1/_1790_ ),
    .A2(\hash/CA1/_0148_ ),
    .B1(\hash/CA1/_1789_ ),
    .Y(\hash/CA1/_0149_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2204_  (.A(\hash/CA1/_0145_ ),
    .B(\hash/CA1/_0149_ ),
    .Y(\hash/CA1/_1157_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2206_  (.A1(\hash/CA1/_1787_ ),
    .A2(\hash/CA1/_0131_ ),
    .B1(\hash/CA1/_1786_ ),
    .X(\hash/CA1/_0151_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2207_  (.A1(\hash/CA1/_1796_ ),
    .A2(\hash/CA1/_0151_ ),
    .B1(\hash/CA1/_1795_ ),
    .X(\hash/CA1/_0152_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2208_  (.A(\hash/CA1/_1805_ ),
    .B(\hash/CA1/_0152_ ),
    .Y(\hash/CA1/_1162_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2209_  (.A(\hash/CA1/_1162_ ),
    .Y(\hash/CA1/_1352_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2210_  (.A0(\hash/g[21] ),
    .A1(\hash/f[21] ),
    .S(\hash/e[21] ),
    .X(\hash/CA1/_1806_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2211_  (.A1(\hash/CA1/_1790_ ),
    .A2(\hash/CA1/_0139_ ),
    .B1(\hash/CA1/_1789_ ),
    .Y(\hash/CA1/_0153_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2212_  (.A1(\hash/CA1/_0145_ ),
    .A2(\hash/CA1/_0153_ ),
    .B1_N(\hash/CA1/_1798_ ),
    .Y(\hash/CA1/_0154_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2213_  (.A(\hash/CA1/_1808_ ),
    .B(\hash/CA1/_0154_ ),
    .X(\hash/CA1/_1355_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2214_  (.A(\hash/CA1/_1355_ ),
    .Y(\hash/CA1/_1161_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2216_  (.A(\hash/CA1/_1795_ ),
    .B(\hash/CA1/_1804_ ),
    .Y(\hash/CA1/_0156_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2217_  (.A1(\hash/CA1/_1796_ ),
    .A2(\hash/CA1/_1795_ ),
    .B1(\hash/CA1/_1805_ ),
    .X(\hash/CA1/_0157_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \hash/CA1/_2218_  (.A1_N(\hash/CA1/_0144_ ),
    .A2_N(\hash/CA1/_0156_ ),
    .B1(\hash/CA1/_0157_ ),
    .B2(\hash/CA1/_1804_ ),
    .Y(\hash/CA1/_0158_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2219_  (.A(\hash/CA1/_1814_ ),
    .B(\hash/CA1/_0158_ ),
    .Y(\hash/CA1/_1358_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2220_  (.A0(\hash/g[22] ),
    .A1(\hash/f[22] ),
    .S(\hash/e[22] ),
    .X(\hash/CA1/_1815_ ));
 sky130_fd_sc_hd__or3_1 \hash/CA1/_2221_  (.A(\hash/CA1/_1780_ ),
    .B(\hash/CA1/_1789_ ),
    .C(\hash/CA1/_1798_ ),
    .X(\hash/CA1/_0159_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2222_  (.A1(\hash/CA1/_0085_ ),
    .A2(\hash/CA1/_0133_ ),
    .B1(\hash/CA1/_0147_ ),
    .C1(\hash/CA1/_0159_ ),
    .Y(\hash/CA1/_0160_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_2223_  (.A(\hash/CA1/_1790_ ),
    .B(\hash/CA1/_1789_ ),
    .X(\hash/CA1/_0161_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2224_  (.A1(\hash/CA1/_1799_ ),
    .A2(\hash/CA1/_0161_ ),
    .B1(\hash/CA1/_1798_ ),
    .Y(\hash/CA1/_0162_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2225_  (.A(\hash/CA1/_0160_ ),
    .B(\hash/CA1/_0162_ ),
    .Y(\hash/CA1/_0163_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2226_  (.A1(\hash/CA1/_1808_ ),
    .A2(\hash/CA1/_0163_ ),
    .B1(\hash/CA1/_1807_ ),
    .Y(\hash/CA1/_0164_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2227_  (.A(\hash/CA1/_1817_ ),
    .B(\hash/CA1/_0164_ ),
    .Y(\hash/CA1/_1361_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2228_  (.A(\hash/CA1/_1361_ ),
    .Y(\hash/CA1/_1166_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2229_  (.A1(\hash/CA1/_1796_ ),
    .A2(\hash/CA1/_1786_ ),
    .B1(\hash/CA1/_1795_ ),
    .X(\hash/CA1/_0165_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2230_  (.A1(\hash/CA1/_1805_ ),
    .A2(\hash/CA1/_0165_ ),
    .B1(\hash/CA1/_1804_ ),
    .X(\hash/CA1/_0166_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2231_  (.A1(\hash/CA1/_1814_ ),
    .A2(\hash/CA1/_0166_ ),
    .B1(\hash/CA1/_1813_ ),
    .Y(\hash/CA1/_0167_ ));
 sky130_fd_sc_hd__and4_1 \hash/CA1/_2232_  (.A(\hash/CA1/_1787_ ),
    .B(\hash/CA1/_1796_ ),
    .C(\hash/CA1/_1805_ ),
    .D(\hash/CA1/_1814_ ),
    .X(\hash/CA1/_0168_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2233_  (.A(\hash/CA1/_0131_ ),
    .B(\hash/CA1/_0168_ ),
    .Y(\hash/CA1/_0169_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2234_  (.A(\hash/CA1/_0167_ ),
    .B(\hash/CA1/_0169_ ),
    .Y(\hash/CA1/_0170_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2235_  (.A(\hash/CA1/_1823_ ),
    .B(\hash/CA1/_0170_ ),
    .Y(\hash/CA1/_1171_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2236_  (.A(\hash/CA1/_1171_ ),
    .Y(\hash/CA1/_1364_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2237_  (.A0(\hash/g[23] ),
    .A1(\hash/f[23] ),
    .S(\hash/e[23] ),
    .X(\hash/CA1/_1824_ ));
 sky130_fd_sc_hd__a211o_1 \hash/CA1/_2238_  (.A1(\hash/CA1/_1817_ ),
    .A2(\hash/CA1/_1807_ ),
    .B1(\hash/CA1/_1816_ ),
    .C1(\hash/CA1/_1798_ ),
    .X(\hash/CA1/_0171_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2239_  (.A1(\hash/CA1/_1799_ ),
    .A2(\hash/CA1/_1789_ ),
    .B1(\hash/CA1/_0171_ ),
    .Y(\hash/CA1/_0172_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2240_  (.A(\hash/CA1/_1790_ ),
    .B(\hash/CA1/_1799_ ),
    .C(\hash/CA1/_0139_ ),
    .Y(\hash/CA1/_0173_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2241_  (.A1(\hash/CA1/_1808_ ),
    .A2(\hash/CA1/_1807_ ),
    .B1(\hash/CA1/_1817_ ),
    .Y(\hash/CA1/_0174_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2242_  (.A_N(\hash/CA1/_1816_ ),
    .B(\hash/CA1/_0174_ ),
    .Y(\hash/CA1/_0175_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA1/_2243_  (.A1(\hash/CA1/_0172_ ),
    .A2(\hash/CA1/_0173_ ),
    .B1_N(\hash/CA1/_0175_ ),
    .Y(\hash/CA1/_0176_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2244_  (.A(\hash/CA1/_1826_ ),
    .B(\hash/CA1/_0176_ ),
    .Y(\hash/CA1/_1172_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2245_  (.A(\hash/CA1/_1769_ ),
    .B(\hash/CA1/_1778_ ),
    .C(\hash/CA1/_0168_ ),
    .Y(\hash/CA1/_0177_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2246_  (.A1(\hash/CA1/_1778_ ),
    .A2(\hash/CA1/_1768_ ),
    .B1(\hash/CA1/_1777_ ),
    .X(\hash/CA1/_0178_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2247_  (.A1(\hash/CA1/_1787_ ),
    .A2(\hash/CA1/_0178_ ),
    .B1(\hash/CA1/_1786_ ),
    .Y(\hash/CA1/_0179_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2248_  (.A(\hash/CA1/_1796_ ),
    .B(\hash/CA1/_1805_ ),
    .Y(\hash/CA1/_0180_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2249_  (.A1(\hash/CA1/_1805_ ),
    .A2(\hash/CA1/_1795_ ),
    .B1(\hash/CA1/_1804_ ),
    .Y(\hash/CA1/_0181_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2250_  (.A1(\hash/CA1/_0179_ ),
    .A2(\hash/CA1/_0180_ ),
    .B1(\hash/CA1/_0181_ ),
    .Y(\hash/CA1/_0182_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2251_  (.A1(\hash/CA1/_1814_ ),
    .A2(\hash/CA1/_0182_ ),
    .B1(\hash/CA1/_1813_ ),
    .Y(\hash/CA1/_0183_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2252_  (.A1(\hash/CA1/_0121_ ),
    .A2(\hash/CA1/_0177_ ),
    .B1(\hash/CA1/_0183_ ),
    .Y(\hash/CA1/_0184_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2253_  (.A1(\hash/CA1/_1823_ ),
    .A2(\hash/CA1/_0184_ ),
    .B1(\hash/CA1/_1822_ ),
    .Y(\hash/CA1/_0185_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2254_  (.A(\hash/CA1/_1832_ ),
    .B(\hash/CA1/_0185_ ),
    .X(\hash/CA1/_1177_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2255_  (.A(\hash/CA1/_1177_ ),
    .Y(\hash/CA1/_1371_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2256_  (.A0(\hash/g[24] ),
    .A1(\hash/f[24] ),
    .S(\hash/e[24] ),
    .X(\hash/CA1/_1833_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2258_  (.A(\hash/CA1/_0145_ ),
    .B(\hash/CA1/_0149_ ),
    .Y(\hash/CA1/_0187_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2259_  (.A(\hash/CA1/_1808_ ),
    .B(\hash/CA1/_1817_ ),
    .C(\hash/CA1/_1826_ ),
    .X(\hash/CA1/_0188_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2260_  (.A1(\hash/CA1/_1808_ ),
    .A2(\hash/CA1/_1798_ ),
    .B1(\hash/CA1/_1807_ ),
    .X(\hash/CA1/_0189_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2261_  (.A1(\hash/CA1/_1817_ ),
    .A2(\hash/CA1/_0189_ ),
    .B1(\hash/CA1/_1816_ ),
    .X(\hash/CA1/_0190_ ));
 sky130_fd_sc_hd__a221o_1 \hash/CA1/_2262_  (.A1(\hash/CA1/_0187_ ),
    .A2(\hash/CA1/_0188_ ),
    .B1(\hash/CA1/_0190_ ),
    .B2(\hash/CA1/_1826_ ),
    .C1(\hash/CA1/_1825_ ),
    .X(\hash/CA1/_0191_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2263_  (.A(\hash/CA1/_1835_ ),
    .B(\hash/CA1/_0191_ ),
    .Y(\hash/CA1/_1176_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2264_  (.A1(\hash/CA1/_1787_ ),
    .A2(\hash/CA1/_0131_ ),
    .B1(\hash/CA1/_1795_ ),
    .C1(\hash/CA1/_1786_ ),
    .Y(\hash/CA1/_0192_ ));
 sky130_fd_sc_hd__o2111ai_1 \hash/CA1/_2265_  (.A1(\hash/CA1/_1796_ ),
    .A2(\hash/CA1/_1795_ ),
    .B1(\hash/CA1/_1823_ ),
    .C1(\hash/CA1/_1814_ ),
    .D1(\hash/CA1/_1805_ ),
    .Y(\hash/CA1/_0193_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2266_  (.A1(\hash/CA1/_1814_ ),
    .A2(\hash/CA1/_1804_ ),
    .B1(\hash/CA1/_1813_ ),
    .X(\hash/CA1/_0194_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2267_  (.A1(\hash/CA1/_1823_ ),
    .A2(\hash/CA1/_0194_ ),
    .B1(\hash/CA1/_1822_ ),
    .Y(\hash/CA1/_0195_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2268_  (.A1(\hash/CA1/_0192_ ),
    .A2(\hash/CA1/_0193_ ),
    .B1(\hash/CA1/_0195_ ),
    .Y(\hash/CA1/_0196_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2269_  (.A1(\hash/CA1/_1832_ ),
    .A2(\hash/CA1/_0196_ ),
    .B1(\hash/CA1/_1831_ ),
    .Y(\hash/CA1/_0197_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2270_  (.A(\hash/CA1/_1841_ ),
    .B(\hash/CA1/_0197_ ),
    .Y(\hash/CA1/_1377_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2271_  (.A0(\hash/g[25] ),
    .A1(\hash/f[25] ),
    .S(\hash/e[25] ),
    .X(\hash/CA1/_1842_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2272_  (.A(\hash/CA1/_1790_ ),
    .B(\hash/CA1/_1799_ ),
    .C(\hash/CA1/_1835_ ),
    .X(\hash/CA1/_0198_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2273_  (.A(\hash/CA1/_1826_ ),
    .B(\hash/CA1/_0175_ ),
    .C(\hash/CA1/_0198_ ),
    .Y(\hash/CA1/_0199_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2274_  (.A1(\hash/CA1/_0135_ ),
    .A2(\hash/CA1/_0136_ ),
    .B1(\hash/CA1/_0199_ ),
    .Y(\hash/CA1/_0200_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2275_  (.A1(\hash/CA1/_1772_ ),
    .A2(\hash/CA1/_0117_ ),
    .B1(\hash/CA1/_1780_ ),
    .C1(\hash/CA1/_1771_ ),
    .Y(\hash/CA1/_0201_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_2276_  (.A1(\hash/CA1/_1781_ ),
    .A2(\hash/CA1/_1780_ ),
    .B1(\hash/CA1/_1790_ ),
    .C1(\hash/CA1/_1799_ ),
    .Y(\hash/CA1/_0202_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2277_  (.A1(\hash/CA1/_0201_ ),
    .A2(\hash/CA1/_0202_ ),
    .B1(\hash/CA1/_0172_ ),
    .Y(\hash/CA1/_0203_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2278_  (.A(\hash/CA1/_1826_ ),
    .B(\hash/CA1/_1835_ ),
    .C(\hash/CA1/_0175_ ),
    .X(\hash/CA1/_0204_ ));
 sky130_fd_sc_hd__a22o_1 \hash/CA1/_2279_  (.A1(\hash/CA1/_1835_ ),
    .A2(\hash/CA1/_1825_ ),
    .B1(\hash/CA1/_0203_ ),
    .B2(\hash/CA1/_0204_ ),
    .X(\hash/CA1/_0205_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2280_  (.A(\hash/CA1/_1834_ ),
    .B(\hash/CA1/_0200_ ),
    .C(\hash/CA1/_0205_ ),
    .Y(\hash/CA1/_0206_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2281_  (.A(\hash/CA1/_1844_ ),
    .B(\hash/CA1/_0206_ ),
    .X(\hash/CA1/_1181_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2283_  (.A(\hash/CA1/_1823_ ),
    .B(\hash/CA1/_1832_ ),
    .Y(\hash/CA1/_0208_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2284_  (.A(\hash/CA1/_0177_ ),
    .B(\hash/CA1/_0208_ ),
    .Y(\hash/CA1/_0209_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2285_  (.A1(\hash/CA1/_1760_ ),
    .A2(\hash/CA1/_0098_ ),
    .A3(\hash/CA1/_0100_ ),
    .B1(\hash/CA1/_0209_ ),
    .Y(\hash/CA1/_0210_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2286_  (.A(\hash/CA1/_0183_ ),
    .B(\hash/CA1/_0208_ ),
    .Y(\hash/CA1/_0211_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2287_  (.A1(\hash/CA1/_1832_ ),
    .A2(\hash/CA1/_1822_ ),
    .B1(\hash/CA1/_0211_ ),
    .Y(\hash/CA1/_0212_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2288_  (.A(\hash/CA1/_0210_ ),
    .B(\hash/CA1/_0212_ ),
    .Y(\hash/CA1/_0213_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2289_  (.A1(\hash/CA1/_1831_ ),
    .A2(\hash/CA1/_0213_ ),
    .B1(\hash/CA1/_1841_ ),
    .Y(\hash/CA1/_0214_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2290_  (.A(\hash/CA1/_1840_ ),
    .B_N(\hash/CA1/_0214_ ),
    .Y(\hash/CA1/_0215_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2291_  (.A(\hash/CA1/_1850_ ),
    .B(\hash/CA1/_0215_ ),
    .Y(\hash/CA1/_1384_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2292_  (.A0(\hash/g[26] ),
    .A1(\hash/f[26] ),
    .S(\hash/e[26] ),
    .X(\hash/CA1/_1851_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2294_  (.A(\hash/CA1/_1835_ ),
    .B(\hash/CA1/_1844_ ),
    .C(\hash/CA1/_0188_ ),
    .Y(\hash/CA1/_0217_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2295_  (.A(\hash/CA1/_0160_ ),
    .B(\hash/CA1/_0162_ ),
    .C(\hash/CA1/_0217_ ),
    .Y(\hash/CA1/_0218_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2296_  (.A1(\hash/CA1/_1826_ ),
    .A2(\hash/CA1/_1816_ ),
    .B1(\hash/CA1/_1825_ ),
    .X(\hash/CA1/_0219_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2297_  (.A1(\hash/CA1/_1835_ ),
    .A2(\hash/CA1/_0219_ ),
    .B1(\hash/CA1/_1834_ ),
    .Y(\hash/CA1/_0220_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2298_  (.A(\hash/CA1/_1817_ ),
    .B(\hash/CA1/_1826_ ),
    .C(\hash/CA1/_1835_ ),
    .D(\hash/CA1/_1807_ ),
    .Y(\hash/CA1/_0221_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA1/_2299_  (.A1(\hash/CA1/_0220_ ),
    .A2(\hash/CA1/_0221_ ),
    .B1_N(\hash/CA1/_1844_ ),
    .Y(\hash/CA1/_0222_ ));
 sky130_fd_sc_hd__or3_1 \hash/CA1/_2300_  (.A(\hash/CA1/_1843_ ),
    .B(\hash/CA1/_0218_ ),
    .C(\hash/CA1/_0222_ ),
    .X(\hash/CA1/_0223_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2301_  (.A(\hash/CA1/_1853_ ),
    .B(\hash/CA1/_0223_ ),
    .X(\hash/CA1/_1387_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2302_  (.A(\hash/CA1/_1387_ ),
    .Y(\hash/CA1/_1186_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2303_  (.A(\hash/CA1/_1823_ ),
    .B(\hash/CA1/_1832_ ),
    .C(\hash/CA1/_1841_ ),
    .D(\hash/CA1/_1850_ ),
    .Y(\hash/CA1/_0224_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2304_  (.A(\hash/CA1/_0224_ ),
    .Y(\hash/CA1/_0225_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2305_  (.A(\hash/CA1/_0168_ ),
    .B(\hash/CA1/_0225_ ),
    .Y(\hash/CA1/_0226_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2306_  (.A1(\hash/CA1/_1832_ ),
    .A2(\hash/CA1/_1822_ ),
    .B1(\hash/CA1/_1831_ ),
    .X(\hash/CA1/_0227_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2307_  (.A1(\hash/CA1/_1841_ ),
    .A2(\hash/CA1/_0227_ ),
    .B1(\hash/CA1/_1840_ ),
    .X(\hash/CA1/_0228_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2308_  (.A1(\hash/CA1/_1850_ ),
    .A2(\hash/CA1/_0228_ ),
    .B1(\hash/CA1/_1849_ ),
    .Y(\hash/CA1/_0229_ ));
 sky130_fd_sc_hd__o221ai_1 \hash/CA1/_2309_  (.A1(\hash/CA1/_0167_ ),
    .A2(\hash/CA1/_0224_ ),
    .B1(\hash/CA1/_0226_ ),
    .B2(\hash/CA1/_0130_ ),
    .C1(\hash/CA1/_0229_ ),
    .Y(\hash/CA1/_0230_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2310_  (.A(\hash/CA1/_1753_ ),
    .B(\hash/CA1/_1761_ ),
    .C(\hash/CA1/_1769_ ),
    .D(\hash/CA1/_1778_ ),
    .Y(\hash/CA1/_0231_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2311_  (.A(\hash/CA1/_0090_ ),
    .B(\hash/CA1/_0226_ ),
    .C(\hash/CA1/_0231_ ),
    .Y(\hash/CA1/_0232_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2312_  (.A(\hash/CA1/_0093_ ),
    .B(\hash/CA1/_0226_ ),
    .C(\hash/CA1/_0231_ ),
    .Y(\hash/CA1/_0233_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2313_  (.A1(\hash/CA1/_0050_ ),
    .A2(\hash/CA1/_0232_ ),
    .B1(\hash/CA1/_0233_ ),
    .Y(\hash/CA1/_0234_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2314_  (.A(\hash/CA1/_0230_ ),
    .B_N(\hash/CA1/_0234_ ),
    .Y(\hash/CA1/_0235_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2315_  (.A(\hash/CA1/_1859_ ),
    .B(\hash/CA1/_0235_ ),
    .Y(\hash/CA1/_1191_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2316_  (.A(\hash/CA1/_1191_ ),
    .Y(\hash/CA1/_1195_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2317_  (.A0(\hash/g[27] ),
    .A1(\hash/f[27] ),
    .S(\hash/e[27] ),
    .X(\hash/CA1/_1860_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2318_  (.A1(\hash/CA1/_1850_ ),
    .A2(\hash/CA1/_1840_ ),
    .B1(\hash/CA1/_1849_ ),
    .Y(\hash/CA1/_0236_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2319_  (.A(\hash/CA1/_1831_ ),
    .B(\hash/CA1/_1858_ ),
    .Y(\hash/CA1/_0237_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2320_  (.A(\hash/CA1/_0210_ ),
    .B(\hash/CA1/_0212_ ),
    .C(\hash/CA1/_0236_ ),
    .D(\hash/CA1/_0237_ ),
    .Y(\hash/CA1/_0238_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2321_  (.A1(\hash/CA1/_1841_ ),
    .A2(\hash/CA1/_1850_ ),
    .B1(\hash/CA1/_1858_ ),
    .Y(\hash/CA1/_0239_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2322_  (.A(\hash/CA1/_0236_ ),
    .B(\hash/CA1/_0239_ ),
    .Y(\hash/CA1/_0240_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_2323_  (.A(\hash/CA1/_1859_ ),
    .B(\hash/CA1/_1858_ ),
    .X(\hash/CA1/_0241_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2324_  (.A(\hash/CA1/_0238_ ),
    .B(\hash/CA1/_0240_ ),
    .C(\hash/CA1/_0241_ ),
    .Y(\hash/CA1/_0242_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2325_  (.A(\hash/CA1/_1867_ ),
    .B(\hash/CA1/_0242_ ),
    .Y(\hash/CA1/_1197_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2326_  (.A(\hash/CA1/_1197_ ),
    .Y(\hash/CA1/_1200_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2327_  (.A0(\hash/g[28] ),
    .A1(\hash/f[28] ),
    .S(\hash/e[28] ),
    .X(\hash/CA1/_1868_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2328_  (.A(\hash/CA1/_1858_ ),
    .B(\hash/CA1/_1866_ ),
    .C(\hash/CA1/_0230_ ),
    .Y(\hash/CA1/_0243_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2329_  (.A1(\hash/CA1/_1867_ ),
    .A2(\hash/CA1/_0241_ ),
    .B1(\hash/CA1/_1866_ ),
    .Y(\hash/CA1/_0244_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2330_  (.A1(\hash/CA1/_0234_ ),
    .A2(\hash/CA1/_0243_ ),
    .B1(\hash/CA1/_0244_ ),
    .Y(\hash/CA1/_0245_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2331_  (.A(\hash/CA1/_1874_ ),
    .B(\hash/CA1/_0245_ ),
    .X(\hash/CA1/_1202_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2332_  (.A(\hash/CA1/_1202_ ),
    .Y(\hash/CA1/_1207_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2333_  (.A0(\hash/g[29] ),
    .A1(\hash/f[29] ),
    .S(\hash/e[29] ),
    .X(\hash/CA1/_1875_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2334_  (.A(\hash/CA1/_1862_ ),
    .B(\hash/CA1/_1861_ ),
    .Y(\hash/CA1/_0246_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2335_  (.A(\hash/CA1/_0246_ ),
    .B_N(\hash/CA1/_1870_ ),
    .Y(\hash/CA1/_0247_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2336_  (.A1(\hash/CA1/_1853_ ),
    .A2(\hash/CA1/_1843_ ),
    .B1(\hash/CA1/_1852_ ),
    .X(\hash/CA1/_0248_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2337_  (.A1(\hash/CA1/_1862_ ),
    .A2(\hash/CA1/_0248_ ),
    .B1(\hash/CA1/_1861_ ),
    .Y(\hash/CA1/_0249_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2338_  (.A(\hash/CA1/_0249_ ),
    .B_N(\hash/CA1/_1870_ ),
    .Y(\hash/CA1/_0250_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2339_  (.A1(\hash/CA1/_1869_ ),
    .A2(\hash/CA1/_0250_ ),
    .B1(\hash/CA1/_1877_ ),
    .Y(\hash/CA1/_0251_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2340_  (.A(\hash/CA1/_1862_ ),
    .B(\hash/CA1/_1870_ ),
    .C(\hash/CA1/_1877_ ),
    .X(\hash/CA1/_0252_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2341_  (.A1(\hash/CA1/_1870_ ),
    .A2(\hash/CA1/_1861_ ),
    .B1(\hash/CA1/_1869_ ),
    .X(\hash/CA1/_0253_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2342_  (.A(\hash/CA1/_1877_ ),
    .B(\hash/CA1/_0248_ ),
    .C(\hash/CA1/_0253_ ),
    .Y(\hash/CA1/_0254_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA1/_2343_  (.A_N(\hash/CA1/_0206_ ),
    .B(\hash/CA1/_1853_ ),
    .C(\hash/CA1/_1844_ ),
    .Y(\hash/CA1/_0255_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA1/_2344_  (.A0(\hash/CA1/_0252_ ),
    .A1(\hash/CA1/_0254_ ),
    .S(\hash/CA1/_0255_ ),
    .Y(\hash/CA1/_0256_ ));
 sky130_fd_sc_hd__o311a_1 \hash/CA1/_2345_  (.A1(\hash/CA1/_1877_ ),
    .A2(\hash/CA1/_1869_ ),
    .A3(\hash/CA1/_0247_ ),
    .B1(\hash/CA1/_0251_ ),
    .C1(\hash/CA1/_0256_ ),
    .X(\hash/CA1/_1203_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2346_  (.A(\hash/CA1/_1203_ ),
    .Y(\hash/CA1/_1208_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA1/_2347_  (.A0(\hash/g[30] ),
    .A1(\hash/f[30] ),
    .S(\hash/e[30] ),
    .X(\hash/CA1/_1882_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2348_  (.A(\hash/CA1/_1519_ ),
    .Y(\hash/CA1/_0993_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2349_  (.A(\k_value1[1] ),
    .Y(\hash/CA1/_1054_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2350_  (.A(\hash/CA1/s1[1] ),
    .Y(\hash/CA1/_1059_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2351_  (.A(\hash/h[4] ),
    .Y(\hash/CA1/_1076_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2352_  (.A(\hash/h[9] ),
    .Y(\hash/CA1/_1099_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2353_  (.A(\hash/h[10] ),
    .Y(\hash/CA1/_1104_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2354_  (.A(\hash/h[11] ),
    .Y(\hash/CA1/_1109_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2355_  (.A(\hash/h[12] ),
    .Y(\hash/CA1/_1114_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2356_  (.A(\hash/h[13] ),
    .Y(\hash/CA1/_1119_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2357_  (.A(\hash/h[14] ),
    .Y(\hash/CA1/_1124_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2358_  (.A(\hash/h[16] ),
    .Y(\hash/CA1/_1135_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2359_  (.A(\hash/h[17] ),
    .Y(\hash/CA1/_1140_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2360_  (.A(\hash/h[18] ),
    .Y(\hash/CA1/_1145_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2361_  (.A(\hash/h[19] ),
    .Y(\hash/CA1/_1150_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2362_  (.A(\hash/h[20] ),
    .Y(\hash/CA1/_1155_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2363_  (.A(\hash/h[21] ),
    .Y(\hash/CA1/_1160_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2364_  (.A(\hash/h[22] ),
    .Y(\hash/CA1/_1165_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2365_  (.A(\hash/h[23] ),
    .Y(\hash/CA1/_1170_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2366_  (.A(\hash/h[24] ),
    .Y(\hash/CA1/_1175_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2367_  (.A(\hash/h[25] ),
    .Y(\hash/CA1/_1180_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2368_  (.A(\hash/h[26] ),
    .Y(\hash/CA1/_1185_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2369_  (.A(\hash/d[0] ),
    .Y(\hash/CA1/_1213_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2370_  (.A(\hash/d[1] ),
    .Y(\hash/CA1/_1218_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2371_  (.A(\hash/d[2] ),
    .Y(\hash/CA1/_1224_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2372_  (.A(\hash/d[3] ),
    .Y(\hash/CA1/_1233_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2373_  (.A(\hash/d[8] ),
    .Y(\hash/CA1/_1270_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2374_  (.A(\hash/d[15] ),
    .Y(\hash/CA1/_1315_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2375_  (.A(\hash/d[27] ),
    .Y(\hash/CA1/_1390_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2376_  (.A(\hash/d[28] ),
    .Y(\hash/CA1/_1396_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2377_  (.A(\hash/d[29] ),
    .Y(\hash/CA1/_1403_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2378_  (.A(\hash/h[0] ),
    .Y(\hash/CA1/_1214_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2379_  (.A(\w_value1[1] ),
    .Y(\hash/CA1/_1055_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2380_  (.A(\hash/h[1] ),
    .Y(\hash/CA1/_1219_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2381_  (.A(\hash/h[2] ),
    .Y(\hash/CA1/_1225_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2382_  (.A(\hash/h[3] ),
    .Y(\hash/CA1/_1234_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2383_  (.A(\hash/h[8] ),
    .Y(\hash/CA1/_1098_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2384_  (.A(\hash/h[15] ),
    .Y(\hash/CA1/_1134_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2385_  (.A(\hash/h[27] ),
    .Y(\hash/CA1/_1194_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2386_  (.A(\hash/h[28] ),
    .Y(\hash/CA1/_1201_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2387_  (.A(\hash/h[29] ),
    .Y(\hash/CA1/_1206_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2388_  (.A(\hash/CA1/_1976_ ),
    .Y(\hash/CA1/_1424_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2389_  (.A(\hash/CA1/_1638_ ),
    .Y(\hash/CA1/_1056_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2390_  (.A(\hash/CA1/_1641_ ),
    .Y(\hash/CA1/_1061_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2391_  (.A(\hash/CA1/_1814_ ),
    .B(\hash/CA1/_0158_ ),
    .X(\hash/CA1/_1167_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2392_  (.A(\hash/CA1/_1841_ ),
    .B(\hash/CA1/_0197_ ),
    .X(\hash/CA1/_1182_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2393_  (.A(\hash/CA1/_1850_ ),
    .B(\hash/CA1/_0215_ ),
    .X(\hash/CA1/_1187_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2394_  (.A(\hash/CA1/_1250_ ),
    .Y(\hash/CA1/_1253_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2395_  (.A(\hash/CA1/_1257_ ),
    .Y(\hash/CA1/_1260_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2396_  (.A(\hash/CA1/_1264_ ),
    .Y(\hash/CA1/_1267_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2397_  (.A(\hash/CA1/_1974_ ),
    .Y(\hash/CA1/_1417_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2398_  (.A(\hash/CA1/_1419_ ),
    .Y(\hash/p2[2] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2399_  (.A(\hash/CA1/_1422_ ),
    .Y(\hash/p3[0] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2400_  (.A(\hash/CA1/_1427_ ),
    .Y(\hash/p3[2] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2401_  (.A(\hash/CA1/_0992_ ),
    .Y(\hash/CA1/_0995_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2402_  (.A(\hash/CA1/_1071_ ),
    .Y(\hash/CA1/_1423_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2403_  (.A(\hash/CA1/_1232_ ),
    .Y(\hash/CA1/_1416_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2404_  (.A(\hash/CA1/_1278_ ),
    .Y(\hash/CA1/_1279_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2405_  (.A(\hash/CA1/_1284_ ),
    .Y(\hash/CA1/_1286_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2406_  (.A(\hash/CA1/_1291_ ),
    .Y(\hash/CA1/_1292_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2407_  (.A(\hash/CA1/_1298_ ),
    .Y(\hash/CA1/_1299_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2408_  (.A(\hash/CA1/_1323_ ),
    .Y(\hash/CA1/_1324_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2409_  (.A(\hash/CA1/_1347_ ),
    .Y(\hash/CA1/_1348_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2410_  (.A(\hash/CA1/_1366_ ),
    .Y(\hash/CA1/_1368_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2411_  (.A(\hash/CA1/_1379_ ),
    .Y(\hash/CA1/_1380_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2412_  (.A(\hash/CA1/_0989_ ),
    .Y(\hash/CA1/_0994_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2413_  (.A(\hash/CA1/_1066_ ),
    .Y(\hash/CA1/_1425_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2414_  (.A(\hash/CA1/_1243_ ),
    .Y(\hash/CA1/_1252_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2415_  (.A(\hash/CA1/_1249_ ),
    .Y(\hash/CA1/_1259_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2416_  (.A(\hash/CA1/_1256_ ),
    .Y(\hash/CA1/_1266_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2417_  (.A(\hash/CA1/_1277_ ),
    .Y(\hash/CA1/_1285_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2418_  (.A(\hash/CA1/_1283_ ),
    .Y(\hash/CA1/_1293_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2419_  (.A(\hash/CA1/_1290_ ),
    .Y(\hash/CA1/_1300_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2420_  (.A(\hash/CA1/_1340_ ),
    .Y(\hash/CA1/_1349_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2421_  (.A(\hash/CA1/_1359_ ),
    .Y(\hash/CA1/_1367_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2422_  (.A(\hash/CA1/_1372_ ),
    .Y(\hash/CA1/_1381_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2423_  (.A(\hash/CA1/_1080_ ),
    .Y(\hash/CA1/_1667_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2424_  (.A(\hash/CA1/_1102_ ),
    .Y(\hash/CA1/_1712_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2425_  (.A(\hash/CA1/_1107_ ),
    .Y(\hash/CA1/_1721_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2426_  (.A(\hash/CA1/_1118_ ),
    .Y(\hash/CA1/_1730_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2427_  (.A(\hash/CA1/_1123_ ),
    .Y(\hash/CA1/_1739_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2428_  (.A(\hash/CA1/_1122_ ),
    .Y(\hash/CA1/_1748_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2429_  (.A(\hash/CA1/_1127_ ),
    .Y(\hash/CA1/_1757_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2430_  (.A(\hash/CA1/_1138_ ),
    .Y(\hash/CA1/_1773_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2431_  (.A(\hash/CA1/_1149_ ),
    .Y(\hash/CA1/_1782_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2432_  (.A(\hash/CA1/_1154_ ),
    .Y(\hash/CA1/_1791_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2433_  (.A(\hash/CA1/_1153_ ),
    .Y(\hash/CA1/_1800_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2434_  (.A(\hash/CA1/_1158_ ),
    .Y(\hash/CA1/_1809_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2435_  (.A(\hash/CA1/_1163_ ),
    .Y(\hash/CA1/_1818_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2436_  (.A(\hash/CA1/_1174_ ),
    .Y(\hash/CA1/_1827_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2437_  (.A(\hash/CA1/_1179_ ),
    .Y(\hash/CA1/_1836_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2438_  (.A(\hash/CA1/_1178_ ),
    .Y(\hash/CA1/_1845_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2439_  (.A(\hash/CA1/_1183_ ),
    .Y(\hash/CA1/_1854_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2440_  (.A1(\hash/CA1/_1853_ ),
    .A2(\hash/CA1/_1843_ ),
    .B1(\hash/CA1/_1852_ ),
    .Y(\hash/CA1/_0257_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2441_  (.A(\hash/CA1/_0257_ ),
    .B(\hash/CA1/_0255_ ),
    .Y(\hash/CA1/_0258_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2442_  (.A(\hash/CA1/_1862_ ),
    .B(\hash/CA1/_0258_ ),
    .X(\hash/CA1/_1190_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2443_  (.A(\hash/CA1/_1188_ ),
    .Y(\hash/CA1/_1863_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2444_  (.A(\hash/CA1/_0218_ ),
    .B(\hash/CA1/_0222_ ),
    .Y(\hash/CA1/_0259_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2445_  (.A(\hash/CA1/_1843_ ),
    .B(\hash/CA1/_1852_ ),
    .C(\hash/CA1/_1861_ ),
    .Y(\hash/CA1/_0260_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2446_  (.A(\hash/CA1/_1853_ ),
    .B(\hash/CA1/_1852_ ),
    .C(\hash/CA1/_1861_ ),
    .Y(\hash/CA1/_0261_ ));
 sky130_fd_sc_hd__a211o_1 \hash/CA1/_2447_  (.A1(\hash/CA1/_0259_ ),
    .A2(\hash/CA1/_0260_ ),
    .B1(\hash/CA1/_0261_ ),
    .C1(\hash/CA1/_0246_ ),
    .X(\hash/CA1/_0262_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2448_  (.A(\hash/CA1/_1870_ ),
    .B(\hash/CA1/_0262_ ),
    .Y(\hash/CA1/_1196_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2449_  (.A(\hash/CA1/_1058_ ),
    .Y(\hash/CA1/_1065_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2450_  (.A(\hash/CA1/_1063_ ),
    .Y(\hash/CA1/_1064_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2451_  (.A(\hash/CA1/_1220_ ),
    .Y(\hash/CA1/_1229_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2452_  (.A(\hash/CA1/_1062_ ),
    .B(\hash/CA1/_1652_ ),
    .Y(\hash/CA1/_1069_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2453_  (.A(\hash/CA1/_1227_ ),
    .Y(\hash/CA1/_1238_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2454_  (.A1(\hash/CA1/_1641_ ),
    .A2(\hash/CA1/_1647_ ),
    .B1(\hash/CA1/_1646_ ),
    .X(\hash/CA1/_0263_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2455_  (.A1(\hash/CA1/_1652_ ),
    .A2(\hash/CA1/_0263_ ),
    .B1(\hash/CA1/_1651_ ),
    .Y(\hash/CA1/_0264_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2456_  (.A(\hash/CA1/_1659_ ),
    .B(\hash/CA1/_0264_ ),
    .Y(\hash/CA1/_1072_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2457_  (.A(\hash/CA1/_1236_ ),
    .Y(\hash/CA1/_1246_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2458_  (.A1(\hash/CA1/_1663_ ),
    .A2(\hash/CA1/_1655_ ),
    .B1(\hash/CA1/_1662_ ),
    .Y(\hash/CA1/_0265_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2459_  (.A1(\hash/CA1/_0001_ ),
    .A2(\hash/CA1/_0021_ ),
    .B1(\hash/CA1/_0265_ ),
    .Y(\hash/CA1/_0266_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2460_  (.A(\hash/CA1/_1671_ ),
    .B(\hash/CA1/_0266_ ),
    .X(\hash/CA1/_1082_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2461_  (.A(\hash/CA1/_0022_ ),
    .B(\hash/CA1/_0265_ ),
    .Y(\hash/CA1/_0267_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2462_  (.A1(\hash/CA1/_1671_ ),
    .A2(\hash/CA1/_0267_ ),
    .B1(\hash/CA1/_1670_ ),
    .Y(\hash/CA1/_0268_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2463_  (.A(\hash/CA1/_1679_ ),
    .B(\hash/CA1/_0268_ ),
    .Y(\hash/CA1/_1086_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2464_  (.A(\hash/CA1/_1254_ ),
    .Y(\hash/CA1/_1897_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2465_  (.A(\hash/CA1/_0028_ ),
    .B(\hash/CA1/_0031_ ),
    .Y(\hash/CA1/_0269_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2466_  (.A(\hash/CA1/_1686_ ),
    .B(\hash/CA1/_0269_ ),
    .Y(\hash/CA1/_1090_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2467_  (.A(\hash/CA1/_1261_ ),
    .Y(\hash/CA1/_1901_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2468_  (.A(\hash/CA1/_1682_ ),
    .Y(\hash/CA1/_0270_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2469_  (.A1(\hash/CA1/_0270_ ),
    .A2(\hash/CA1/_0014_ ),
    .B1(\hash/CA1/_0015_ ),
    .Y(\hash/CA1/_0271_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2470_  (.A1(\hash/CA1/_1689_ ),
    .A2(\hash/CA1/_0271_ ),
    .B1(\hash/CA1/_1688_ ),
    .Y(\hash/CA1/_0272_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2471_  (.A(\hash/CA1/_1696_ ),
    .B(\hash/CA1/_0272_ ),
    .Y(\hash/CA1/_1094_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2472_  (.A(\hash/CA1/_1280_ ),
    .Y(\hash/CA1/_1911_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2473_  (.A(\hash/CA1/_1287_ ),
    .Y(\hash/CA1/_1915_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2474_  (.A(\hash/CA1/_1294_ ),
    .Y(\hash/CA1/_1919_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2475_  (.A(\hash/CA1/_1301_ ),
    .Y(\hash/CA1/_1923_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2476_  (.A(\hash/CA1/_1326_ ),
    .Y(\hash/CA1/_1930_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2477_  (.A(\hash/CA1/_1350_ ),
    .Y(\hash/CA1/_1943_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2478_  (.A(\hash/CA1/_1370_ ),
    .Y(\hash/CA1/_1948_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2479_  (.A(\hash/CA1/_1392_ ),
    .Y(\hash/CA1/_1393_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2480_  (.A(\hash/CA1/_1391_ ),
    .Y(\hash/CA1/_1399_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2481_  (.A(\hash/CA1/_1407_ ),
    .Y(\hash/CA1/_1964_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2482_  (.A(\hash/CA1/_1223_ ),
    .Y(\hash/CA1/_1973_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2483_  (.A(\hash/CA1/_1421_ ),
    .Y(\hash/CA1/_1975_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2484_  (.A(\hash/b[1] ),
    .B(\hash/a[1] ),
    .C(\hash/c[1] ),
    .X(\hash/CA1/_1413_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2485_  (.A(\hash/b[2] ),
    .B(\hash/a[2] ),
    .C(\hash/c[2] ),
    .X(\hash/CA1/_1432_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2486_  (.A(\hash/b[3] ),
    .B(\hash/a[3] ),
    .C(\hash/c[3] ),
    .X(\hash/CA1/_1435_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2487_  (.A(\hash/b[4] ),
    .B(\hash/a[4] ),
    .C(\hash/c[4] ),
    .X(\hash/CA1/_1438_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2488_  (.A(\hash/b[5] ),
    .B(\hash/a[5] ),
    .C(\hash/c[5] ),
    .X(\hash/CA1/_1441_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2489_  (.A(\hash/b[6] ),
    .B(\hash/a[6] ),
    .C(\hash/c[6] ),
    .X(\hash/CA1/_1444_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2490_  (.A(\hash/b[7] ),
    .B(\hash/a[7] ),
    .C(\hash/c[7] ),
    .X(\hash/CA1/_1447_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2491_  (.A(\hash/b[8] ),
    .B(\hash/a[8] ),
    .C(\hash/c[8] ),
    .X(\hash/CA1/_1450_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2492_  (.A(\hash/b[9] ),
    .B(\hash/a[9] ),
    .C(\hash/c[9] ),
    .X(\hash/CA1/_1453_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2493_  (.A(\hash/b[10] ),
    .B(\hash/a[10] ),
    .C(\hash/c[10] ),
    .X(\hash/CA1/_1456_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2494_  (.A(\hash/b[11] ),
    .B(\hash/a[11] ),
    .C(\hash/c[11] ),
    .X(\hash/CA1/_1459_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2495_  (.A(\hash/b[12] ),
    .B(\hash/a[12] ),
    .C(\hash/c[12] ),
    .X(\hash/CA1/_1462_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2496_  (.A(\hash/b[13] ),
    .B(\hash/a[13] ),
    .C(\hash/c[13] ),
    .X(\hash/CA1/_1465_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2497_  (.A(\hash/b[14] ),
    .B(\hash/a[14] ),
    .C(\hash/c[14] ),
    .X(\hash/CA1/_1468_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2498_  (.A(\hash/b[15] ),
    .B(\hash/a[15] ),
    .C(\hash/c[15] ),
    .X(\hash/CA1/_1471_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2499_  (.A(\hash/b[16] ),
    .B(\hash/a[16] ),
    .C(\hash/c[16] ),
    .X(\hash/CA1/_1474_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2500_  (.A(\hash/b[17] ),
    .B(\hash/a[17] ),
    .C(\hash/c[17] ),
    .X(\hash/CA1/_1477_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2501_  (.A(\hash/b[18] ),
    .B(\hash/a[18] ),
    .C(\hash/c[18] ),
    .X(\hash/CA1/_1480_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2502_  (.A(\hash/b[19] ),
    .B(\hash/a[19] ),
    .C(\hash/c[19] ),
    .X(\hash/CA1/_1483_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2503_  (.A(\hash/b[20] ),
    .B(\hash/a[20] ),
    .C(\hash/c[20] ),
    .X(\hash/CA1/_1486_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2504_  (.A(\hash/b[21] ),
    .B(\hash/a[21] ),
    .C(\hash/c[21] ),
    .X(\hash/CA1/_1489_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2505_  (.A(\hash/b[22] ),
    .B(\hash/a[22] ),
    .C(\hash/c[22] ),
    .X(\hash/CA1/_1492_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2506_  (.A(\hash/b[23] ),
    .B(\hash/a[23] ),
    .C(\hash/c[23] ),
    .X(\hash/CA1/_1495_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2507_  (.A(\hash/b[24] ),
    .B(\hash/a[24] ),
    .C(\hash/c[24] ),
    .X(\hash/CA1/_1498_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2508_  (.A(\hash/b[25] ),
    .B(\hash/a[25] ),
    .C(\hash/c[25] ),
    .X(\hash/CA1/_1501_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2509_  (.A(\hash/b[26] ),
    .B(\hash/a[26] ),
    .C(\hash/c[26] ),
    .X(\hash/CA1/_1504_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2510_  (.A(\hash/b[27] ),
    .B(\hash/a[27] ),
    .C(\hash/c[27] ),
    .X(\hash/CA1/_1507_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2511_  (.A(\hash/b[28] ),
    .B(\hash/a[28] ),
    .C(\hash/c[28] ),
    .X(\hash/CA1/_1510_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2512_  (.A(\hash/b[29] ),
    .B(\hash/a[29] ),
    .C(\hash/c[29] ),
    .X(\hash/CA1/_1513_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2513_  (.A(\hash/b[30] ),
    .B(\hash/a[30] ),
    .C(\hash/c[30] ),
    .X(\hash/CA1/_1516_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2514_  (.A(\hash/CA1/_0997_ ),
    .Y(\hash/p4[2] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2515_  (.A(\hash/CA1/_0996_ ),
    .B(\hash/CA1/_1523_ ),
    .Y(\hash/p4[3] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2516_  (.A1(\hash/CA1/_1519_ ),
    .A2(\hash/CA1/_1521_ ),
    .B1(\hash/CA1/_1520_ ),
    .X(\hash/CA1/_0273_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2517_  (.A1(\hash/CA1/_1523_ ),
    .A2(\hash/CA1/_0273_ ),
    .B1(\hash/CA1/_1522_ ),
    .Y(\hash/CA1/_0274_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2518_  (.A(\hash/CA1/_1525_ ),
    .B(\hash/CA1/_0274_ ),
    .Y(\hash/p4[4] ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2519_  (.A_N(\hash/CA1/_0996_ ),
    .B(\hash/CA1/_1523_ ),
    .Y(\hash/CA1/_0275_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2520_  (.A_N(\hash/CA1/_1522_ ),
    .B(\hash/CA1/_0275_ ),
    .Y(\hash/CA1/_0276_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2521_  (.A1(\hash/CA1/_1525_ ),
    .A2(\hash/CA1/_0276_ ),
    .B1(\hash/CA1/_1524_ ),
    .Y(\hash/CA1/_0277_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2522_  (.A(\hash/CA1/_1527_ ),
    .B(\hash/CA1/_0277_ ),
    .Y(\hash/p4[5] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2523_  (.A(\hash/CA1/_1525_ ),
    .Y(\hash/CA1/_0278_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2524_  (.A1(\hash/CA1/_0278_ ),
    .A2(\hash/CA1/_0274_ ),
    .B1_N(\hash/CA1/_1524_ ),
    .Y(\hash/CA1/_0279_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2525_  (.A1(\hash/CA1/_1527_ ),
    .A2(\hash/CA1/_0279_ ),
    .B1(\hash/CA1/_1526_ ),
    .Y(\hash/CA1/_0280_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2526_  (.A(\hash/CA1/_1529_ ),
    .B(\hash/CA1/_0280_ ),
    .Y(\hash/p4[6] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2527_  (.A(\hash/CA1/_1522_ ),
    .B(\hash/CA1/_1524_ ),
    .Y(\hash/CA1/_0281_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_2528_  (.A1(\hash/CA1/_1525_ ),
    .A2(\hash/CA1/_1524_ ),
    .B1(\hash/CA1/_1529_ ),
    .C1(\hash/CA1/_1527_ ),
    .Y(\hash/CA1/_0282_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2529_  (.A1(\hash/CA1/_0275_ ),
    .A2(\hash/CA1/_0281_ ),
    .B1(\hash/CA1/_0282_ ),
    .Y(\hash/CA1/_0283_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2530_  (.A1(\hash/CA1/_1529_ ),
    .A2(\hash/CA1/_1526_ ),
    .B1(\hash/CA1/_1528_ ),
    .X(\hash/CA1/_0284_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2531_  (.A(\hash/CA1/_0283_ ),
    .B(\hash/CA1/_0284_ ),
    .Y(\hash/CA1/_0285_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2532_  (.A(\hash/CA1/_1531_ ),
    .B(\hash/CA1/_0285_ ),
    .Y(\hash/p4[7] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2533_  (.A(\hash/CA1/_1529_ ),
    .Y(\hash/CA1/_0286_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2534_  (.A1(\hash/CA1/_0286_ ),
    .A2(\hash/CA1/_0280_ ),
    .B1_N(\hash/CA1/_1528_ ),
    .Y(\hash/CA1/_0287_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2535_  (.A1(\hash/CA1/_1531_ ),
    .A2(\hash/CA1/_0287_ ),
    .B1(\hash/CA1/_1530_ ),
    .Y(\hash/CA1/_0288_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2536_  (.A(\hash/CA1/_1533_ ),
    .B(\hash/CA1/_0288_ ),
    .Y(\hash/p4[8] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2537_  (.A(\hash/CA1/_1531_ ),
    .B(\hash/CA1/_1533_ ),
    .Y(\hash/CA1/_0289_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2538_  (.A1(\hash/CA1/_1533_ ),
    .A2(\hash/CA1/_1530_ ),
    .B1(\hash/CA1/_1532_ ),
    .X(\hash/CA1/_0290_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2539_  (.A1(\hash/CA1/_0285_ ),
    .A2(\hash/CA1/_0289_ ),
    .B1_N(\hash/CA1/_0290_ ),
    .Y(\hash/CA1/_0291_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2540_  (.A(\hash/CA1/_1535_ ),
    .B(\hash/CA1/_0291_ ),
    .X(\hash/p4[9] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2541_  (.A(\hash/CA1/_1537_ ),
    .Y(\hash/CA1/_0292_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2542_  (.A1(\hash/CA1/_1535_ ),
    .A2(\hash/CA1/_0290_ ),
    .B1(\hash/CA1/_1534_ ),
    .Y(\hash/CA1/_0293_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2543_  (.A(\hash/CA1/_1526_ ),
    .B(\hash/CA1/_1528_ ),
    .Y(\hash/CA1/_0294_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2544_  (.A(\hash/CA1/_0293_ ),
    .B(\hash/CA1/_0294_ ),
    .Y(\hash/CA1/_0295_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2545_  (.A1(\hash/CA1/_1527_ ),
    .A2(\hash/CA1/_0279_ ),
    .B1(\hash/CA1/_0295_ ),
    .Y(\hash/CA1/_0296_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2546_  (.A(\hash/CA1/_1531_ ),
    .B(\hash/CA1/_1533_ ),
    .C(\hash/CA1/_1535_ ),
    .Y(\hash/CA1/_0297_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2547_  (.A(\hash/CA1/_1529_ ),
    .B(\hash/CA1/_1528_ ),
    .Y(\hash/CA1/_0298_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2548_  (.A1(\hash/CA1/_0297_ ),
    .A2(\hash/CA1/_0298_ ),
    .B1(\hash/CA1/_0293_ ),
    .X(\hash/CA1/_0299_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2549_  (.A(\hash/CA1/_0296_ ),
    .B(\hash/CA1/_0299_ ),
    .Y(\hash/CA1/_0300_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2550_  (.A(\hash/CA1/_0292_ ),
    .B(\hash/CA1/_0300_ ),
    .Y(\hash/p4[10] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2551_  (.A1(\hash/CA1/_1537_ ),
    .A2(\hash/CA1/_1534_ ),
    .B1(\hash/CA1/_1536_ ),
    .X(\hash/CA1/_0301_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2552_  (.A(\hash/CA1/_0292_ ),
    .B(\hash/CA1/_0297_ ),
    .Y(\hash/CA1/_0302_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2553_  (.A1(\hash/CA1/_0283_ ),
    .A2(\hash/CA1/_0284_ ),
    .B1(\hash/CA1/_0302_ ),
    .X(\hash/CA1/_0303_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2554_  (.A(\hash/CA1/_1535_ ),
    .B(\hash/CA1/_1537_ ),
    .C(\hash/CA1/_0290_ ),
    .X(\hash/CA1/_0304_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2555_  (.A(\hash/CA1/_0301_ ),
    .B(\hash/CA1/_0303_ ),
    .C(\hash/CA1/_0304_ ),
    .Y(\hash/CA1/_0305_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2556_  (.A(\hash/CA1/_1539_ ),
    .B(\hash/CA1/_0305_ ),
    .Y(\hash/p4[11] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2557_  (.A(\hash/CA1/_1537_ ),
    .B(\hash/CA1/_1539_ ),
    .Y(\hash/CA1/_0306_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2558_  (.A1(\hash/CA1/_1539_ ),
    .A2(\hash/CA1/_1536_ ),
    .B1(\hash/CA1/_1538_ ),
    .Y(\hash/CA1/_0307_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2559_  (.A1(\hash/CA1/_0296_ ),
    .A2(\hash/CA1/_0299_ ),
    .A3(\hash/CA1/_0306_ ),
    .B1(\hash/CA1/_0307_ ),
    .Y(\hash/CA1/_0308_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2560_  (.A(\hash/CA1/_1541_ ),
    .B(\hash/CA1/_0308_ ),
    .X(\hash/p4[12] ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2561_  (.A(\hash/CA1/_0305_ ),
    .B_N(\hash/CA1/_1539_ ),
    .Y(\hash/CA1/_0309_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2562_  (.A1(\hash/CA1/_1538_ ),
    .A2(\hash/CA1/_0309_ ),
    .B1(\hash/CA1/_1541_ ),
    .X(\hash/CA1/_0310_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2563_  (.A(\hash/CA1/_1540_ ),
    .B(\hash/CA1/_0310_ ),
    .Y(\hash/CA1/_0311_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2564_  (.A(\hash/CA1/_1543_ ),
    .B(\hash/CA1/_0311_ ),
    .Y(\hash/p4[13] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2565_  (.A1(\hash/CA1/_1541_ ),
    .A2(\hash/CA1/_1540_ ),
    .B1(\hash/CA1/_1543_ ),
    .Y(\hash/CA1/_0312_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2566_  (.A_N(\hash/CA1/_1542_ ),
    .B(\hash/CA1/_0312_ ),
    .Y(\hash/CA1/_0313_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2567_  (.A(\hash/CA1/_1540_ ),
    .B(\hash/CA1/_1542_ ),
    .Y(\hash/CA1/_0314_ ));
 sky130_fd_sc_hd__o311ai_1 \hash/CA1/_2568_  (.A1(\hash/CA1/_0296_ ),
    .A2(\hash/CA1/_0299_ ),
    .A3(\hash/CA1/_0306_ ),
    .B1(\hash/CA1/_0314_ ),
    .C1(\hash/CA1/_0307_ ),
    .Y(\hash/CA1/_0315_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2569_  (.A(\hash/CA1/_0313_ ),
    .B(\hash/CA1/_0315_ ),
    .Y(\hash/CA1/_0316_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2570_  (.A(\hash/CA1/_1545_ ),
    .B(\hash/CA1/_0316_ ),
    .Y(\hash/p4[14] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2571_  (.A1(\hash/CA1/_1543_ ),
    .A2(\hash/CA1/_1540_ ),
    .B1(\hash/CA1/_1542_ ),
    .X(\hash/CA1/_0317_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2572_  (.A1(\hash/CA1/_1545_ ),
    .A2(\hash/CA1/_0317_ ),
    .B1(\hash/CA1/_1544_ ),
    .Y(\hash/CA1/_0318_ ));
 sky130_fd_sc_hd__and4_1 \hash/CA1/_2573_  (.A(\hash/CA1/_1539_ ),
    .B(\hash/CA1/_1541_ ),
    .C(\hash/CA1/_1543_ ),
    .D(\hash/CA1/_1545_ ),
    .X(\hash/CA1/_0319_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2574_  (.A1(\hash/CA1/_0301_ ),
    .A2(\hash/CA1/_0303_ ),
    .A3(\hash/CA1/_0304_ ),
    .B1(\hash/CA1/_0319_ ),
    .Y(\hash/CA1/_0320_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2575_  (.A(\hash/CA1/_1541_ ),
    .B(\hash/CA1/_1543_ ),
    .C(\hash/CA1/_1545_ ),
    .D(\hash/CA1/_1538_ ),
    .Y(\hash/CA1/_0321_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2576_  (.A(\hash/CA1/_0318_ ),
    .B(\hash/CA1/_0320_ ),
    .C(\hash/CA1/_0321_ ),
    .Y(\hash/CA1/_0322_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2577_  (.A(\hash/CA1/_1547_ ),
    .B(\hash/CA1/_0322_ ),
    .X(\hash/p4[15] ));
 sky130_fd_sc_hd__a31o_2 \hash/CA1/_2578_  (.A1(\hash/CA1/_1545_ ),
    .A2(\hash/CA1/_0313_ ),
    .A3(\hash/CA1/_0315_ ),
    .B1(\hash/CA1/_1544_ ),
    .X(\hash/CA1/_0323_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2579_  (.A1(\hash/CA1/_1547_ ),
    .A2(\hash/CA1/_0323_ ),
    .B1(\hash/CA1/_1546_ ),
    .Y(\hash/CA1/_0324_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2580_  (.A(\hash/CA1/_1549_ ),
    .B(\hash/CA1/_0324_ ),
    .Y(\hash/p4[16] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2581_  (.A(\hash/CA1/_1549_ ),
    .Y(\hash/CA1/_0325_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2582_  (.A1(\hash/CA1/_1547_ ),
    .A2(\hash/CA1/_0322_ ),
    .B1(\hash/CA1/_1546_ ),
    .Y(\hash/CA1/_0326_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2583_  (.A(\hash/CA1/_0325_ ),
    .B(\hash/CA1/_0326_ ),
    .Y(\hash/CA1/_0327_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2584_  (.A(\hash/CA1/_1548_ ),
    .B(\hash/CA1/_0327_ ),
    .Y(\hash/CA1/_0328_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2585_  (.A(\hash/CA1/_1551_ ),
    .B(\hash/CA1/_0328_ ),
    .Y(\hash/p4[17] ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2586_  (.A1(\hash/CA1/_0325_ ),
    .A2(\hash/CA1/_0324_ ),
    .B1_N(\hash/CA1/_1548_ ),
    .Y(\hash/CA1/_0329_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2587_  (.A1(\hash/CA1/_1551_ ),
    .A2(\hash/CA1/_0329_ ),
    .B1(\hash/CA1/_1550_ ),
    .Y(\hash/CA1/_0330_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2588_  (.A(\hash/CA1/_1553_ ),
    .B(\hash/CA1/_0330_ ),
    .Y(\hash/p4[18] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2589_  (.A1(\hash/CA1/_1547_ ),
    .A2(\hash/CA1/_1546_ ),
    .B1(\hash/CA1/_1549_ ),
    .X(\hash/CA1/_0331_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2590_  (.A1(\hash/CA1/_1548_ ),
    .A2(\hash/CA1/_0331_ ),
    .B1(\hash/CA1/_1551_ ),
    .X(\hash/CA1/_0332_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2591_  (.A1(\hash/CA1/_1550_ ),
    .A2(\hash/CA1/_0332_ ),
    .B1(\hash/CA1/_1553_ ),
    .Y(\hash/CA1/_0333_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2592_  (.A1(\hash/CA1/_1549_ ),
    .A2(\hash/CA1/_1546_ ),
    .B1(\hash/CA1/_1548_ ),
    .Y(\hash/CA1/_0334_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2593_  (.A(\hash/CA1/_0334_ ),
    .B_N(\hash/CA1/_1551_ ),
    .Y(\hash/CA1/_0335_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2594_  (.A1(\hash/CA1/_1550_ ),
    .A2(\hash/CA1/_0335_ ),
    .B1(\hash/CA1/_1553_ ),
    .Y(\hash/CA1/_0336_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2595_  (.A(\hash/CA1/_0322_ ),
    .B_N(\hash/CA1/_0336_ ),
    .Y(\hash/CA1/_0337_ ));
 sky130_fd_sc_hd__o21ba_2 \hash/CA1/_2596_  (.A1(\hash/CA1/_0333_ ),
    .A2(\hash/CA1/_0337_ ),
    .B1_N(\hash/CA1/_1552_ ),
    .X(\hash/CA1/_0338_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2597_  (.A(\hash/CA1/_1555_ ),
    .B(\hash/CA1/_0338_ ),
    .Y(\hash/p4[19] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2598_  (.A(\hash/CA1/_1555_ ),
    .Y(\hash/CA1/_0339_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2599_  (.A1(\hash/CA1/_1555_ ),
    .A2(\hash/CA1/_1552_ ),
    .B1(\hash/CA1/_1554_ ),
    .Y(\hash/CA1/_0340_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2600_  (.A1(\hash/CA1/_0339_ ),
    .A2(\hash/CA1/_0333_ ),
    .B1(\hash/CA1/_0340_ ),
    .Y(\hash/CA1/_0341_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2601_  (.A(\hash/CA1/_0341_ ),
    .Y(\hash/CA1/_0342_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2602_  (.A1(\hash/CA1/_1551_ ),
    .A2(\hash/CA1/_1548_ ),
    .B1(\hash/CA1/_1546_ ),
    .C1(\hash/CA1/_1544_ ),
    .Y(\hash/CA1/_0343_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA1/_2603_  (.A_N(\hash/CA1/_1550_ ),
    .B(\hash/CA1/_0340_ ),
    .C(\hash/CA1/_0343_ ),
    .Y(\hash/CA1/_0344_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_2604_  (.A1(\hash/CA1/_1545_ ),
    .A2(\hash/CA1/_0313_ ),
    .A3(\hash/CA1/_0315_ ),
    .B1(\hash/CA1/_0344_ ),
    .Y(\hash/CA1/_0345_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2605_  (.A(\hash/CA1/_0342_ ),
    .B(\hash/CA1/_0345_ ),
    .Y(\hash/CA1/_0346_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2606_  (.A(\hash/CA1/_1557_ ),
    .B(\hash/CA1/_0346_ ),
    .X(\hash/p4[20] ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2607_  (.A1(\hash/CA1/_0339_ ),
    .A2(\hash/CA1/_0338_ ),
    .B1_N(\hash/CA1/_1554_ ),
    .Y(\hash/CA1/_0347_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2608_  (.A1(\hash/CA1/_1557_ ),
    .A2(\hash/CA1/_0347_ ),
    .B1(\hash/CA1/_1556_ ),
    .Y(\hash/CA1/_0348_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2609_  (.A(\hash/CA1/_1559_ ),
    .B(\hash/CA1/_0348_ ),
    .Y(\hash/p4[21] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2610_  (.A1(\hash/CA1/_1557_ ),
    .A2(\hash/CA1/_0346_ ),
    .B1(\hash/CA1/_1556_ ),
    .X(\hash/CA1/_0349_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2611_  (.A1(\hash/CA1/_1559_ ),
    .A2(\hash/CA1/_0349_ ),
    .B1(\hash/CA1/_1558_ ),
    .Y(\hash/CA1/_0350_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2612_  (.A(\hash/CA1/_1561_ ),
    .B(\hash/CA1/_0350_ ),
    .Y(\hash/p4[22] ));
 sky130_fd_sc_hd__a2111oi_0 \hash/CA1/_2613_  (.A1(\hash/CA1/_1557_ ),
    .A2(\hash/CA1/_1554_ ),
    .B1(\hash/CA1/_1556_ ),
    .C1(\hash/CA1/_1558_ ),
    .D1(\hash/CA1/_1552_ ),
    .Y(\hash/CA1/_0351_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2614_  (.A(\hash/CA1/_0336_ ),
    .B(\hash/CA1/_0351_ ),
    .Y(\hash/CA1/_0352_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2615_  (.A(\hash/CA1/_0322_ ),
    .B(\hash/CA1/_0352_ ),
    .Y(\hash/CA1/_0353_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2616_  (.A1(\hash/CA1/_1555_ ),
    .A2(\hash/CA1/_1554_ ),
    .B1(\hash/CA1/_1557_ ),
    .X(\hash/CA1/_0354_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2617_  (.A1(\hash/CA1/_1556_ ),
    .A2(\hash/CA1/_0354_ ),
    .B1(\hash/CA1/_1559_ ),
    .X(\hash/CA1/_0355_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2618_  (.A1(\hash/CA1/_1558_ ),
    .A2(\hash/CA1/_0355_ ),
    .B1(\hash/CA1/_1561_ ),
    .Y(\hash/CA1/_0356_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2619_  (.A1(\hash/CA1/_0333_ ),
    .A2(\hash/CA1/_0351_ ),
    .B1(\hash/CA1/_0356_ ),
    .X(\hash/CA1/_0357_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2620_  (.A(\hash/CA1/_0353_ ),
    .B(\hash/CA1/_0357_ ),
    .Y(\hash/CA1/_0358_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2621_  (.A(\hash/CA1/_1560_ ),
    .B(\hash/CA1/_0358_ ),
    .Y(\hash/CA1/_0359_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2622_  (.A(\hash/CA1/_1563_ ),
    .B(\hash/CA1/_0359_ ),
    .Y(\hash/p4[23] ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2623_  (.A(\hash/CA1/_1557_ ),
    .B(\hash/CA1/_1559_ ),
    .C(\hash/CA1/_1561_ ),
    .D(\hash/CA1/_0341_ ),
    .Y(\hash/CA1/_0360_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2624_  (.A1(\hash/CA1/_1559_ ),
    .A2(\hash/CA1/_1556_ ),
    .B1(\hash/CA1/_1558_ ),
    .X(\hash/CA1/_0361_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2625_  (.A1(\hash/CA1/_1561_ ),
    .A2(\hash/CA1/_0361_ ),
    .B1(\hash/CA1/_1560_ ),
    .Y(\hash/CA1/_0362_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_2626_  (.A1(\hash/CA1/_0345_ ),
    .A2(\hash/CA1/_0360_ ),
    .B1(\hash/CA1/_0362_ ),
    .Y(\hash/CA1/_0363_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2627_  (.A1(\hash/CA1/_1563_ ),
    .A2(\hash/CA1/_0363_ ),
    .B1(\hash/CA1/_1562_ ),
    .Y(\hash/CA1/_0364_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2628_  (.A(\hash/CA1/_1565_ ),
    .B(\hash/CA1/_0364_ ),
    .Y(\hash/p4[24] ));
 sky130_fd_sc_hd__and2_1 \hash/CA1/_2629_  (.A(\hash/CA1/_1563_ ),
    .B(\hash/CA1/_1565_ ),
    .X(\hash/CA1/_0365_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2630_  (.A(\hash/CA1/_0357_ ),
    .B_N(\hash/CA1/_0365_ ),
    .Y(\hash/CA1/_0366_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2631_  (.A1(\hash/CA1/_0322_ ),
    .A2(\hash/CA1/_0352_ ),
    .B1(\hash/CA1/_0366_ ),
    .Y(\hash/CA1/_0367_ ));
 sky130_fd_sc_hd__a22oi_1 \hash/CA1/_2632_  (.A1(\hash/CA1/_1565_ ),
    .A2(\hash/CA1/_1562_ ),
    .B1(\hash/CA1/_0365_ ),
    .B2(\hash/CA1/_1560_ ),
    .Y(\hash/CA1/_0368_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2633_  (.A(\hash/CA1/_0367_ ),
    .B(\hash/CA1/_0368_ ),
    .Y(\hash/CA1/_0369_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2634_  (.A(\hash/CA1/_1564_ ),
    .B(\hash/CA1/_0369_ ),
    .Y(\hash/CA1/_0370_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2635_  (.A(\hash/CA1/_1567_ ),
    .B(\hash/CA1/_0370_ ),
    .Y(\hash/p4[25] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2636_  (.A(\hash/CA1/_1567_ ),
    .B(\hash/CA1/_1564_ ),
    .Y(\hash/CA1/_0371_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2637_  (.A(\hash/CA1/_1565_ ),
    .B(\hash/CA1/_1567_ ),
    .C(\hash/CA1/_1562_ ),
    .Y(\hash/CA1/_0372_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2638_  (.A(\hash/CA1/_0371_ ),
    .B(\hash/CA1/_0372_ ),
    .Y(\hash/CA1/_0373_ ));
 sky130_fd_sc_hd__a311o_1 \hash/CA1/_2639_  (.A1(\hash/CA1/_1567_ ),
    .A2(\hash/CA1/_0363_ ),
    .A3(\hash/CA1/_0365_ ),
    .B1(\hash/CA1/_0373_ ),
    .C1(\hash/CA1/_1566_ ),
    .X(\hash/CA1/_0374_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2640_  (.A(\hash/CA1/_1569_ ),
    .B(\hash/CA1/_0374_ ),
    .X(\hash/p4[26] ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2641_  (.A(\hash/CA1/_1564_ ),
    .B(\hash/CA1/_1566_ ),
    .C(\hash/CA1/_1568_ ),
    .Y(\hash/CA1/_0375_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_2642_  (.A(\hash/CA1/_1569_ ),
    .B(\hash/CA1/_1568_ ),
    .X(\hash/CA1/_0376_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2643_  (.A1(\hash/CA1/_1567_ ),
    .A2(\hash/CA1/_1566_ ),
    .A3(\hash/CA1/_1568_ ),
    .B1(\hash/CA1/_0376_ ),
    .Y(\hash/CA1/_0377_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_2644_  (.A1(\hash/CA1/_0367_ ),
    .A2(\hash/CA1/_0368_ ),
    .A3(\hash/CA1/_0375_ ),
    .B1(\hash/CA1/_0377_ ),
    .Y(\hash/CA1/_0378_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2645_  (.A(\hash/CA1/_1571_ ),
    .B(\hash/CA1/_0378_ ),
    .X(\hash/p4[27] ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_2646_  (.A1(\hash/CA1/_1567_ ),
    .A2(\hash/CA1/_0363_ ),
    .A3(\hash/CA1/_0365_ ),
    .B1(\hash/CA1/_0373_ ),
    .Y(\hash/CA1/_0379_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2647_  (.A(\hash/CA1/_1566_ ),
    .B(\hash/CA1/_1568_ ),
    .C(\hash/CA1/_1570_ ),
    .Y(\hash/CA1/_0380_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2648_  (.A1(\hash/CA1/_1571_ ),
    .A2(\hash/CA1/_0376_ ),
    .B1(\hash/CA1/_1570_ ),
    .Y(\hash/CA1/_0381_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2649_  (.A1(\hash/CA1/_0379_ ),
    .A2(\hash/CA1/_0380_ ),
    .B1(\hash/CA1/_0381_ ),
    .Y(\hash/CA1/_0382_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2650_  (.A(\hash/CA1/_1573_ ),
    .B(\hash/CA1/_0382_ ),
    .X(\hash/p4[28] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2651_  (.A1(\hash/CA1/_1571_ ),
    .A2(\hash/CA1/_0378_ ),
    .B1(\hash/CA1/_1570_ ),
    .X(\hash/CA1/_0383_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2652_  (.A1(\hash/CA1/_1573_ ),
    .A2(\hash/CA1/_0383_ ),
    .B1(\hash/CA1/_1572_ ),
    .Y(\hash/CA1/_0384_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2653_  (.A(\hash/CA1/_1575_ ),
    .B(\hash/CA1/_0384_ ),
    .Y(\hash/p4[29] ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2654_  (.A(\hash/CA1/_1571_ ),
    .B(\hash/CA1/_1573_ ),
    .C(\hash/CA1/_1575_ ),
    .X(\hash/CA1/_0385_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2655_  (.A1(\hash/CA1/_1571_ ),
    .A2(\hash/CA1/_1568_ ),
    .B1(\hash/CA1/_1570_ ),
    .X(\hash/CA1/_0386_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2656_  (.A1(\hash/CA1/_1573_ ),
    .A2(\hash/CA1/_0386_ ),
    .B1(\hash/CA1/_1572_ ),
    .Y(\hash/CA1/_0387_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2657_  (.A(\hash/CA1/_0387_ ),
    .B_N(\hash/CA1/_1575_ ),
    .Y(\hash/CA1/_0388_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/CA1/_2658_  (.A1(\hash/CA1/_1569_ ),
    .A2(\hash/CA1/_0374_ ),
    .A3(\hash/CA1/_0385_ ),
    .B1(\hash/CA1/_0388_ ),
    .C1(\hash/CA1/_1574_ ),
    .Y(\hash/CA1/_0389_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2659_  (.A(\hash/CA1/_1577_ ),
    .B(\hash/CA1/_0389_ ),
    .Y(\hash/p4[30] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2660_  (.A(\hash/CA1/_1079_ ),
    .Y(\hash/CA1/_1675_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2661_  (.A(\hash/CA1/_1103_ ),
    .Y(\hash/CA1/_1704_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2662_  (.A(\hash/CA1/_1108_ ),
    .Y(\hash/CA1/_1713_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2663_  (.A(\hash/CA1/_1113_ ),
    .Y(\hash/CA1/_1722_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2664_  (.A(\hash/CA1/_1112_ ),
    .Y(\hash/CA1/_1731_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2665_  (.A(\hash/CA1/_1117_ ),
    .Y(\hash/CA1/_1740_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2666_  (.A(\hash/CA1/_1128_ ),
    .Y(\hash/CA1/_1749_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2667_  (.A(\hash/CA1/_1139_ ),
    .Y(\hash/CA1/_1765_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2668_  (.A(\hash/CA1/_1144_ ),
    .Y(\hash/CA1/_1774_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2669_  (.A(\hash/CA1/_1143_ ),
    .Y(\hash/CA1/_1783_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2670_  (.A(\hash/CA1/_1148_ ),
    .Y(\hash/CA1/_1792_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2671_  (.A(\hash/CA1/_1159_ ),
    .Y(\hash/CA1/_1801_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2672_  (.A(\hash/CA1/_1164_ ),
    .Y(\hash/CA1/_1810_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2673_  (.A(\hash/CA1/_1169_ ),
    .Y(\hash/CA1/_1819_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2674_  (.A(\hash/CA1/_1168_ ),
    .Y(\hash/CA1/_1828_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2675_  (.A(\hash/CA1/_1173_ ),
    .Y(\hash/CA1/_1837_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2676_  (.A(\hash/CA1/_1184_ ),
    .Y(\hash/CA1/_1846_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2677_  (.A(\hash/CA1/_1189_ ),
    .Y(\hash/CA1/_1855_ ));
 sky130_fd_sc_hd__a41o_1 \hash/CA1/_2678_  (.A1(\hash/CA1/_1867_ ),
    .A2(\hash/CA1/_0238_ ),
    .A3(\hash/CA1/_0240_ ),
    .A4(\hash/CA1/_0241_ ),
    .B1(\hash/CA1/_1866_ ),
    .X(\hash/CA1/_0390_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2679_  (.A1(\hash/CA1/_1874_ ),
    .A2(\hash/CA1/_0390_ ),
    .B1(\hash/CA1/_1873_ ),
    .Y(\hash/CA1/_0391_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2680_  (.A(\hash/CA1/_1881_ ),
    .B(\hash/CA1/_0391_ ),
    .Y(\hash/CA1/_1209_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2681_  (.A1(\hash/CA1/_1862_ ),
    .A2(\hash/CA1/_1852_ ),
    .B1(\hash/CA1/_1861_ ),
    .X(\hash/CA1/_0392_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2682_  (.A1(\hash/CA1/_1870_ ),
    .A2(\hash/CA1/_0392_ ),
    .B1(\hash/CA1/_1869_ ),
    .Y(\hash/CA1/_0393_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2683_  (.A(\hash/CA1/_0393_ ),
    .B_N(\hash/CA1/_1877_ ),
    .Y(\hash/CA1/_0394_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/CA1/_2684_  (.A1(\hash/CA1/_1853_ ),
    .A2(\hash/CA1/_0223_ ),
    .A3(\hash/CA1/_0252_ ),
    .B1(\hash/CA1/_0394_ ),
    .C1(\hash/CA1/_1876_ ),
    .Y(\hash/CA1/_0395_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2685_  (.A(\hash/CA1/_1884_ ),
    .B(\hash/CA1/_0395_ ),
    .Y(\hash/CA1/_1210_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2686_  (.A(\hash/CA1/_1228_ ),
    .Y(\hash/CA1/_1230_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2687_  (.A(\hash/CA1/_1222_ ),
    .Y(\hash/CA1/_1887_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2688_  (.A(\hash/CA1/_1237_ ),
    .Y(\hash/CA1/_1239_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2689_  (.A(\hash/CA1/_1255_ ),
    .Y(\hash/CA1/_1894_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2690_  (.A(\hash/CA1/_1262_ ),
    .Y(\hash/CA1/_1898_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2691_  (.A(\hash/CA1/_1269_ ),
    .Y(\hash/CA1/_1902_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2692_  (.A(\hash/CA1/_1272_ ),
    .Y(\hash/CA1/_1273_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2693_  (.A(\hash/CA1/_1268_ ),
    .Y(\hash/CA1/_1905_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2694_  (.A(\hash/CA1/_1281_ ),
    .Y(\hash/CA1/_1908_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2695_  (.A(\hash/CA1/_1288_ ),
    .Y(\hash/CA1/_1912_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2696_  (.A(\hash/CA1/_1295_ ),
    .Y(\hash/CA1/_1916_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2697_  (.A(\hash/CA1/_1302_ ),
    .Y(\hash/CA1/_1920_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2698_  (.A(\hash/CA1/_1317_ ),
    .Y(\hash/CA1/_1318_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2699_  (.A(\hash/CA1/_1756_ ),
    .B(\hash/CA1/_0115_ ),
    .Y(\hash/CA1/_1129_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2700_  (.A(\hash/CA1/_1325_ ),
    .Y(\hash/CA1/_1933_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2701_  (.A(\hash/CA1/_1351_ ),
    .Y(\hash/CA1/_1940_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2702_  (.A(\hash/CA1/_1835_ ),
    .B(\hash/CA1/_0191_ ),
    .X(\hash/CA1/_1374_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2703_  (.A(\hash/CA1/_1369_ ),
    .Y(\hash/CA1/_1951_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2704_  (.A(\hash/CA1/_1383_ ),
    .Y(\hash/CA1/_1954_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2705_  (.A(\hash/CA1/_1382_ ),
    .Y(\hash/CA1/_1957_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2706_  (.A(\hash/CA1/_1398_ ),
    .Y(\hash/CA1/_1400_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2707_  (.A(\hash/CA1/_1404_ ),
    .Y(\hash/CA1/_1410_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2708_  (.A(\hash/CA1/_1406_ ),
    .Y(\hash/CA1/_1967_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2709_  (.A(\hash/b[0] ),
    .B(\hash/a[0] ),
    .C(\hash/c[0] ),
    .X(\hash/CA1/_1970_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2710_  (.A(\hash/CA1/_1217_ ),
    .Y(\hash/CA1/_1971_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2711_  (.A(\hash/CA1/_1639_ ),
    .Y(\hash/CA1/_1215_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2712_  (.A(\hash/CA1/_1642_ ),
    .Y(\hash/CA1/_1420_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2713_  (.A1(\hash/CA1/_1415_ ),
    .A2(\hash/CA1/_1434_ ),
    .B1(\hash/CA1/_1433_ ),
    .X(\hash/CA1/_0396_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2714_  (.A1(\hash/CA1/_1437_ ),
    .A2(\hash/CA1/_0396_ ),
    .B1(\hash/CA1/_1436_ ),
    .Y(\hash/CA1/_0397_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2715_  (.A(\hash/CA1/_0397_ ),
    .B_N(\hash/CA1/_1440_ ),
    .Y(\hash/CA1/_0398_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2716_  (.A1(\hash/CA1/_1439_ ),
    .A2(\hash/CA1/_0398_ ),
    .B1(\hash/CA1/_1443_ ),
    .X(\hash/CA1/_0399_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_2717_  (.A(\hash/CA1/_1442_ ),
    .B(\hash/CA1/_1445_ ),
    .X(\hash/CA1/_0400_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA1/_2718_  (.A1(\hash/CA1/_1446_ ),
    .A2(\hash/CA1/_1445_ ),
    .B1(\hash/CA1/_0399_ ),
    .B2(\hash/CA1/_0400_ ),
    .Y(\hash/CA1/_0401_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2719_  (.A(\hash/CA1/_1449_ ),
    .B(\hash/CA1/_1452_ ),
    .C(\hash/CA1/_1455_ ),
    .Y(\hash/CA1/_0402_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2720_  (.A1(\hash/CA1/_1452_ ),
    .A2(\hash/CA1/_1448_ ),
    .B1(\hash/CA1/_1451_ ),
    .X(\hash/CA1/_0403_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2721_  (.A(\hash/CA1/_1455_ ),
    .B(\hash/CA1/_0403_ ),
    .Y(\hash/CA1/_0404_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2722_  (.A1(\hash/CA1/_0401_ ),
    .A2(\hash/CA1/_0402_ ),
    .B1(\hash/CA1/_0404_ ),
    .Y(\hash/CA1/_0405_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2723_  (.A(\hash/CA1/_1454_ ),
    .B(\hash/CA1/_0405_ ),
    .Y(\hash/CA1/_0406_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2724_  (.A(\hash/CA1/_1458_ ),
    .B(\hash/CA1/_0406_ ),
    .Y(\hash/p1[10] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2725_  (.A(\hash/CA1/_1454_ ),
    .Y(\hash/CA1/_0407_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2726_  (.A1(\hash/CA1/_1414_ ),
    .A2(\hash/CA1/_1431_ ),
    .B1(\hash/CA1/_1430_ ),
    .C1(\hash/CA1/_1433_ ),
    .Y(\hash/CA1/_0408_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2727_  (.A1(\hash/CA1/_1434_ ),
    .A2(\hash/CA1/_1433_ ),
    .B1(\hash/CA1/_1437_ ),
    .Y(\hash/CA1/_0409_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2728_  (.A(\hash/CA1/_1436_ ),
    .B(\hash/CA1/_1439_ ),
    .C(\hash/CA1/_1442_ ),
    .Y(\hash/CA1/_0410_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2729_  (.A1(\hash/CA1/_0408_ ),
    .A2(\hash/CA1/_0409_ ),
    .B1(\hash/CA1/_0410_ ),
    .X(\hash/CA1/_0411_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2730_  (.A1(\hash/CA1/_1440_ ),
    .A2(\hash/CA1/_1439_ ),
    .B1(\hash/CA1/_1443_ ),
    .X(\hash/CA1/_0412_ ));
 sky130_fd_sc_hd__o2111ai_1 \hash/CA1/_2731_  (.A1(\hash/CA1/_1442_ ),
    .A2(\hash/CA1/_0412_ ),
    .B1(\hash/CA1/_1446_ ),
    .C1(\hash/CA1/_1449_ ),
    .D1(\hash/CA1/_1452_ ),
    .Y(\hash/CA1/_0413_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2732_  (.A1(\hash/CA1/_1449_ ),
    .A2(\hash/CA1/_1445_ ),
    .B1(\hash/CA1/_1448_ ),
    .X(\hash/CA1/_0414_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2733_  (.A1(\hash/CA1/_1452_ ),
    .A2(\hash/CA1/_0414_ ),
    .B1(\hash/CA1/_1451_ ),
    .Y(\hash/CA1/_0415_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2734_  (.A1(\hash/CA1/_0411_ ),
    .A2(\hash/CA1/_0413_ ),
    .B1(\hash/CA1/_0415_ ),
    .Y(\hash/CA1/_0416_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2735_  (.A(\hash/CA1/_1455_ ),
    .B(\hash/CA1/_0416_ ),
    .Y(\hash/CA1/_0417_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2736_  (.A(\hash/CA1/_0407_ ),
    .B(\hash/CA1/_0417_ ),
    .Y(\hash/CA1/_0418_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2737_  (.A1(\hash/CA1/_1458_ ),
    .A2(\hash/CA1/_0418_ ),
    .B1(\hash/CA1/_1457_ ),
    .Y(\hash/CA1/_0419_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2738_  (.A(\hash/CA1/_1461_ ),
    .B(\hash/CA1/_0419_ ),
    .Y(\hash/p1[11] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2739_  (.A1(\hash/CA1/_1454_ ),
    .A2(\hash/CA1/_0405_ ),
    .B1(\hash/CA1/_1458_ ),
    .Y(\hash/CA1/_0420_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2740_  (.A_N(\hash/CA1/_1457_ ),
    .B(\hash/CA1/_0420_ ),
    .Y(\hash/CA1/_0421_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2741_  (.A1(\hash/CA1/_1461_ ),
    .A2(\hash/CA1/_0421_ ),
    .B1(\hash/CA1/_1460_ ),
    .Y(\hash/CA1/_0422_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2742_  (.A(\hash/CA1/_1464_ ),
    .B(\hash/CA1/_0422_ ),
    .Y(\hash/p1[12] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2743_  (.A1(\hash/CA1/_1461_ ),
    .A2(\hash/CA1/_1457_ ),
    .B1(\hash/CA1/_1460_ ),
    .X(\hash/CA1/_0423_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2744_  (.A1(\hash/CA1/_1464_ ),
    .A2(\hash/CA1/_0423_ ),
    .B1(\hash/CA1/_1463_ ),
    .Y(\hash/CA1/_0424_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2745_  (.A(\hash/CA1/_1458_ ),
    .B(\hash/CA1/_1461_ ),
    .C(\hash/CA1/_1464_ ),
    .X(\hash/CA1/_0425_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2746_  (.A1(\hash/CA1/_1455_ ),
    .A2(\hash/CA1/_1454_ ),
    .B1(\hash/CA1/_0425_ ),
    .Y(\hash/CA1/_0426_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2747_  (.A(\hash/CA1/_0424_ ),
    .B(\hash/CA1/_0426_ ),
    .Y(\hash/CA1/_0427_ ));
 sky130_fd_sc_hd__o2111ai_1 \hash/CA1/_2748_  (.A1(\hash/CA1/_0411_ ),
    .A2(\hash/CA1/_0413_ ),
    .B1(\hash/CA1/_0415_ ),
    .C1(\hash/CA1/_0424_ ),
    .D1(\hash/CA1/_0407_ ),
    .Y(\hash/CA1/_0428_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2749_  (.A(\hash/CA1/_0427_ ),
    .B(\hash/CA1/_0428_ ),
    .Y(\hash/CA1/_0429_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2750_  (.A(\hash/CA1/_1467_ ),
    .B(\hash/CA1/_0429_ ),
    .Y(\hash/p1[13] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2751_  (.A(\hash/CA1/_1454_ ),
    .B(\hash/CA1/_0425_ ),
    .Y(\hash/CA1/_0430_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2752_  (.A(\hash/CA1/_0424_ ),
    .B(\hash/CA1/_0430_ ),
    .Y(\hash/CA1/_0431_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2753_  (.A1(\hash/CA1/_1467_ ),
    .A2(\hash/CA1/_0431_ ),
    .B1(\hash/CA1/_1466_ ),
    .Y(\hash/CA1/_0432_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2754_  (.A(\hash/CA1/_0432_ ),
    .Y(\hash/CA1/_0433_ ));
 sky130_fd_sc_hd__a31o_2 \hash/CA1/_2755_  (.A1(\hash/CA1/_1467_ ),
    .A2(\hash/CA1/_0405_ ),
    .A3(\hash/CA1/_0425_ ),
    .B1(\hash/CA1/_0433_ ),
    .X(\hash/CA1/_0434_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2756_  (.A(\hash/CA1/_1470_ ),
    .B(\hash/CA1/_0434_ ),
    .X(\hash/p1[14] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2757_  (.A1(\hash/CA1/_1470_ ),
    .A2(\hash/CA1/_1466_ ),
    .B1(\hash/CA1/_1469_ ),
    .X(\hash/CA1/_0435_ ));
 sky130_fd_sc_hd__a41oi_2 \hash/CA1/_2758_  (.A1(\hash/CA1/_1467_ ),
    .A2(\hash/CA1/_1470_ ),
    .A3(\hash/CA1/_0427_ ),
    .A4(\hash/CA1/_0428_ ),
    .B1(\hash/CA1/_0435_ ),
    .Y(\hash/CA1/_0436_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2759_  (.A(\hash/CA1/_1473_ ),
    .B(\hash/CA1/_0436_ ),
    .Y(\hash/p1[15] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2760_  (.A1(\hash/CA1/_1470_ ),
    .A2(\hash/CA1/_0434_ ),
    .B1(\hash/CA1/_1469_ ),
    .X(\hash/CA1/_0437_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2761_  (.A1(\hash/CA1/_1473_ ),
    .A2(\hash/CA1/_0437_ ),
    .B1(\hash/CA1/_1472_ ),
    .Y(\hash/CA1/_0438_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2762_  (.A(\hash/CA1/_1476_ ),
    .B(\hash/CA1/_0438_ ),
    .Y(\hash/p1[16] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2763_  (.A(\hash/CA1/_1473_ ),
    .Y(\hash/CA1/_0439_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2764_  (.A1(\hash/CA1/_0439_ ),
    .A2(\hash/CA1/_0436_ ),
    .B1_N(\hash/CA1/_1472_ ),
    .Y(\hash/CA1/_0440_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2765_  (.A1(\hash/CA1/_1476_ ),
    .A2(\hash/CA1/_0440_ ),
    .B1(\hash/CA1/_1475_ ),
    .Y(\hash/CA1/_0441_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2766_  (.A(\hash/CA1/_1479_ ),
    .B(\hash/CA1/_0441_ ),
    .Y(\hash/p1[17] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2767_  (.A(\hash/CA1/_1467_ ),
    .B(\hash/CA1/_0425_ ),
    .Y(\hash/CA1/_0442_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2768_  (.A(\hash/CA1/_1473_ ),
    .B(\hash/CA1/_1476_ ),
    .C(\hash/CA1/_1479_ ),
    .X(\hash/CA1/_0443_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2769_  (.A(\hash/CA1/_1470_ ),
    .B(\hash/CA1/_0443_ ),
    .Y(\hash/CA1/_0444_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2770_  (.A(\hash/CA1/_0442_ ),
    .B(\hash/CA1/_0444_ ),
    .Y(\hash/CA1/_0445_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2771_  (.A1(\hash/CA1/_1473_ ),
    .A2(\hash/CA1/_1469_ ),
    .B1(\hash/CA1/_1472_ ),
    .X(\hash/CA1/_0446_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2772_  (.A1(\hash/CA1/_1476_ ),
    .A2(\hash/CA1/_0446_ ),
    .B1(\hash/CA1/_1475_ ),
    .X(\hash/CA1/_0447_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2773_  (.A1(\hash/CA1/_1479_ ),
    .A2(\hash/CA1/_0447_ ),
    .B1(\hash/CA1/_1478_ ),
    .Y(\hash/CA1/_0448_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2774_  (.A1(\hash/CA1/_0432_ ),
    .A2(\hash/CA1/_0444_ ),
    .B1(\hash/CA1/_0448_ ),
    .Y(\hash/CA1/_0449_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2775_  (.A1(\hash/CA1/_0405_ ),
    .A2(\hash/CA1/_0445_ ),
    .B1(\hash/CA1/_0449_ ),
    .Y(\hash/CA1/_0450_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2776_  (.A(\hash/CA1/_1482_ ),
    .B(\hash/CA1/_0450_ ),
    .Y(\hash/p1[18] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2777_  (.A(\hash/CA1/_1482_ ),
    .B(\hash/CA1/_0443_ ),
    .Y(\hash/CA1/_0451_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2778_  (.A1(\hash/CA1/_1476_ ),
    .A2(\hash/CA1/_1472_ ),
    .B1(\hash/CA1/_1475_ ),
    .X(\hash/CA1/_0452_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2779_  (.A1(\hash/CA1/_1479_ ),
    .A2(\hash/CA1/_0452_ ),
    .B1(\hash/CA1/_1478_ ),
    .X(\hash/CA1/_0453_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2780_  (.A1(\hash/CA1/_1482_ ),
    .A2(\hash/CA1/_0453_ ),
    .B1(\hash/CA1/_1481_ ),
    .X(\hash/CA1/_0454_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2781_  (.A1(\hash/CA1/_0436_ ),
    .A2(\hash/CA1/_0451_ ),
    .B1_N(\hash/CA1/_0454_ ),
    .Y(\hash/CA1/_0455_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2782_  (.A(\hash/CA1/_1485_ ),
    .B(\hash/CA1/_0455_ ),
    .X(\hash/p1[19] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2783_  (.A(\hash/CA1/_1488_ ),
    .Y(\hash/CA1/_0456_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2784_  (.A(\hash/CA1/_1481_ ),
    .B(\hash/CA1/_1484_ ),
    .Y(\hash/CA1/_0457_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2785_  (.A1(\hash/CA1/_1482_ ),
    .A2(\hash/CA1/_1481_ ),
    .B1(\hash/CA1/_1485_ ),
    .X(\hash/CA1/_0458_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2786_  (.A(\hash/CA1/_1484_ ),
    .B(\hash/CA1/_0458_ ),
    .Y(\hash/CA1/_0459_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2787_  (.A1(\hash/CA1/_0450_ ),
    .A2(\hash/CA1/_0457_ ),
    .B1(\hash/CA1/_0459_ ),
    .Y(\hash/CA1/_0460_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2788_  (.A(\hash/CA1/_0456_ ),
    .B(\hash/CA1/_0460_ ),
    .Y(\hash/p1[20] ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_2789_  (.A(\hash/CA1/_1482_ ),
    .B(\hash/CA1/_1485_ ),
    .C(\hash/CA1/_1488_ ),
    .D(\hash/CA1/_0443_ ),
    .Y(\hash/CA1/_0461_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2790_  (.A1(\hash/CA1/_1485_ ),
    .A2(\hash/CA1/_0454_ ),
    .B1(\hash/CA1/_1484_ ),
    .Y(\hash/CA1/_0462_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2791_  (.A(\hash/CA1/_1487_ ),
    .Y(\hash/CA1/_0463_ ));
 sky130_fd_sc_hd__o221ai_1 \hash/CA1/_2792_  (.A1(\hash/CA1/_0436_ ),
    .A2(\hash/CA1/_0461_ ),
    .B1(\hash/CA1/_0462_ ),
    .B2(\hash/CA1/_0456_ ),
    .C1(\hash/CA1/_0463_ ),
    .Y(\hash/CA1/_0464_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2793_  (.A(\hash/CA1/_1491_ ),
    .B(\hash/CA1/_0464_ ),
    .X(\hash/p1[21] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2794_  (.A1(\hash/CA1/_1491_ ),
    .A2(\hash/CA1/_1487_ ),
    .B1(\hash/CA1/_1490_ ),
    .X(\hash/CA1/_0465_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_2795_  (.A1(\hash/CA1/_1488_ ),
    .A2(\hash/CA1/_1491_ ),
    .A3(\hash/CA1/_0460_ ),
    .B1(\hash/CA1/_0465_ ),
    .Y(\hash/CA1/_0466_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2796_  (.A(\hash/CA1/_1494_ ),
    .B(\hash/CA1/_0466_ ),
    .Y(\hash/p1[22] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2797_  (.A(\hash/CA1/_1487_ ),
    .B(\hash/CA1/_1490_ ),
    .Y(\hash/CA1/_0467_ ));
 sky130_fd_sc_hd__o221ai_1 \hash/CA1/_2798_  (.A1(\hash/CA1/_0436_ ),
    .A2(\hash/CA1/_0461_ ),
    .B1(\hash/CA1/_0462_ ),
    .B2(\hash/CA1/_0456_ ),
    .C1(\hash/CA1/_0467_ ),
    .Y(\hash/CA1/_0468_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2799_  (.A(\hash/CA1/_1494_ ),
    .Y(\hash/CA1/_0469_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2800_  (.A(\hash/CA1/_1491_ ),
    .B(\hash/CA1/_1490_ ),
    .Y(\hash/CA1/_0470_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2801_  (.A(\hash/CA1/_0469_ ),
    .B(\hash/CA1/_0470_ ),
    .Y(\hash/CA1/_0471_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2802_  (.A1(\hash/CA1/_0468_ ),
    .A2(\hash/CA1/_0471_ ),
    .B1(\hash/CA1/_1493_ ),
    .Y(\hash/CA1/_0472_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2803_  (.A(\hash/CA1/_1497_ ),
    .B(\hash/CA1/_0472_ ),
    .Y(\hash/p1[23] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2804_  (.A(\hash/CA1/_1497_ ),
    .Y(\hash/CA1/_0473_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2805_  (.A(\hash/CA1/_1488_ ),
    .B(\hash/CA1/_1491_ ),
    .Y(\hash/CA1/_0474_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2806_  (.A(\hash/CA1/_0469_ ),
    .B(\hash/CA1/_0473_ ),
    .C(\hash/CA1/_0474_ ),
    .Y(\hash/CA1/_0475_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2807_  (.A1(\hash/CA1/_1494_ ),
    .A2(\hash/CA1/_0465_ ),
    .B1(\hash/CA1/_1493_ ),
    .Y(\hash/CA1/_0476_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2808_  (.A1(\hash/CA1/_0473_ ),
    .A2(\hash/CA1/_0476_ ),
    .B1_N(\hash/CA1/_1496_ ),
    .Y(\hash/CA1/_0477_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2809_  (.A1(\hash/CA1/_0460_ ),
    .A2(\hash/CA1/_0475_ ),
    .B1(\hash/CA1/_0477_ ),
    .Y(\hash/CA1/_0478_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2810_  (.A(\hash/CA1/_1500_ ),
    .B(\hash/CA1/_0478_ ),
    .Y(\hash/p1[24] ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2811_  (.A1(\hash/CA1/_0473_ ),
    .A2(\hash/CA1/_0472_ ),
    .B1_N(\hash/CA1/_1496_ ),
    .Y(\hash/CA1/_0479_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2812_  (.A1(\hash/CA1/_1500_ ),
    .A2(\hash/CA1/_0479_ ),
    .B1(\hash/CA1/_1499_ ),
    .Y(\hash/CA1/_0480_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2813_  (.A(\hash/CA1/_1503_ ),
    .B(\hash/CA1/_0480_ ),
    .Y(\hash/p1[25] ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2814_  (.A(\hash/CA1/_1497_ ),
    .B(\hash/CA1/_1500_ ),
    .C(\hash/CA1/_1503_ ),
    .Y(\hash/CA1/_0481_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2815_  (.A(\hash/CA1/_0469_ ),
    .B(\hash/CA1/_0474_ ),
    .C(\hash/CA1/_0481_ ),
    .Y(\hash/CA1/_0482_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2816_  (.A1(\hash/CA1/_1500_ ),
    .A2(\hash/CA1/_0477_ ),
    .B1(\hash/CA1/_1499_ ),
    .X(\hash/CA1/_0483_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2817_  (.A1(\hash/CA1/_1503_ ),
    .A2(\hash/CA1/_0483_ ),
    .B1(\hash/CA1/_1502_ ),
    .X(\hash/CA1/_0484_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2818_  (.A1(\hash/CA1/_0460_ ),
    .A2(\hash/CA1/_0482_ ),
    .B1(\hash/CA1/_0484_ ),
    .Y(\hash/CA1/_0485_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2819_  (.A(\hash/CA1/_1506_ ),
    .B(\hash/CA1/_0485_ ),
    .Y(\hash/p1[26] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2820_  (.A1(\hash/CA1/_1500_ ),
    .A2(\hash/CA1/_1496_ ),
    .B1(\hash/CA1/_1499_ ),
    .X(\hash/CA1/_0486_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2821_  (.A1(\hash/CA1/_1503_ ),
    .A2(\hash/CA1/_0486_ ),
    .B1(\hash/CA1/_1502_ ),
    .Y(\hash/CA1/_0487_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_2822_  (.A1(\hash/CA1/_0472_ ),
    .A2(\hash/CA1/_0481_ ),
    .B1(\hash/CA1/_0487_ ),
    .Y(\hash/CA1/_0488_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2823_  (.A1(\hash/CA1/_1506_ ),
    .A2(\hash/CA1/_0488_ ),
    .B1(\hash/CA1/_1505_ ),
    .Y(\hash/CA1/_0489_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2824_  (.A(\hash/CA1/_1509_ ),
    .B(\hash/CA1/_0489_ ),
    .Y(\hash/p1[27] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2825_  (.A1(\hash/CA1/_1506_ ),
    .A2(\hash/CA1/_1505_ ),
    .B1(\hash/CA1/_1509_ ),
    .Y(\hash/CA1/_0490_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2826_  (.A(\hash/CA1/_1512_ ),
    .B(\hash/CA1/_0490_ ),
    .Y(\hash/CA1/_0491_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2827_  (.A(\hash/CA1/_0460_ ),
    .B(\hash/CA1/_0482_ ),
    .C(\hash/CA1/_0491_ ),
    .Y(\hash/CA1/_0492_ ));
 sky130_fd_sc_hd__or4b_2 \hash/CA1/_2828_  (.A(\hash/CA1/_1505_ ),
    .B(\hash/CA1/_1508_ ),
    .C(\hash/CA1/_0484_ ),
    .D_N(\hash/CA1/_1512_ ),
    .X(\hash/CA1/_0493_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2829_  (.A1(\hash/CA1/_0460_ ),
    .A2(\hash/CA1/_0482_ ),
    .B1(\hash/CA1/_0493_ ),
    .X(\hash/CA1/_0494_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA1/_2830_  (.A_N(\hash/CA1/_1508_ ),
    .B(\hash/CA1/_0490_ ),
    .C(\hash/CA1/_1512_ ),
    .Y(\hash/CA1/_0495_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA1/_2831_  (.A_N(\hash/CA1/_1512_ ),
    .B(\hash/CA1/_1505_ ),
    .C(\hash/CA1/_1509_ ),
    .Y(\hash/CA1/_0496_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2832_  (.A_N(\hash/CA1/_1512_ ),
    .B(\hash/CA1/_1508_ ),
    .Y(\hash/CA1/_0497_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2833_  (.A(\hash/CA1/_0495_ ),
    .B(\hash/CA1/_0496_ ),
    .C(\hash/CA1/_0497_ ),
    .Y(\hash/CA1/_0498_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2834_  (.A1(\hash/CA1/_0484_ ),
    .A2(\hash/CA1/_0491_ ),
    .B1(\hash/CA1/_0498_ ),
    .Y(\hash/CA1/_0499_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2835_  (.A(\hash/CA1/_0492_ ),
    .B(\hash/CA1/_0494_ ),
    .C(\hash/CA1/_0499_ ),
    .Y(\hash/p1[28] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2836_  (.A(\hash/CA1/_1511_ ),
    .Y(\hash/CA1/_0500_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2837_  (.A1(\hash/CA1/_1509_ ),
    .A2(\hash/CA1/_1508_ ),
    .B1(\hash/CA1/_1512_ ),
    .Y(\hash/CA1/_0501_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2838_  (.A(\hash/CA1/_1508_ ),
    .B(\hash/CA1/_1511_ ),
    .Y(\hash/CA1/_0502_ ));
 sky130_fd_sc_hd__a22oi_1 \hash/CA1/_2839_  (.A1(\hash/CA1/_0500_ ),
    .A2(\hash/CA1/_0501_ ),
    .B1(\hash/CA1/_0502_ ),
    .B2(\hash/CA1/_0489_ ),
    .Y(\hash/CA1/_0503_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2840_  (.A(\hash/CA1/_1515_ ),
    .B(\hash/CA1/_0503_ ),
    .X(\hash/p1[29] ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2841_  (.A(\hash/CA1/_1415_ ),
    .B(\hash/CA1/_1434_ ),
    .X(\hash/p1[2] ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2842_  (.A(\hash/CA1/_1509_ ),
    .B(\hash/CA1/_1512_ ),
    .C(\hash/CA1/_1515_ ),
    .X(\hash/CA1/_0504_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA1/_2843_  (.A(\hash/CA1/_1506_ ),
    .B(\hash/CA1/_0504_ ),
    .X(\hash/CA1/_0505_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2844_  (.A(\hash/CA1/_1512_ ),
    .B(\hash/CA1/_1508_ ),
    .Y(\hash/CA1/_0506_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2845_  (.A(\hash/CA1/_0500_ ),
    .B(\hash/CA1/_0506_ ),
    .Y(\hash/CA1/_0507_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA1/_2846_  (.A1(\hash/CA1/_1515_ ),
    .A2(\hash/CA1/_0507_ ),
    .B1(\hash/CA1/_0504_ ),
    .B2(\hash/CA1/_1505_ ),
    .C1(\hash/CA1/_1514_ ),
    .Y(\hash/CA1/_0508_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2847_  (.A(\hash/CA1/_0484_ ),
    .B(\hash/CA1/_0505_ ),
    .Y(\hash/CA1/_0509_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2848_  (.A(\hash/CA1/_0508_ ),
    .B(\hash/CA1/_0509_ ),
    .Y(\hash/CA1/_0510_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_2849_  (.A1(\hash/CA1/_0460_ ),
    .A2(\hash/CA1/_0482_ ),
    .A3(\hash/CA1/_0505_ ),
    .B1(\hash/CA1/_0510_ ),
    .Y(\hash/CA1/_0511_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2850_  (.A(\hash/CA1/_1518_ ),
    .B(\hash/CA1/_0511_ ),
    .Y(\hash/p1[30] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA1/_2851_  (.A(\hash/b[31] ),
    .B(\hash/a[31] ),
    .C(\hash/c[31] ),
    .X(\hash/CA1/_0512_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2852_  (.A(\hash/CA1/s0[31] ),
    .B(\hash/CA1/_0512_ ),
    .X(\hash/CA1/_0513_ ));
 sky130_fd_sc_hd__a21bo_2 \hash/CA1/_2853_  (.A1(\hash/CA1/_0488_ ),
    .A2(\hash/CA1/_0505_ ),
    .B1_N(\hash/CA1/_0508_ ),
    .X(\hash/CA1/_0514_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2854_  (.A1(\hash/CA1/_1518_ ),
    .A2(\hash/CA1/_0514_ ),
    .B1(\hash/CA1/_1517_ ),
    .Y(\hash/CA1/_0515_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2855_  (.A(\hash/CA1/_0513_ ),
    .B(\hash/CA1/_0515_ ),
    .Y(\hash/p1[31] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2856_  (.A(\hash/CA1/_0408_ ),
    .B(\hash/CA1/_0409_ ),
    .Y(\hash/CA1/_0516_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2857_  (.A1(\hash/CA1/_1414_ ),
    .A2(\hash/CA1/_1431_ ),
    .B1(\hash/CA1/_1430_ ),
    .X(\hash/CA1/_0517_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2858_  (.A1(\hash/CA1/_1434_ ),
    .A2(\hash/CA1/_0517_ ),
    .B1(\hash/CA1/_1433_ ),
    .C1(\hash/CA1/_1437_ ),
    .Y(\hash/CA1/_0518_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2859_  (.A(\hash/CA1/_0516_ ),
    .B(\hash/CA1/_0518_ ),
    .Y(\hash/p1[3] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2860_  (.A(\hash/CA1/_1440_ ),
    .B(\hash/CA1/_0397_ ),
    .Y(\hash/p1[4] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2861_  (.A1(\hash/CA1/_1436_ ),
    .A2(\hash/CA1/_0516_ ),
    .B1(\hash/CA1/_1440_ ),
    .X(\hash/CA1/_0519_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2862_  (.A(\hash/CA1/_1439_ ),
    .B(\hash/CA1/_0519_ ),
    .Y(\hash/CA1/_0520_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2863_  (.A(\hash/CA1/_1443_ ),
    .B(\hash/CA1/_0520_ ),
    .Y(\hash/p1[5] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2864_  (.A(\hash/CA1/_1442_ ),
    .B(\hash/CA1/_0399_ ),
    .Y(\hash/CA1/_0521_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2865_  (.A(\hash/CA1/_1446_ ),
    .B(\hash/CA1/_0521_ ),
    .Y(\hash/p1[6] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2866_  (.A1(\hash/CA1/_1442_ ),
    .A2(\hash/CA1/_0412_ ),
    .B1(\hash/CA1/_1446_ ),
    .Y(\hash/CA1/_0522_ ));
 sky130_fd_sc_hd__o21ba_2 \hash/CA1/_2867_  (.A1(\hash/CA1/_0411_ ),
    .A2(\hash/CA1/_0522_ ),
    .B1_N(\hash/CA1/_1445_ ),
    .X(\hash/CA1/_0523_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2868_  (.A(\hash/CA1/_1449_ ),
    .B(\hash/CA1/_0523_ ),
    .Y(\hash/p1[7] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2869_  (.A(\hash/CA1/_1449_ ),
    .Y(\hash/CA1/_0524_ ));
 sky130_fd_sc_hd__o21ba_2 \hash/CA1/_2870_  (.A1(\hash/CA1/_0524_ ),
    .A2(\hash/CA1/_0401_ ),
    .B1_N(\hash/CA1/_1448_ ),
    .X(\hash/CA1/_0525_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2871_  (.A(\hash/CA1/_1452_ ),
    .B(\hash/CA1/_0525_ ),
    .Y(\hash/p1[8] ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2872_  (.A(\hash/CA1/_1455_ ),
    .B(\hash/CA1/_0416_ ),
    .X(\hash/p1[9] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2873_  (.A1(\hash/CA1/_1904_ ),
    .A2(\hash/CA1/_1903_ ),
    .B1(\hash/CA1/_1907_ ),
    .X(\hash/CA1/_0526_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2874_  (.A1(\hash/CA1/_1906_ ),
    .A2(\hash/CA1/_0526_ ),
    .B1(\hash/CA1/_1910_ ),
    .X(\hash/CA1/_0527_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2875_  (.A(\hash/CA1/_1900_ ),
    .Y(\hash/CA1/_0528_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2876_  (.A(\hash/CA1/_1893_ ),
    .Y(\hash/CA1/_0529_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2877_  (.A1(\hash/CA1/_1974_ ),
    .A2(\hash/CA1/_1889_ ),
    .B1(\hash/CA1/_1888_ ),
    .X(\hash/CA1/_0530_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2878_  (.A1(\hash/CA1/_1891_ ),
    .A2(\hash/CA1/_0530_ ),
    .B1(\hash/CA1/_1890_ ),
    .Y(\hash/CA1/_0531_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2879_  (.A1(\hash/CA1/_0529_ ),
    .A2(\hash/CA1/_0531_ ),
    .B1_N(\hash/CA1/_1892_ ),
    .Y(\hash/CA1/_0532_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2880_  (.A1(\hash/CA1/_1896_ ),
    .A2(\hash/CA1/_0532_ ),
    .B1(\hash/CA1/_1895_ ),
    .Y(\hash/CA1/_0533_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2881_  (.A(\hash/CA1/_1899_ ),
    .B(\hash/CA1/_1903_ ),
    .C(\hash/CA1/_1906_ ),
    .Y(\hash/CA1/_0534_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2882_  (.A1(\hash/CA1/_0528_ ),
    .A2(\hash/CA1/_0533_ ),
    .B1(\hash/CA1/_0534_ ),
    .Y(\hash/CA1/_0535_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2883_  (.A1(\hash/CA1/_0527_ ),
    .A2(\hash/CA1/_0535_ ),
    .B1(\hash/CA1/_1909_ ),
    .Y(\hash/CA1/_0536_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2884_  (.A(\hash/CA1/_1914_ ),
    .B(\hash/CA1/_0536_ ),
    .Y(\hash/p2[10] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2885_  (.A1(\hash/CA1/_1914_ ),
    .A2(\hash/CA1/_1909_ ),
    .B1(\hash/CA1/_1913_ ),
    .X(\hash/CA1/_0537_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2886_  (.A1(\hash/CA1/_1914_ ),
    .A2(\hash/CA1/_0527_ ),
    .B1(\hash/CA1/_0537_ ),
    .X(\hash/CA1/_0538_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2887_  (.A(\hash/CA1/_1418_ ),
    .B_N(\hash/CA1/_1891_ ),
    .Y(\hash/CA1/_0539_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_2888_  (.A1(\hash/CA1/_1890_ ),
    .A2(\hash/CA1/_0539_ ),
    .B1(\hash/CA1/_1893_ ),
    .Y(\hash/CA1/_0540_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2889_  (.A(\hash/CA1/_1900_ ),
    .B(\hash/CA1/_1896_ ),
    .Y(\hash/CA1/_0541_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2890_  (.A1(\hash/CA1/_1896_ ),
    .A2(\hash/CA1/_1892_ ),
    .B1(\hash/CA1/_1895_ ),
    .X(\hash/CA1/_0542_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2891_  (.A(\hash/CA1/_1900_ ),
    .B(\hash/CA1/_0542_ ),
    .Y(\hash/CA1/_0543_ ));
 sky130_fd_sc_hd__nor4_1 \hash/CA1/_2892_  (.A(\hash/CA1/_1899_ ),
    .B(\hash/CA1/_1903_ ),
    .C(\hash/CA1/_1906_ ),
    .D(\hash/CA1/_0537_ ),
    .Y(\hash/CA1/_0544_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_2893_  (.A1(\hash/CA1/_0540_ ),
    .A2(\hash/CA1/_0541_ ),
    .B1(\hash/CA1/_0543_ ),
    .C1(\hash/CA1/_0544_ ),
    .Y(\hash/CA1/_0545_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2894_  (.A(\hash/CA1/_0538_ ),
    .B(\hash/CA1/_0545_ ),
    .Y(\hash/CA1/_0546_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2895_  (.A(\hash/CA1/_1918_ ),
    .B(\hash/CA1/_0546_ ),
    .Y(\hash/p2[11] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2896_  (.A(\hash/CA1/_1914_ ),
    .Y(\hash/CA1/_0547_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2897_  (.A1(\hash/CA1/_0547_ ),
    .A2(\hash/CA1/_0536_ ),
    .B1_N(\hash/CA1/_1913_ ),
    .Y(\hash/CA1/_0548_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2898_  (.A1(\hash/CA1/_1918_ ),
    .A2(\hash/CA1/_0548_ ),
    .B1(\hash/CA1/_1917_ ),
    .Y(\hash/CA1/_0549_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2899_  (.A(\hash/CA1/_1922_ ),
    .B(\hash/CA1/_0549_ ),
    .Y(\hash/p2[12] ));
 sky130_fd_sc_hd__a31o_2 \hash/CA1/_2900_  (.A1(\hash/CA1/_1918_ ),
    .A2(\hash/CA1/_0538_ ),
    .A3(\hash/CA1/_0545_ ),
    .B1(\hash/CA1/_1917_ ),
    .X(\hash/CA1/_0550_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2901_  (.A1(\hash/CA1/_1922_ ),
    .A2(\hash/CA1/_0550_ ),
    .B1(\hash/CA1/_1921_ ),
    .Y(\hash/CA1/_0551_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2902_  (.A(\hash/CA1/_1925_ ),
    .B(\hash/CA1/_0551_ ),
    .Y(\hash/p2[13] ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2903_  (.A(\hash/CA1/_1918_ ),
    .B(\hash/CA1/_1922_ ),
    .C(\hash/CA1/_1925_ ),
    .X(\hash/CA1/_0552_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_2904_  (.A(\hash/CA1/_1914_ ),
    .B(\hash/CA1/_0527_ ),
    .C(\hash/CA1/_0552_ ),
    .X(\hash/CA1/_0553_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2905_  (.A1(\hash/CA1/_1918_ ),
    .A2(\hash/CA1/_1913_ ),
    .B1(\hash/CA1/_1917_ ),
    .X(\hash/CA1/_0554_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2906_  (.A1(\hash/CA1/_1922_ ),
    .A2(\hash/CA1/_0554_ ),
    .B1(\hash/CA1/_1921_ ),
    .X(\hash/CA1/_0555_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2907_  (.A1(\hash/CA1/_1925_ ),
    .A2(\hash/CA1/_0555_ ),
    .B1(\hash/CA1/_1924_ ),
    .Y(\hash/CA1/_0556_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2908_  (.A(\hash/CA1/_1914_ ),
    .B(\hash/CA1/_1909_ ),
    .C(\hash/CA1/_0552_ ),
    .Y(\hash/CA1/_0557_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2909_  (.A(\hash/CA1/_0556_ ),
    .B(\hash/CA1/_0557_ ),
    .Y(\hash/CA1/_0558_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2910_  (.A1(\hash/CA1/_0535_ ),
    .A2(\hash/CA1/_0553_ ),
    .B1(\hash/CA1/_0558_ ),
    .X(\hash/CA1/_0559_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2911_  (.A(\hash/CA1/_1927_ ),
    .B(\hash/CA1/_0559_ ),
    .X(\hash/p2[14] ));
 sky130_fd_sc_hd__a211o_1 \hash/CA1/_2912_  (.A1(\hash/CA1/_1927_ ),
    .A2(\hash/CA1/_1924_ ),
    .B1(\hash/CA1/_1926_ ),
    .C1(\hash/CA1/_1921_ ),
    .X(\hash/CA1/_0560_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_2913_  (.A1(\hash/CA1/_1922_ ),
    .A2(\hash/CA1/_1921_ ),
    .B1(\hash/CA1/_1927_ ),
    .C1(\hash/CA1/_1925_ ),
    .Y(\hash/CA1/_0561_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2914_  (.A1(\hash/CA1/_1927_ ),
    .A2(\hash/CA1/_1924_ ),
    .B1(\hash/CA1/_1926_ ),
    .Y(\hash/CA1/_0562_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2915_  (.A(\hash/CA1/_0561_ ),
    .B(\hash/CA1/_0562_ ),
    .Y(\hash/CA1/_0563_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2916_  (.A1(\hash/CA1/_0550_ ),
    .A2(\hash/CA1/_0560_ ),
    .B1(\hash/CA1/_0563_ ),
    .Y(\hash/CA1/_0564_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2917_  (.A(\hash/CA1/_1929_ ),
    .B(\hash/CA1/_0564_ ),
    .Y(\hash/p2[15] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2918_  (.A1(\hash/CA1/_1927_ ),
    .A2(\hash/CA1/_1926_ ),
    .B1(\hash/CA1/_1929_ ),
    .Y(\hash/CA1/_0565_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2919_  (.A_N(\hash/CA1/_1928_ ),
    .B(\hash/CA1/_0565_ ),
    .Y(\hash/CA1/_0566_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2920_  (.A1(\hash/CA1/_1926_ ),
    .A2(\hash/CA1/_1928_ ),
    .A3(\hash/CA1/_0559_ ),
    .B1(\hash/CA1/_0566_ ),
    .Y(\hash/CA1/_0567_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2921_  (.A(\hash/CA1/_1932_ ),
    .B(\hash/CA1/_0567_ ),
    .Y(\hash/p2[16] ));
 sky130_fd_sc_hd__a311oi_2 \hash/CA1/_2922_  (.A1(\hash/CA1/_1918_ ),
    .A2(\hash/CA1/_0538_ ),
    .A3(\hash/CA1/_0545_ ),
    .B1(\hash/CA1/_0560_ ),
    .C1(\hash/CA1/_1917_ ),
    .Y(\hash/CA1/_0568_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2923_  (.A(\hash/CA1/_1929_ ),
    .B(\hash/CA1/_1932_ ),
    .C(\hash/CA1/_0563_ ),
    .Y(\hash/CA1/_0569_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2924_  (.A1(\hash/CA1/_1932_ ),
    .A2(\hash/CA1/_1928_ ),
    .B1(\hash/CA1/_1931_ ),
    .Y(\hash/CA1/_0570_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2925_  (.A1(\hash/CA1/_0568_ ),
    .A2(\hash/CA1/_0569_ ),
    .B1(\hash/CA1/_0570_ ),
    .Y(\hash/CA1/_0571_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2926_  (.A(\hash/CA1/_1935_ ),
    .B(\hash/CA1/_0571_ ),
    .X(\hash/p2[17] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2927_  (.A(\hash/CA1/_1932_ ),
    .Y(\hash/CA1/_0572_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_2928_  (.A1(\hash/CA1/_0572_ ),
    .A2(\hash/CA1/_0567_ ),
    .B1_N(\hash/CA1/_1931_ ),
    .Y(\hash/CA1/_0573_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2929_  (.A1(\hash/CA1/_1935_ ),
    .A2(\hash/CA1/_0573_ ),
    .B1(\hash/CA1/_1934_ ),
    .Y(\hash/CA1/_0574_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2930_  (.A(\hash/CA1/_1937_ ),
    .B(\hash/CA1/_0574_ ),
    .Y(\hash/p2[18] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2931_  (.A(\hash/CA1/_1935_ ),
    .B(\hash/CA1/_1937_ ),
    .Y(\hash/CA1/_0575_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2932_  (.A(\hash/CA1/_0570_ ),
    .B(\hash/CA1/_0575_ ),
    .Y(\hash/CA1/_0576_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2933_  (.A1(\hash/CA1/_1937_ ),
    .A2(\hash/CA1/_1934_ ),
    .B1(\hash/CA1/_1936_ ),
    .C1(\hash/CA1/_0576_ ),
    .Y(\hash/CA1/_0577_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2934_  (.A1(\hash/CA1/_0569_ ),
    .A2(\hash/CA1/_0575_ ),
    .B1(\hash/CA1/_0577_ ),
    .X(\hash/CA1/_0578_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2935_  (.A1(\hash/CA1/_0568_ ),
    .A2(\hash/CA1/_0577_ ),
    .B1(\hash/CA1/_0578_ ),
    .Y(\hash/CA1/_0579_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2936_  (.A(\hash/CA1/_1939_ ),
    .B(\hash/CA1/_0579_ ),
    .X(\hash/p2[19] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2937_  (.A(\hash/CA1/_0572_ ),
    .B(\hash/CA1/_0575_ ),
    .Y(\hash/CA1/_0580_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2938_  (.A1(\hash/CA1/_1935_ ),
    .A2(\hash/CA1/_1931_ ),
    .B1(\hash/CA1/_1934_ ),
    .X(\hash/CA1/_0581_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2939_  (.A1(\hash/CA1/_1937_ ),
    .A2(\hash/CA1/_0581_ ),
    .B1(\hash/CA1/_1936_ ),
    .Y(\hash/CA1/_0582_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2940_  (.A(\hash/CA1/_1926_ ),
    .B(\hash/CA1/_1928_ ),
    .Y(\hash/CA1/_0583_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2941_  (.A(\hash/CA1/_0583_ ),
    .B(\hash/CA1/_0575_ ),
    .Y(\hash/CA1/_0584_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2942_  (.A(\hash/CA1/_1932_ ),
    .B(\hash/CA1/_0566_ ),
    .C(\hash/CA1/_0584_ ),
    .Y(\hash/CA1/_0585_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2943_  (.A(\hash/CA1/_0582_ ),
    .B(\hash/CA1/_0585_ ),
    .Y(\hash/CA1/_0586_ ));
 sky130_fd_sc_hd__a31o_2 \hash/CA1/_2944_  (.A1(\hash/CA1/_0559_ ),
    .A2(\hash/CA1/_0566_ ),
    .A3(\hash/CA1/_0580_ ),
    .B1(\hash/CA1/_0586_ ),
    .X(\hash/CA1/_0587_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2945_  (.A1(\hash/CA1/_1939_ ),
    .A2(\hash/CA1/_0587_ ),
    .B1(\hash/CA1/_1938_ ),
    .Y(\hash/CA1/_0588_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2946_  (.A(\hash/CA1/_1942_ ),
    .B(\hash/CA1/_0588_ ),
    .Y(\hash/p2[20] ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2947_  (.A(\hash/CA1/_1939_ ),
    .B(\hash/CA1/_1942_ ),
    .C(\hash/CA1/_1945_ ),
    .Y(\hash/CA1/_0589_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2948_  (.A1(\hash/CA1/_0568_ ),
    .A2(\hash/CA1/_0577_ ),
    .B1(\hash/CA1/_0578_ ),
    .C1(\hash/CA1/_0589_ ),
    .Y(\hash/CA1/_0590_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2949_  (.A(\hash/CA1/_1945_ ),
    .B(\hash/CA1/_1941_ ),
    .Y(\hash/CA1/_0591_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2950_  (.A(\hash/CA1/_1942_ ),
    .B(\hash/CA1/_1945_ ),
    .C(\hash/CA1/_1938_ ),
    .Y(\hash/CA1/_0592_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2951_  (.A(\hash/CA1/_0591_ ),
    .B(\hash/CA1/_0592_ ),
    .Y(\hash/CA1/_0593_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2952_  (.A1(\hash/CA1/_1939_ ),
    .A2(\hash/CA1/_0579_ ),
    .B1(\hash/CA1/_1938_ ),
    .X(\hash/CA1/_0594_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2953_  (.A1(\hash/CA1/_1942_ ),
    .A2(\hash/CA1/_0594_ ),
    .B1(\hash/CA1/_1941_ ),
    .C1(\hash/CA1/_1945_ ),
    .Y(\hash/CA1/_0595_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2954_  (.A(\hash/CA1/_0590_ ),
    .B(\hash/CA1/_0593_ ),
    .C(\hash/CA1/_0595_ ),
    .Y(\hash/p2[21] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2955_  (.A(\hash/CA1/_1942_ ),
    .B(\hash/CA1/_1945_ ),
    .Y(\hash/CA1/_0596_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2956_  (.A1(\hash/CA1/_1945_ ),
    .A2(\hash/CA1/_1941_ ),
    .B1(\hash/CA1/_1944_ ),
    .Y(\hash/CA1/_0597_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2957_  (.A1(\hash/CA1/_0588_ ),
    .A2(\hash/CA1/_0596_ ),
    .B1(\hash/CA1/_0597_ ),
    .Y(\hash/CA1/_0598_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_2958_  (.A(\hash/CA1/_1947_ ),
    .B(\hash/CA1/_0598_ ),
    .X(\hash/p2[22] ));
 sky130_fd_sc_hd__or3_1 \hash/CA1/_2959_  (.A(\hash/CA1/_1944_ ),
    .B(\hash/CA1/_0590_ ),
    .C(\hash/CA1/_0593_ ),
    .X(\hash/CA1/_0599_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2960_  (.A1(\hash/CA1/_1947_ ),
    .A2(\hash/CA1/_0599_ ),
    .B1(\hash/CA1/_1946_ ),
    .Y(\hash/CA1/_0600_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2961_  (.A(\hash/CA1/_1950_ ),
    .B(\hash/CA1/_0600_ ),
    .Y(\hash/p2[23] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2962_  (.A(\hash/CA1/_1953_ ),
    .Y(\hash/CA1/_0601_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2963_  (.A(\hash/CA1/_1947_ ),
    .B(\hash/CA1/_1950_ ),
    .Y(\hash/CA1/_0602_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_2964_  (.A_N(\hash/CA1/_1944_ ),
    .B(\hash/CA1/_0591_ ),
    .Y(\hash/CA1/_0603_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2965_  (.A1(\hash/CA1/_1947_ ),
    .A2(\hash/CA1/_0603_ ),
    .B1(\hash/CA1/_1946_ ),
    .X(\hash/CA1/_0604_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2966_  (.A1(\hash/CA1/_1950_ ),
    .A2(\hash/CA1/_0604_ ),
    .B1(\hash/CA1/_1949_ ),
    .Y(\hash/CA1/_0605_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2967_  (.A1(\hash/CA1/_0588_ ),
    .A2(\hash/CA1/_0596_ ),
    .A3(\hash/CA1/_0602_ ),
    .B1(\hash/CA1/_0605_ ),
    .Y(\hash/CA1/_0606_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2968_  (.A(\hash/CA1/_0601_ ),
    .B(\hash/CA1/_0606_ ),
    .Y(\hash/p2[24] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2969_  (.A(\hash/CA1/_1949_ ),
    .Y(\hash/CA1/_0607_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_2970_  (.A1(\hash/CA1/_1947_ ),
    .A2(\hash/CA1/_1946_ ),
    .B1(\hash/CA1/_1950_ ),
    .X(\hash/CA1/_0608_ ));
 sky130_fd_sc_hd__o41ai_2 \hash/CA1/_2971_  (.A1(\hash/CA1/_1944_ ),
    .A2(\hash/CA1/_1946_ ),
    .A3(\hash/CA1/_0590_ ),
    .A4(\hash/CA1/_0593_ ),
    .B1(\hash/CA1/_0608_ ),
    .Y(\hash/CA1/_0609_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2972_  (.A1(\hash/CA1/_0607_ ),
    .A2(\hash/CA1/_0609_ ),
    .B1(\hash/CA1/_0601_ ),
    .Y(\hash/CA1/_0610_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2973_  (.A(\hash/CA1/_1952_ ),
    .B(\hash/CA1/_0610_ ),
    .Y(\hash/CA1/_0611_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_2974_  (.A(\hash/CA1/_1956_ ),
    .B(\hash/CA1/_0611_ ),
    .Y(\hash/p2[25] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2976_  (.A(\hash/CA1/_1950_ ),
    .B(\hash/CA1/_1946_ ),
    .Y(\hash/CA1/_0613_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2977_  (.A(\hash/CA1/_1953_ ),
    .B(\hash/CA1/_1956_ ),
    .Y(\hash/CA1/_0614_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_2978_  (.A1(\hash/CA1/_1953_ ),
    .A2(\hash/CA1/_1949_ ),
    .B1(\hash/CA1/_1952_ ),
    .X(\hash/CA1/_0615_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2979_  (.A1(\hash/CA1/_1956_ ),
    .A2(\hash/CA1/_0615_ ),
    .B1(\hash/CA1/_1955_ ),
    .Y(\hash/CA1/_0616_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2980_  (.A1(\hash/CA1/_0613_ ),
    .A2(\hash/CA1/_0614_ ),
    .B1(\hash/CA1/_0616_ ),
    .Y(\hash/CA1/_0617_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2981_  (.A(\hash/CA1/_1959_ ),
    .B(\hash/CA1/_0603_ ),
    .C(\hash/CA1/_0617_ ),
    .Y(\hash/CA1/_0618_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_2982_  (.A(\hash/CA1/_1959_ ),
    .Y(\hash/CA1/_0619_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2983_  (.A(\hash/CA1/_0619_ ),
    .B(\hash/CA1/_0596_ ),
    .C(\hash/CA1/_0597_ ),
    .Y(\hash/CA1/_0620_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2984_  (.A(\hash/CA1/_0602_ ),
    .B(\hash/CA1/_0614_ ),
    .Y(\hash/CA1/_0621_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2985_  (.A(\hash/CA1/_1959_ ),
    .B(\hash/CA1/_0603_ ),
    .C(\hash/CA1/_0621_ ),
    .Y(\hash/CA1/_0622_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_2986_  (.A(\hash/CA1/_1959_ ),
    .B(\hash/CA1/_0617_ ),
    .C(\hash/CA1/_0621_ ),
    .Y(\hash/CA1/_0623_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2987_  (.A1(\hash/CA1/_1959_ ),
    .A2(\hash/CA1/_0617_ ),
    .B1(\hash/CA1/_0623_ ),
    .Y(\hash/CA1/_0624_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_2988_  (.A1(\hash/CA1/_0617_ ),
    .A2(\hash/CA1/_0620_ ),
    .B1(\hash/CA1/_0622_ ),
    .C1(\hash/CA1/_0624_ ),
    .Y(\hash/CA1/_0625_ ));
 sky130_fd_sc_hd__nor4b_1 \hash/CA1/_2989_  (.A(\hash/CA1/_0619_ ),
    .B(\hash/CA1/_0588_ ),
    .C(\hash/CA1/_0596_ ),
    .D_N(\hash/CA1/_0621_ ),
    .Y(\hash/CA1/_0626_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_2990_  (.A1(\hash/CA1/_0588_ ),
    .A2(\hash/CA1/_0618_ ),
    .B1(\hash/CA1/_0625_ ),
    .C1(\hash/CA1/_0626_ ),
    .Y(\hash/p2[26] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_2991_  (.A(\hash/CA1/_1959_ ),
    .B(\hash/CA1/_1961_ ),
    .Y(\hash/CA1/_0627_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2992_  (.A(\hash/CA1/_0616_ ),
    .B(\hash/CA1/_0627_ ),
    .Y(\hash/CA1/_0628_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2993_  (.A1(\hash/CA1/_1961_ ),
    .A2(\hash/CA1/_1958_ ),
    .B1(\hash/CA1/_0628_ ),
    .Y(\hash/CA1/_0629_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_2994_  (.A1(\hash/CA1/_0609_ ),
    .A2(\hash/CA1/_0614_ ),
    .A3(\hash/CA1/_0627_ ),
    .B1(\hash/CA1/_0629_ ),
    .Y(\hash/CA1/_0630_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_2995_  (.A1(\hash/CA1/_0599_ ),
    .A2(\hash/CA1/_0621_ ),
    .B1(\hash/CA1/_0617_ ),
    .Y(\hash/CA1/_0631_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_2996_  (.A(\hash/CA1/_1961_ ),
    .B(\hash/CA1/_1958_ ),
    .Y(\hash/CA1/_0632_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_2997_  (.A1(\hash/CA1/_0619_ ),
    .A2(\hash/CA1/_0631_ ),
    .B1(\hash/CA1/_0632_ ),
    .Y(\hash/CA1/_0633_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_2998_  (.A(\hash/CA1/_0630_ ),
    .B_N(\hash/CA1/_0633_ ),
    .Y(\hash/p2[27] ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_2999_  (.A(\hash/CA1/_1959_ ),
    .B(\hash/CA1/_1961_ ),
    .C(\hash/CA1/_0621_ ),
    .Y(\hash/CA1/_0634_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3000_  (.A1(\hash/CA1/_0601_ ),
    .A2(\hash/CA1/_0605_ ),
    .B1_N(\hash/CA1/_1952_ ),
    .Y(\hash/CA1/_0635_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3001_  (.A1(\hash/CA1/_1956_ ),
    .A2(\hash/CA1/_0635_ ),
    .B1(\hash/CA1/_1955_ ),
    .Y(\hash/CA1/_0636_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3002_  (.A1(\hash/CA1/_0619_ ),
    .A2(\hash/CA1/_0636_ ),
    .B1_N(\hash/CA1/_1958_ ),
    .Y(\hash/CA1/_0637_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3003_  (.A1(\hash/CA1/_1961_ ),
    .A2(\hash/CA1/_0637_ ),
    .B1(\hash/CA1/_1960_ ),
    .Y(\hash/CA1/_0638_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_3004_  (.A1(\hash/CA1/_0588_ ),
    .A2(\hash/CA1/_0596_ ),
    .A3(\hash/CA1/_0634_ ),
    .B1(\hash/CA1/_0638_ ),
    .Y(\hash/CA1/_0639_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3005_  (.A(\hash/CA1/_1963_ ),
    .B(\hash/CA1/_0639_ ),
    .X(\hash/p2[28] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3006_  (.A1(\hash/CA1/_1960_ ),
    .A2(\hash/CA1/_0630_ ),
    .B1(\hash/CA1/_1963_ ),
    .X(\hash/CA1/_0640_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3007_  (.A(\hash/CA1/_1962_ ),
    .B(\hash/CA1/_0640_ ),
    .Y(\hash/CA1/_0641_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3008_  (.A(\hash/CA1/_1966_ ),
    .B(\hash/CA1/_0641_ ),
    .Y(\hash/p2[29] ));
 sky130_fd_sc_hd__nor3b_1 \hash/CA1/_3009_  (.A(\hash/CA1/_0589_ ),
    .B(\hash/CA1/_0634_ ),
    .C_N(\hash/CA1/_0587_ ),
    .Y(\hash/CA1/_0642_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3010_  (.A1(\hash/CA1/_0592_ ),
    .A2(\hash/CA1/_0597_ ),
    .B1(\hash/CA1/_0634_ ),
    .Y(\hash/CA1/_0643_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3011_  (.A1(\hash/CA1/_1963_ ),
    .A2(\hash/CA1/_1962_ ),
    .B1(\hash/CA1/_1966_ ),
    .Y(\hash/CA1/_0644_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3012_  (.A(\hash/CA1/_1969_ ),
    .B(\hash/CA1/_0644_ ),
    .Y(\hash/CA1/_0645_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3013_  (.A1(\hash/CA1/_0642_ ),
    .A2(\hash/CA1/_0643_ ),
    .B1(\hash/CA1/_0645_ ),
    .Y(\hash/CA1/_0646_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3014_  (.A1(\hash/CA1/_1959_ ),
    .A2(\hash/CA1/_0617_ ),
    .B1(\hash/CA1/_1958_ ),
    .X(\hash/CA1/_0647_ ));
 sky130_fd_sc_hd__a211o_1 \hash/CA1/_3015_  (.A1(\hash/CA1/_1961_ ),
    .A2(\hash/CA1/_0647_ ),
    .B1(\hash/CA1/_1962_ ),
    .C1(\hash/CA1/_1960_ ),
    .X(\hash/CA1/_0648_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3016_  (.A(\hash/CA1/_1965_ ),
    .Y(\hash/CA1/_0649_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3017_  (.A(\hash/CA1/_1969_ ),
    .B(\hash/CA1/_0649_ ),
    .Y(\hash/CA1/_0650_ ));
 sky130_fd_sc_hd__or4_1 \hash/CA1/_3018_  (.A(\hash/CA1/_0648_ ),
    .B(\hash/CA1/_0642_ ),
    .C(\hash/CA1/_0643_ ),
    .D(\hash/CA1/_0650_ ),
    .X(\hash/CA1/_0651_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3019_  (.A(\hash/CA1/_1969_ ),
    .Y(\hash/CA1/_0652_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_3020_  (.A(\hash/CA1/_1969_ ),
    .B(\hash/CA1/_0649_ ),
    .C(\hash/CA1/_0644_ ),
    .X(\hash/CA1/_0653_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA1/_3021_  (.A1(\hash/CA1/_0652_ ),
    .A2(\hash/CA1/_1965_ ),
    .B1(\hash/CA1/_0648_ ),
    .B2(\hash/CA1/_0645_ ),
    .C1(\hash/CA1/_0653_ ),
    .Y(\hash/CA1/_0654_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3022_  (.A(\hash/CA1/_0646_ ),
    .B(\hash/CA1/_0651_ ),
    .C(\hash/CA1/_0654_ ),
    .Y(\hash/p2[30] ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3023_  (.A(\hash/h[31] ),
    .B(\hash/CA1/s1[31] ),
    .X(\hash/CA1/_0655_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3024_  (.A(\k_value1[31] ),
    .B(\w_value1[31] ),
    .Y(\hash/CA1/_0656_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3025_  (.A(\hash/CA1/_0655_ ),
    .B(\hash/CA1/_0656_ ),
    .Y(\hash/CA1/_0657_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA1/_3026_  (.A0(\hash/g[31] ),
    .A1(\hash/f[31] ),
    .S(\hash/e[31] ),
    .Y(\hash/CA1/_0658_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3027_  (.A(\hash/CA1/_0657_ ),
    .B(\hash/CA1/_0658_ ),
    .Y(\hash/CA1/_0659_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3028_  (.A1(\hash/CA1/_1877_ ),
    .A2(\hash/CA1/_0253_ ),
    .B1(\hash/CA1/_1876_ ),
    .Y(\hash/CA1/_0660_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3029_  (.A(\hash/CA1/_0206_ ),
    .B(\hash/CA1/_0257_ ),
    .C(\hash/CA1/_0660_ ),
    .Y(\hash/CA1/_0661_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3030_  (.A(\hash/CA1/_1862_ ),
    .B(\hash/CA1/_1870_ ),
    .C(\hash/CA1/_1877_ ),
    .Y(\hash/CA1/_0662_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3031_  (.A1(\hash/CA1/_1844_ ),
    .A2(\hash/CA1/_1853_ ),
    .B1(\hash/CA1/_0248_ ),
    .Y(\hash/CA1/_0663_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3032_  (.A1(\hash/CA1/_0662_ ),
    .A2(\hash/CA1/_0663_ ),
    .B1(\hash/CA1/_0660_ ),
    .Y(\hash/CA1/_0664_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_3033_  (.A1(\hash/CA1/_1884_ ),
    .A2(\hash/CA1/_0661_ ),
    .A3(\hash/CA1/_0664_ ),
    .B1(\hash/CA1/_1883_ ),
    .Y(\hash/CA1/_0665_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3034_  (.A(\hash/CA1/_0659_ ),
    .B(\hash/CA1/_0665_ ),
    .Y(\hash/CA1/_0666_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3035_  (.A1(\hash/CA1/_1874_ ),
    .A2(\hash/CA1/_0245_ ),
    .B1(\hash/CA1/_1873_ ),
    .X(\hash/CA1/_0667_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3036_  (.A1(\hash/CA1/_1881_ ),
    .A2(\hash/CA1/_0667_ ),
    .B1(\hash/CA1/_1880_ ),
    .Y(\hash/CA1/_0668_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3037_  (.A(\hash/CA1/_0666_ ),
    .B(\hash/CA1/_0668_ ),
    .Y(\hash/CA1/_0669_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3038_  (.A1(\hash/CA1/_0649_ ),
    .A2(\hash/CA1/_0644_ ),
    .B1(\hash/CA1/_0652_ ),
    .Y(\hash/CA1/_0670_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3039_  (.A(\hash/CA1/_1960_ ),
    .B(\hash/CA1/_1962_ ),
    .C(\hash/CA1/_1968_ ),
    .Y(\hash/CA1/_0671_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3040_  (.A1(\hash/CA1/_0652_ ),
    .A2(\hash/CA1/_0649_ ),
    .B1(\hash/CA1/_0671_ ),
    .Y(\hash/CA1/_0672_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA1/_3041_  (.A1(\hash/CA1/_1968_ ),
    .A2(\hash/CA1/_0670_ ),
    .B1(\hash/CA1/_0672_ ),
    .B2(\hash/CA1/_0630_ ),
    .Y(\hash/CA1/_0673_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3042_  (.A(\hash/CA1/_1408_ ),
    .B(\hash/CA1/_1411_ ),
    .X(\hash/CA1/_0674_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3043_  (.A(\hash/d[31] ),
    .B(\hash/CA1/_0674_ ),
    .Y(\hash/CA1/_0675_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3044_  (.A(\hash/CA1/_0673_ ),
    .B(\hash/CA1/_0675_ ),
    .Y(\hash/CA1/_0676_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3045_  (.A(\hash/CA1/_0669_ ),
    .B(\hash/CA1/_0676_ ),
    .Y(\hash/p2[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3046_  (.A(\hash/CA1/_1418_ ),
    .B(\hash/CA1/_1891_ ),
    .Y(\hash/p2[3] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3047_  (.A(\hash/CA1/_1893_ ),
    .B(\hash/CA1/_0531_ ),
    .Y(\hash/p2[4] ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3048_  (.A(\hash/CA1/_1892_ ),
    .B_N(\hash/CA1/_0540_ ),
    .Y(\hash/CA1/_0677_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3049_  (.A(\hash/CA1/_1896_ ),
    .B(\hash/CA1/_0677_ ),
    .Y(\hash/p2[5] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3050_  (.A(\hash/CA1/_1900_ ),
    .B(\hash/CA1/_0533_ ),
    .Y(\hash/p2[6] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3051_  (.A1(\hash/CA1/_0540_ ),
    .A2(\hash/CA1/_0541_ ),
    .B1(\hash/CA1/_0543_ ),
    .Y(\hash/CA1/_0678_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3052_  (.A(\hash/CA1/_1899_ ),
    .B(\hash/CA1/_0678_ ),
    .Y(\hash/CA1/_0679_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3053_  (.A(\hash/CA1/_1904_ ),
    .B(\hash/CA1/_0679_ ),
    .Y(\hash/p2[7] ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3054_  (.A1(\hash/CA1/_0528_ ),
    .A2(\hash/CA1/_0533_ ),
    .B1_N(\hash/CA1/_1899_ ),
    .Y(\hash/CA1/_0680_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3055_  (.A1(\hash/CA1/_1904_ ),
    .A2(\hash/CA1/_0680_ ),
    .B1(\hash/CA1/_1903_ ),
    .Y(\hash/CA1/_0681_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3056_  (.A(\hash/CA1/_1907_ ),
    .B(\hash/CA1/_0681_ ),
    .Y(\hash/p2[8] ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3057_  (.A_N(\hash/CA1/_0678_ ),
    .B(\hash/CA1/_0534_ ),
    .Y(\hash/CA1/_0682_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3058_  (.A1(\hash/CA1/_1906_ ),
    .A2(\hash/CA1/_0526_ ),
    .B1(\hash/CA1/_0682_ ),
    .Y(\hash/CA1/_0683_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3059_  (.A(\hash/CA1/_1910_ ),
    .B(\hash/CA1/_0683_ ),
    .Y(\hash/p2[9] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3060_  (.A(\hash/CA1/_1669_ ),
    .Y(\hash/CA1/_0684_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3061_  (.A1(\hash/CA1/_1976_ ),
    .A2(\hash/CA1/_1654_ ),
    .B1(\hash/CA1/_1653_ ),
    .X(\hash/CA1/_0685_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3062_  (.A1(\hash/CA1/_1661_ ),
    .A2(\hash/CA1/_0685_ ),
    .B1(\hash/CA1/_1660_ ),
    .Y(\hash/CA1/_0686_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3063_  (.A(\hash/CA1/_1668_ ),
    .B(\hash/CA1/_1676_ ),
    .Y(\hash/CA1/_0687_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3064_  (.A1(\hash/CA1/_0684_ ),
    .A2(\hash/CA1/_0686_ ),
    .B1(\hash/CA1/_0687_ ),
    .Y(\hash/CA1/_0688_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3065_  (.A1(\hash/CA1/_1677_ ),
    .A2(\hash/CA1/_1676_ ),
    .B1(\hash/CA1/_1684_ ),
    .X(\hash/CA1/_0689_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3066_  (.A1(\hash/CA1/_0688_ ),
    .A2(\hash/CA1/_0689_ ),
    .B1(\hash/CA1/_1683_ ),
    .X(\hash/CA1/_0690_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3067_  (.A1(\hash/CA1/_1691_ ),
    .A2(\hash/CA1/_0690_ ),
    .B1(\hash/CA1/_1690_ ),
    .Y(\hash/CA1/_0691_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3068_  (.A(\hash/CA1/_0691_ ),
    .B_N(\hash/CA1/_1698_ ),
    .Y(\hash/CA1/_0692_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3070_  (.A1(\hash/CA1/_1697_ ),
    .A2(\hash/CA1/_0692_ ),
    .B1(\hash/CA1/_1706_ ),
    .X(\hash/CA1/_0694_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3071_  (.A(\hash/CA1/_1705_ ),
    .B(\hash/CA1/_0694_ ),
    .Y(\hash/CA1/_0695_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3072_  (.A(\hash/CA1/_1715_ ),
    .B(\hash/CA1/_0695_ ),
    .Y(\hash/p3[10] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3073_  (.A1(\hash/CA1/_1684_ ),
    .A2(\hash/CA1/_1683_ ),
    .B1(\hash/CA1/_1691_ ),
    .X(\hash/CA1/_0696_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3074_  (.A1(\hash/CA1/_1690_ ),
    .A2(\hash/CA1/_0696_ ),
    .B1(\hash/CA1/_1698_ ),
    .Y(\hash/CA1/_0697_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_3075_  (.A(\hash/CA1/_1683_ ),
    .B(\hash/CA1/_1690_ ),
    .X(\hash/CA1/_0698_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3076_  (.A(\hash/CA1/_1668_ ),
    .Y(\hash/CA1/_0699_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3077_  (.A(\hash/CA1/_1426_ ),
    .B_N(\hash/CA1/_1661_ ),
    .Y(\hash/CA1/_0700_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3078_  (.A1(\hash/CA1/_1660_ ),
    .A2(\hash/CA1/_0700_ ),
    .B1(\hash/CA1/_1669_ ),
    .Y(\hash/CA1/_0701_ ));
 sky130_fd_sc_hd__a21boi_1 \hash/CA1/_3079_  (.A1(\hash/CA1/_0699_ ),
    .A2(\hash/CA1/_0701_ ),
    .B1_N(\hash/CA1/_1677_ ),
    .Y(\hash/CA1/_0702_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3080_  (.A(\hash/CA1/_1676_ ),
    .B(\hash/CA1/_0698_ ),
    .C(\hash/CA1/_0702_ ),
    .Y(\hash/CA1/_0703_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3081_  (.A(\hash/CA1/_0697_ ),
    .B(\hash/CA1/_0703_ ),
    .Y(\hash/CA1/_0704_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3082_  (.A1(\hash/CA1/_1697_ ),
    .A2(\hash/CA1/_0704_ ),
    .B1(\hash/CA1/_1706_ ),
    .Y(\hash/CA1/_0705_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3083_  (.A_N(\hash/CA1/_1705_ ),
    .B(\hash/CA1/_0705_ ),
    .Y(\hash/CA1/_0706_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3084_  (.A1(\hash/CA1/_1715_ ),
    .A2(\hash/CA1/_0706_ ),
    .B1(\hash/CA1/_1714_ ),
    .Y(\hash/CA1/_0707_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3085_  (.A(\hash/CA1/_1724_ ),
    .B(\hash/CA1/_0707_ ),
    .Y(\hash/p3[11] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3086_  (.A1(\hash/CA1/_1698_ ),
    .A2(\hash/CA1/_1697_ ),
    .B1(\hash/CA1/_1706_ ),
    .X(\hash/CA1/_0708_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3087_  (.A1(\hash/CA1/_1705_ ),
    .A2(\hash/CA1/_0708_ ),
    .B1(\hash/CA1/_1715_ ),
    .X(\hash/CA1/_0709_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3088_  (.A1(\hash/CA1/_1714_ ),
    .A2(\hash/CA1/_0709_ ),
    .B1(\hash/CA1/_1724_ ),
    .Y(\hash/CA1/_0710_ ));
 sky130_fd_sc_hd__a211o_1 \hash/CA1/_3089_  (.A1(\hash/CA1/_1706_ ),
    .A2(\hash/CA1/_1697_ ),
    .B1(\hash/CA1/_1705_ ),
    .C1(\hash/CA1/_1714_ ),
    .X(\hash/CA1/_0711_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_3090_  (.A1(\hash/CA1/_1691_ ),
    .A2(\hash/CA1/_0690_ ),
    .B1(\hash/CA1/_0711_ ),
    .C1(\hash/CA1/_1690_ ),
    .Y(\hash/CA1/_0712_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3091_  (.A1(\hash/CA1/_0710_ ),
    .A2(\hash/CA1/_0712_ ),
    .B1_N(\hash/CA1/_1723_ ),
    .Y(\hash/CA1/_0713_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3092_  (.A(\hash/CA1/_1733_ ),
    .B(\hash/CA1/_0713_ ),
    .X(\hash/p3[12] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3093_  (.A1(\hash/CA1/_1715_ ),
    .A2(\hash/CA1/_1705_ ),
    .B1(\hash/CA1/_1714_ ),
    .X(\hash/CA1/_0714_ ));
 sky130_fd_sc_hd__a41o_1 \hash/CA1/_3094_  (.A1(\hash/CA1/_1706_ ),
    .A2(\hash/CA1/_1715_ ),
    .A3(\hash/CA1/_1724_ ),
    .A4(\hash/CA1/_1697_ ),
    .B1(\hash/CA1/_1723_ ),
    .X(\hash/CA1/_0715_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3095_  (.A1(\hash/CA1/_1724_ ),
    .A2(\hash/CA1/_0714_ ),
    .B1(\hash/CA1/_0715_ ),
    .Y(\hash/CA1/_0716_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3096_  (.A(\hash/CA1/_1706_ ),
    .B(\hash/CA1/_1715_ ),
    .C(\hash/CA1/_1724_ ),
    .Y(\hash/CA1/_0717_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3097_  (.A(\hash/CA1/_0697_ ),
    .B(\hash/CA1/_0717_ ),
    .Y(\hash/CA1/_0718_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_3098_  (.A1(\hash/CA1/_1676_ ),
    .A2(\hash/CA1/_0698_ ),
    .A3(\hash/CA1/_0702_ ),
    .B1(\hash/CA1/_0718_ ),
    .Y(\hash/CA1/_0719_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3099_  (.A(\hash/CA1/_0716_ ),
    .B(\hash/CA1/_0719_ ),
    .Y(\hash/CA1/_0720_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3100_  (.A1(\hash/CA1/_1733_ ),
    .A2(\hash/CA1/_0720_ ),
    .B1(\hash/CA1/_1732_ ),
    .Y(\hash/CA1/_0721_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3101_  (.A(\hash/CA1/_1742_ ),
    .B(\hash/CA1/_0721_ ),
    .Y(\hash/p3[13] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3102_  (.A(\hash/CA1/_1751_ ),
    .Y(\hash/CA1/_0722_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3103_  (.A(\hash/CA1/_1742_ ),
    .B(\hash/CA1/_1741_ ),
    .Y(\hash/CA1/_0723_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3104_  (.A(\hash/CA1/_1732_ ),
    .B(\hash/CA1/_1741_ ),
    .Y(\hash/CA1/_0724_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA1/_3105_  (.A1(\hash/CA1/_1733_ ),
    .A2(\hash/CA1/_0713_ ),
    .B1_N(\hash/CA1/_0724_ ),
    .Y(\hash/CA1/_0725_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3106_  (.A(\hash/CA1/_0723_ ),
    .B(\hash/CA1/_0725_ ),
    .Y(\hash/CA1/_0726_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3107_  (.A(\hash/CA1/_0722_ ),
    .B(\hash/CA1/_0726_ ),
    .Y(\hash/p3[14] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3108_  (.A1(\hash/CA1/_1733_ ),
    .A2(\hash/CA1/_1732_ ),
    .B1(\hash/CA1/_1742_ ),
    .X(\hash/CA1/_0727_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3109_  (.A1(\hash/CA1/_1741_ ),
    .A2(\hash/CA1/_0727_ ),
    .B1(\hash/CA1/_1751_ ),
    .Y(\hash/CA1/_0728_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3110_  (.A(\hash/CA1/_1732_ ),
    .B(\hash/CA1/_1741_ ),
    .C(\hash/CA1/_0720_ ),
    .Y(\hash/CA1/_0729_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3111_  (.A(\hash/CA1/_1750_ ),
    .Y(\hash/CA1/_0730_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3112_  (.A1(\hash/CA1/_0728_ ),
    .A2(\hash/CA1/_0729_ ),
    .B1(\hash/CA1/_0730_ ),
    .Y(\hash/CA1/_0731_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3113_  (.A(\hash/CA1/_1759_ ),
    .B(\hash/CA1/_0731_ ),
    .X(\hash/p3[15] ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_3114_  (.A1(\hash/CA1/_0722_ ),
    .A2(\hash/CA1/_0723_ ),
    .A3(\hash/CA1/_0725_ ),
    .B1(\hash/CA1/_0730_ ),
    .Y(\hash/CA1/_0732_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3115_  (.A1(\hash/CA1/_1759_ ),
    .A2(\hash/CA1/_0732_ ),
    .B1(\hash/CA1/_1758_ ),
    .Y(\hash/CA1/_0733_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3116_  (.A(\hash/CA1/_1767_ ),
    .B(\hash/CA1/_0733_ ),
    .Y(\hash/p3[16] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3117_  (.A1(\hash/CA1/_1767_ ),
    .A2(\hash/CA1/_1758_ ),
    .B1(\hash/CA1/_1766_ ),
    .X(\hash/CA1/_0734_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3118_  (.A1(\hash/CA1/_1776_ ),
    .A2(\hash/CA1/_0734_ ),
    .B1(\hash/CA1/_1750_ ),
    .Y(\hash/CA1/_0735_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_3119_  (.A(\hash/CA1/_0716_ ),
    .B(\hash/CA1/_0724_ ),
    .C(\hash/CA1/_0735_ ),
    .X(\hash/CA1/_0736_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3120_  (.A1(\hash/CA1/_1759_ ),
    .A2(\hash/CA1/_1758_ ),
    .B1(\hash/CA1/_1767_ ),
    .X(\hash/CA1/_0737_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3121_  (.A(\hash/CA1/_0728_ ),
    .B(\hash/CA1/_0735_ ),
    .Y(\hash/CA1/_0738_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_3122_  (.A1(\hash/CA1/_1766_ ),
    .A2(\hash/CA1/_0737_ ),
    .B1(\hash/CA1/_0738_ ),
    .C1(\hash/CA1/_1776_ ),
    .Y(\hash/CA1/_0739_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3123_  (.A1(\hash/CA1/_0719_ ),
    .A2(\hash/CA1/_0736_ ),
    .B1(\hash/CA1/_0739_ ),
    .Y(\hash/CA1/_0740_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3124_  (.A1(\hash/CA1/_1759_ ),
    .A2(\hash/CA1/_0731_ ),
    .B1(\hash/CA1/_1758_ ),
    .X(\hash/CA1/_0741_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_3125_  (.A1(\hash/CA1/_1767_ ),
    .A2(\hash/CA1/_0741_ ),
    .B1(\hash/CA1/_1766_ ),
    .C1(\hash/CA1/_1776_ ),
    .Y(\hash/CA1/_0742_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3126_  (.A(\hash/CA1/_0740_ ),
    .B(\hash/CA1/_0742_ ),
    .Y(\hash/p3[17] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3127_  (.A1(\hash/CA1/_1733_ ),
    .A2(\hash/CA1/_1723_ ),
    .B1(\hash/CA1/_1732_ ),
    .X(\hash/CA1/_0743_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3128_  (.A1(\hash/CA1/_1742_ ),
    .A2(\hash/CA1/_0743_ ),
    .B1(\hash/CA1/_1741_ ),
    .Y(\hash/CA1/_0744_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3129_  (.A1(\hash/CA1/_0722_ ),
    .A2(\hash/CA1/_0744_ ),
    .B1(\hash/CA1/_0730_ ),
    .Y(\hash/CA1/_0745_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3130_  (.A1(\hash/CA1/_1759_ ),
    .A2(\hash/CA1/_0745_ ),
    .B1(\hash/CA1/_1758_ ),
    .X(\hash/CA1/_0746_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3131_  (.A1(\hash/CA1/_1767_ ),
    .A2(\hash/CA1/_0746_ ),
    .B1(\hash/CA1/_1766_ ),
    .Y(\hash/CA1/_0747_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3132_  (.A(\hash/CA1/_1733_ ),
    .B(\hash/CA1/_1742_ ),
    .Y(\hash/CA1/_0748_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3133_  (.A(\hash/CA1/_1751_ ),
    .B(\hash/CA1/_1759_ ),
    .C(\hash/CA1/_1767_ ),
    .Y(\hash/CA1/_0749_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3134_  (.A(\hash/CA1/_1691_ ),
    .B(\hash/CA1/_1690_ ),
    .C(\hash/CA1/_0711_ ),
    .Y(\hash/CA1/_0750_ ));
 sky130_fd_sc_hd__nor4_1 \hash/CA1/_3135_  (.A(\hash/CA1/_0710_ ),
    .B(\hash/CA1/_0748_ ),
    .C(\hash/CA1/_0749_ ),
    .D(\hash/CA1/_0750_ ),
    .Y(\hash/CA1/_0751_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA1/_3136_  (.A1(\hash/CA1/_1690_ ),
    .A2(\hash/CA1/_0690_ ),
    .A3(\hash/CA1/_0711_ ),
    .B1(\hash/CA1/_0751_ ),
    .Y(\hash/CA1/_0752_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3137_  (.A(\hash/CA1/_0747_ ),
    .B(\hash/CA1/_0752_ ),
    .Y(\hash/CA1/_0753_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3138_  (.A1(\hash/CA1/_1776_ ),
    .A2(\hash/CA1/_0753_ ),
    .B1(\hash/CA1/_1775_ ),
    .Y(\hash/CA1/_0754_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3139_  (.A(\hash/CA1/_1785_ ),
    .B(\hash/CA1/_0754_ ),
    .Y(\hash/p3[18] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3140_  (.A1(\hash/CA1/_1785_ ),
    .A2(\hash/CA1/_1784_ ),
    .B1(\hash/CA1/_1794_ ),
    .X(\hash/CA1/_0755_ ));
 sky130_fd_sc_hd__o31a_1 \hash/CA1/_3141_  (.A1(\hash/CA1/_1775_ ),
    .A2(\hash/CA1/_1784_ ),
    .A3(\hash/CA1/_0740_ ),
    .B1(\hash/CA1/_0755_ ),
    .X(\hash/CA1/_0756_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3142_  (.A1(\hash/CA1/_1775_ ),
    .A2(\hash/CA1/_0740_ ),
    .B1(\hash/CA1/_1785_ ),
    .X(\hash/CA1/_0757_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3143_  (.A(\hash/CA1/_1794_ ),
    .B(\hash/CA1/_1784_ ),
    .C(\hash/CA1/_0757_ ),
    .Y(\hash/CA1/_0758_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3144_  (.A(\hash/CA1/_0756_ ),
    .B(\hash/CA1/_0758_ ),
    .Y(\hash/p3[19] ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3145_  (.A(\hash/CA1/_1775_ ),
    .B(\hash/CA1/_1784_ ),
    .C(\hash/CA1/_1793_ ),
    .Y(\hash/CA1/_0759_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3146_  (.A1(\hash/CA1/_1776_ ),
    .A2(\hash/CA1/_1775_ ),
    .B1(\hash/CA1/_1785_ ),
    .X(\hash/CA1/_0760_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3147_  (.A1(\hash/CA1/_1784_ ),
    .A2(\hash/CA1/_0760_ ),
    .B1(\hash/CA1/_1794_ ),
    .Y(\hash/CA1/_0761_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3148_  (.A_N(\hash/CA1/_1793_ ),
    .B(\hash/CA1/_0761_ ),
    .Y(\hash/CA1/_0762_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3149_  (.A(\hash/CA1/_0762_ ),
    .Y(\hash/CA1/_0763_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_3150_  (.A1(\hash/CA1/_0747_ ),
    .A2(\hash/CA1/_0752_ ),
    .A3(\hash/CA1/_0759_ ),
    .B1(\hash/CA1/_0763_ ),
    .Y(\hash/CA1/_0764_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3151_  (.A(\hash/CA1/_1803_ ),
    .B(\hash/CA1/_0764_ ),
    .X(\hash/p3[20] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3152_  (.A1(\hash/CA1/_1793_ ),
    .A2(\hash/CA1/_0756_ ),
    .B1(\hash/CA1/_1803_ ),
    .X(\hash/CA1/_0765_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3153_  (.A(\hash/CA1/_1802_ ),
    .B(\hash/CA1/_0765_ ),
    .Y(\hash/CA1/_0766_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3154_  (.A(\hash/CA1/_1812_ ),
    .B(\hash/CA1/_0766_ ),
    .Y(\hash/p3[21] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3155_  (.A1(\hash/CA1/_1803_ ),
    .A2(\hash/CA1/_0764_ ),
    .B1(\hash/CA1/_1802_ ),
    .X(\hash/CA1/_0767_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3156_  (.A1(\hash/CA1/_1812_ ),
    .A2(\hash/CA1/_0767_ ),
    .B1(\hash/CA1/_1811_ ),
    .Y(\hash/CA1/_0768_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3157_  (.A(\hash/CA1/_1821_ ),
    .B(\hash/CA1/_0768_ ),
    .Y(\hash/p3[22] ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3158_  (.A1(\hash/CA1/_1821_ ),
    .A2(\hash/CA1/_1811_ ),
    .B1(\hash/CA1/_1820_ ),
    .Y(\hash/CA1/_0769_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3159_  (.A(\hash/CA1/_1793_ ),
    .B(\hash/CA1/_1802_ ),
    .Y(\hash/CA1/_0770_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3160_  (.A(\hash/CA1/_0769_ ),
    .B(\hash/CA1/_0770_ ),
    .Y(\hash/CA1/_0771_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3161_  (.A(\hash/CA1/_1812_ ),
    .B(\hash/CA1/_1821_ ),
    .Y(\hash/CA1/_0772_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3162_  (.A(\hash/CA1/_1803_ ),
    .B(\hash/CA1/_1802_ ),
    .Y(\hash/CA1/_0773_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3163_  (.A1(\hash/CA1/_0772_ ),
    .A2(\hash/CA1/_0773_ ),
    .B1(\hash/CA1/_0769_ ),
    .Y(\hash/CA1/_0774_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_3164_  (.A1(\hash/CA1/_0756_ ),
    .A2(\hash/CA1/_0771_ ),
    .B1(\hash/CA1/_0774_ ),
    .Y(\hash/CA1/_0775_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3165_  (.A(\hash/CA1/_1830_ ),
    .B(\hash/CA1/_0775_ ),
    .Y(\hash/p3[23] ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_3166_  (.A(\hash/CA1/_1803_ ),
    .B(\hash/CA1/_1812_ ),
    .C(\hash/CA1/_1821_ ),
    .X(\hash/CA1/_0776_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3167_  (.A(\hash/CA1/_1821_ ),
    .B(\hash/CA1/_1811_ ),
    .Y(\hash/CA1/_0777_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3168_  (.A(\hash/CA1/_1812_ ),
    .B(\hash/CA1/_1821_ ),
    .C(\hash/CA1/_1802_ ),
    .Y(\hash/CA1/_0778_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3169_  (.A(\hash/CA1/_0777_ ),
    .B(\hash/CA1/_0778_ ),
    .Y(\hash/CA1/_0779_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3170_  (.A1(\hash/CA1/_0764_ ),
    .A2(\hash/CA1/_0776_ ),
    .B1(\hash/CA1/_0779_ ),
    .X(\hash/CA1/_0780_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3171_  (.A1(\hash/CA1/_1820_ ),
    .A2(\hash/CA1/_0780_ ),
    .B1(\hash/CA1/_1830_ ),
    .X(\hash/CA1/_0781_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3172_  (.A(\hash/CA1/_1829_ ),
    .B(\hash/CA1/_0781_ ),
    .Y(\hash/CA1/_0782_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3173_  (.A(\hash/CA1/_1839_ ),
    .B(\hash/CA1/_0782_ ),
    .Y(\hash/p3[24] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3174_  (.A(\hash/CA1/_1830_ ),
    .Y(\hash/CA1/_0783_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3175_  (.A1(\hash/CA1/_0783_ ),
    .A2(\hash/CA1/_0775_ ),
    .B1_N(\hash/CA1/_1829_ ),
    .Y(\hash/CA1/_0784_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3176_  (.A1(\hash/CA1/_1839_ ),
    .A2(\hash/CA1/_0784_ ),
    .B1(\hash/CA1/_1838_ ),
    .Y(\hash/CA1/_0785_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3177_  (.A(\hash/CA1/_1848_ ),
    .B(\hash/CA1/_0785_ ),
    .Y(\hash/p3[25] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3178_  (.A1(\hash/CA1/_1830_ ),
    .A2(\hash/CA1/_1820_ ),
    .B1(\hash/CA1/_1829_ ),
    .X(\hash/CA1/_0786_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3179_  (.A1(\hash/CA1/_1839_ ),
    .A2(\hash/CA1/_0786_ ),
    .B1(\hash/CA1/_1838_ ),
    .Y(\hash/CA1/_0787_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3180_  (.A(\hash/CA1/_0787_ ),
    .Y(\hash/CA1/_0788_ ));
 sky130_fd_sc_hd__a31o_2 \hash/CA1/_3181_  (.A1(\hash/CA1/_1830_ ),
    .A2(\hash/CA1/_1839_ ),
    .A3(\hash/CA1/_0780_ ),
    .B1(\hash/CA1/_0788_ ),
    .X(\hash/CA1/_0789_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3182_  (.A1(\hash/CA1/_1848_ ),
    .A2(\hash/CA1/_0789_ ),
    .B1(\hash/CA1/_1847_ ),
    .Y(\hash/CA1/_0790_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3183_  (.A(\hash/CA1/_1857_ ),
    .B(\hash/CA1/_0790_ ),
    .Y(\hash/p3[26] ));
 sky130_fd_sc_hd__and4_1 \hash/CA1/_3185_  (.A(\hash/CA1/_1830_ ),
    .B(\hash/CA1/_1839_ ),
    .C(\hash/CA1/_1848_ ),
    .D(\hash/CA1/_1857_ ),
    .X(\hash/CA1/_0792_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_3186_  (.A1(\hash/CA1/_0756_ ),
    .A2(\hash/CA1/_0771_ ),
    .B1(\hash/CA1/_0774_ ),
    .C1(\hash/CA1/_0792_ ),
    .Y(\hash/CA1/_0793_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3187_  (.A1(\hash/CA1/_1839_ ),
    .A2(\hash/CA1/_1829_ ),
    .B1(\hash/CA1/_1838_ ),
    .X(\hash/CA1/_0794_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3188_  (.A1(\hash/CA1/_1848_ ),
    .A2(\hash/CA1/_0794_ ),
    .B1(\hash/CA1/_1847_ ),
    .X(\hash/CA1/_0795_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3189_  (.A1(\hash/CA1/_1857_ ),
    .A2(\hash/CA1/_0795_ ),
    .B1(\hash/CA1/_1856_ ),
    .Y(\hash/CA1/_0796_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3190_  (.A(\hash/CA1/_0793_ ),
    .B(\hash/CA1/_0796_ ),
    .Y(\hash/CA1/_0797_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3191_  (.A(\hash/CA1/_1865_ ),
    .B(\hash/CA1/_0797_ ),
    .X(\hash/p3[27] ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3192_  (.A(\hash/CA1/_1872_ ),
    .B_N(\hash/CA1/_1865_ ),
    .Y(\hash/CA1/_0798_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3193_  (.A(\hash/CA1/_1872_ ),
    .Y(\hash/CA1/_0799_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3194_  (.A(\hash/CA1/_0799_ ),
    .B(\hash/CA1/_1856_ ),
    .C(\hash/CA1/_1864_ ),
    .Y(\hash/CA1/_0800_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA1/_3195_  (.A(\hash/CA1/_1848_ ),
    .B(\hash/CA1/_1857_ ),
    .C(\hash/CA1/_0788_ ),
    .X(\hash/CA1/_0801_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA1/_3196_  (.A1(\hash/CA1/_1857_ ),
    .A2(\hash/CA1/_1847_ ),
    .B1(\hash/CA1/_0780_ ),
    .B2(\hash/CA1/_0792_ ),
    .C1(\hash/CA1/_0801_ ),
    .Y(\hash/CA1/_0802_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA1/_3197_  (.A0(\hash/CA1/_0798_ ),
    .A1(\hash/CA1/_0800_ ),
    .S(\hash/CA1/_0802_ ),
    .Y(\hash/CA1/_0803_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3198_  (.A(\hash/CA1/_1865_ ),
    .B(\hash/CA1/_0799_ ),
    .C(\hash/CA1/_1864_ ),
    .Y(\hash/CA1/_0804_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA1/_3199_  (.A1(\hash/CA1/_0799_ ),
    .A2(\hash/CA1/_1864_ ),
    .B1(\hash/CA1/_0798_ ),
    .B2(\hash/CA1/_1856_ ),
    .C1(\hash/CA1/_0804_ ),
    .Y(\hash/CA1/_0805_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3200_  (.A(\hash/CA1/_0803_ ),
    .B(\hash/CA1/_0805_ ),
    .Y(\hash/p3[28] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3201_  (.A(\hash/CA1/_1879_ ),
    .Y(\hash/CA1/_0806_ ));
 sky130_fd_sc_hd__a2111o_1 \hash/CA1/_3202_  (.A1(\hash/CA1/_1865_ ),
    .A2(\hash/CA1/_0797_ ),
    .B1(\hash/CA1/_1871_ ),
    .C1(\hash/CA1/_1864_ ),
    .D1(\hash/CA1/_0806_ ),
    .X(\hash/CA1/_0807_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3203_  (.A(\hash/CA1/_0799_ ),
    .B(\hash/CA1/_1879_ ),
    .Y(\hash/CA1/_0808_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3204_  (.A(\hash/CA1/_1865_ ),
    .B(\hash/CA1/_0797_ ),
    .C(\hash/CA1/_0808_ ),
    .Y(\hash/CA1/_0809_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3205_  (.A(\hash/CA1/_1872_ ),
    .B(\hash/CA1/_0806_ ),
    .C(\hash/CA1/_1871_ ),
    .Y(\hash/CA1/_0810_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA1/_3206_  (.A1(\hash/CA1/_0806_ ),
    .A2(\hash/CA1/_1871_ ),
    .B1(\hash/CA1/_0808_ ),
    .B2(\hash/CA1/_1864_ ),
    .C1(\hash/CA1/_0810_ ),
    .Y(\hash/CA1/_0811_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3207_  (.A(\hash/CA1/_0807_ ),
    .B(\hash/CA1/_0809_ ),
    .C(\hash/CA1/_0811_ ),
    .Y(\hash/p3[29] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3208_  (.A(\hash/CA1/_1886_ ),
    .Y(\hash/CA1/_0812_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3209_  (.A(\hash/CA1/_1865_ ),
    .B(\hash/CA1/_1872_ ),
    .C(\hash/CA1/_1879_ ),
    .Y(\hash/CA1/_0813_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3210_  (.A1(\hash/CA1/_1865_ ),
    .A2(\hash/CA1/_1856_ ),
    .B1(\hash/CA1/_1864_ ),
    .Y(\hash/CA1/_0814_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3211_  (.A1(\hash/CA1/_0799_ ),
    .A2(\hash/CA1/_0814_ ),
    .B1_N(\hash/CA1/_1871_ ),
    .Y(\hash/CA1/_0815_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3212_  (.A1(\hash/CA1/_1879_ ),
    .A2(\hash/CA1/_0815_ ),
    .B1(\hash/CA1/_1878_ ),
    .Y(\hash/CA1/_0816_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3213_  (.A1(\hash/CA1/_0802_ ),
    .A2(\hash/CA1/_0813_ ),
    .B1(\hash/CA1/_0816_ ),
    .Y(\hash/CA1/_0817_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3214_  (.A(\hash/CA1/_0812_ ),
    .B(\hash/CA1/_0817_ ),
    .Y(\hash/p3[30] ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3215_  (.A1(\hash/CA1/_1872_ ),
    .A2(\hash/CA1/_1864_ ),
    .B1(\hash/CA1/_1871_ ),
    .Y(\hash/CA1/_0818_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3216_  (.A1(\hash/CA1/_0806_ ),
    .A2(\hash/CA1/_0818_ ),
    .B1_N(\hash/CA1/_1878_ ),
    .Y(\hash/CA1/_0819_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3217_  (.A1(\hash/CA1/_1886_ ),
    .A2(\hash/CA1/_0819_ ),
    .B1(\hash/CA1/_1885_ ),
    .Y(\hash/CA1/_0820_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3218_  (.A(\hash/CA1/_0796_ ),
    .B(\hash/CA1/_0820_ ),
    .Y(\hash/CA1/_0821_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3219_  (.A(\hash/CA1/_1211_ ),
    .B(\hash/CA1/_0821_ ),
    .Y(\hash/CA1/_0822_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3220_  (.A(\hash/CA1/_0812_ ),
    .B(\hash/CA1/_0813_ ),
    .Y(\hash/CA1/_0823_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3221_  (.A(\hash/CA1/_1211_ ),
    .B(\hash/CA1/_0792_ ),
    .C(\hash/CA1/_0823_ ),
    .Y(\hash/CA1/_0824_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3222_  (.A(\hash/CA1/_0775_ ),
    .B(\hash/CA1/_0824_ ),
    .Y(\hash/CA1/_0825_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3223_  (.A(\hash/CA1/_1211_ ),
    .B(\hash/CA1/_0823_ ),
    .Y(\hash/CA1/_0826_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA1/_3224_  (.A0(\hash/CA1/_1211_ ),
    .A1(\hash/CA1/_0826_ ),
    .S(\hash/CA1/_0820_ ),
    .Y(\hash/CA1/_0827_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA1/_3225_  (.A_N(\hash/CA1/_0796_ ),
    .B(\hash/CA1/_0823_ ),
    .C(\hash/CA1/_1211_ ),
    .Y(\hash/CA1/_0828_ ));
 sky130_fd_sc_hd__o311ai_0 \hash/CA1/_3226_  (.A1(\hash/CA1/_1211_ ),
    .A2(\hash/CA1/_0792_ ),
    .A3(\hash/CA1/_0821_ ),
    .B1(\hash/CA1/_0827_ ),
    .C1(\hash/CA1/_0828_ ),
    .Y(\hash/CA1/_0829_ ));
 sky130_fd_sc_hd__a211o_1 \hash/CA1/_3227_  (.A1(\hash/CA1/_0775_ ),
    .A2(\hash/CA1/_0822_ ),
    .B1(\hash/CA1/_0825_ ),
    .C1(\hash/CA1/_0829_ ),
    .X(\hash/CA1/_0830_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3228_  (.A(\hash/CA1/_0669_ ),
    .B(\hash/CA1/_0830_ ),
    .Y(\hash/p3[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3229_  (.A(\hash/CA1/_1426_ ),
    .B(\hash/CA1/_1661_ ),
    .Y(\hash/p3[3] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3230_  (.A(\hash/CA1/_1669_ ),
    .B(\hash/CA1/_0686_ ),
    .Y(\hash/p3[4] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3231_  (.A(\hash/CA1/_0699_ ),
    .B(\hash/CA1/_0701_ ),
    .Y(\hash/CA1/_0831_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3232_  (.A(\hash/CA1/_1677_ ),
    .B(\hash/CA1/_0831_ ),
    .Y(\hash/CA1/_0832_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3233_  (.A(\hash/CA1/_0702_ ),
    .B(\hash/CA1/_0832_ ),
    .Y(\hash/p3[5] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3234_  (.A1(\hash/CA1/_0684_ ),
    .A2(\hash/CA1/_0686_ ),
    .B1(\hash/CA1/_0699_ ),
    .Y(\hash/CA1/_0833_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3235_  (.A1(\hash/CA1/_1677_ ),
    .A2(\hash/CA1/_0833_ ),
    .B1(\hash/CA1/_1676_ ),
    .Y(\hash/CA1/_0834_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3236_  (.A(\hash/CA1/_1684_ ),
    .B(\hash/CA1/_0834_ ),
    .Y(\hash/p3[6] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3237_  (.A1(\hash/CA1/_1676_ ),
    .A2(\hash/CA1/_0702_ ),
    .B1(\hash/CA1/_1684_ ),
    .X(\hash/CA1/_0835_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3238_  (.A(\hash/CA1/_1683_ ),
    .B(\hash/CA1/_0835_ ),
    .Y(\hash/CA1/_0836_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3239_  (.A(\hash/CA1/_1691_ ),
    .B(\hash/CA1/_0836_ ),
    .Y(\hash/p3[7] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3240_  (.A(\hash/CA1/_1698_ ),
    .B(\hash/CA1/_0691_ ),
    .Y(\hash/p3[8] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3241_  (.A(\hash/CA1/_1697_ ),
    .B(\hash/CA1/_0704_ ),
    .Y(\hash/CA1/_0837_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3242_  (.A(\hash/CA1/_1706_ ),
    .B(\hash/CA1/_0837_ ),
    .Y(\hash/p3[9] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3243_  (.A(\w_value2[31] ),
    .B(\hash/CA1/_1052_ ),
    .Y(\hash/CA1/_0838_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3244_  (.A(\k_value2[31] ),
    .B(\hash/g[31] ),
    .Y(\hash/CA1/_0839_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3245_  (.A(\hash/CA1/_0838_ ),
    .B(\hash/CA1/_0839_ ),
    .Y(\hash/CA1/_0840_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3246_  (.A1(\hash/CA1/_1573_ ),
    .A2(\hash/CA1/_1570_ ),
    .B1(\hash/CA1/_1572_ ),
    .X(\hash/CA1/_0841_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3247_  (.A1(\hash/CA1/_1575_ ),
    .A2(\hash/CA1/_0841_ ),
    .B1(\hash/CA1/_1574_ ),
    .Y(\hash/CA1/_0842_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3248_  (.A(\hash/CA1/_0840_ ),
    .B(\hash/CA1/_0842_ ),
    .Y(\hash/CA1/_0843_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_3249_  (.A(\hash/CA1/_1576_ ),
    .B(\hash/CA1/_0843_ ),
    .X(\hash/CA1/_0844_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA1/_3250_  (.A_N(\hash/CA1/_0840_ ),
    .B(\hash/CA1/_0385_ ),
    .C(\hash/CA1/_1577_ ),
    .Y(\hash/CA1/_0845_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA1/_3251_  (.A0(\hash/CA1/_0844_ ),
    .A1(\hash/CA1/_0845_ ),
    .S(\hash/CA1/_0378_ ),
    .Y(\hash/CA1/_0846_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3252_  (.A(\hash/CA1/_0840_ ),
    .B(\hash/CA1/_0842_ ),
    .Y(\hash/CA1/_0847_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3253_  (.A(\hash/CA1/_1577_ ),
    .B(\hash/CA1/_0847_ ),
    .Y(\hash/CA1/_0848_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3254_  (.A(\hash/CA1/_1577_ ),
    .B(\hash/CA1/_1576_ ),
    .Y(\hash/CA1/_0849_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA1/_3255_  (.A0(\hash/CA1/_1576_ ),
    .A1(\hash/CA1/_0849_ ),
    .S(\hash/CA1/_0840_ ),
    .Y(\hash/CA1/_0850_ ));
 sky130_fd_sc_hd__o311ai_0 \hash/CA1/_3256_  (.A1(\hash/CA1/_1576_ ),
    .A2(\hash/CA1/_0385_ ),
    .A3(\hash/CA1/_0843_ ),
    .B1(\hash/CA1/_0848_ ),
    .C1(\hash/CA1/_0850_ ),
    .Y(\hash/CA1/_0851_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3257_  (.A(\hash/CA1/_0846_ ),
    .B(\hash/CA1/_0851_ ),
    .Y(\hash/p4[31] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3258_  (.A1(\hash/CA1/_1593_ ),
    .A2(\hash/CA1/_1590_ ),
    .B1(\hash/CA1/_1592_ ),
    .X(\hash/CA1/_0852_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3259_  (.A(\hash/CA1/_1585_ ),
    .Y(\hash/CA1/_0853_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3260_  (.A1(\hash/CA1/_1429_ ),
    .A2(\hash/CA1/_1581_ ),
    .B1(\hash/CA1/_1580_ ),
    .X(\hash/CA1/_0854_ ));
 sky130_fd_sc_hd__a21oi_2 \hash/CA1/_3261_  (.A1(\hash/CA1/_1583_ ),
    .A2(\hash/CA1/_0854_ ),
    .B1(\hash/CA1/_1582_ ),
    .Y(\hash/CA1/_0855_ ));
 sky130_fd_sc_hd__or3_4 \hash/CA1/_3262_  (.A(\hash/CA1/_1584_ ),
    .B(\hash/CA1/_1586_ ),
    .C(\hash/CA1/_1588_ ),
    .X(\hash/CA1/_0856_ ));
 sky130_fd_sc_hd__o21bai_4 \hash/CA1/_3263_  (.A1(\hash/CA1/_0853_ ),
    .A2(\hash/CA1/_0855_ ),
    .B1_N(\hash/CA1/_0856_ ),
    .Y(\hash/CA1/_0857_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_3264_  (.A1(\hash/CA1/_1587_ ),
    .A2(\hash/CA1/_1586_ ),
    .B1(\hash/CA1/_1589_ ),
    .Y(\hash/CA1/_0858_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3265_  (.A_N(\hash/CA1/_1588_ ),
    .B(\hash/CA1/_0858_ ),
    .Y(\hash/CA1/_0859_ ));
 sky130_fd_sc_hd__and4_1 \hash/CA1/_3266_  (.A(\hash/CA1/_1591_ ),
    .B(\hash/CA1/_1593_ ),
    .C(\hash/CA1/_1595_ ),
    .D(\hash/CA1/_0859_ ),
    .X(\hash/CA1/_0860_ ));
 sky130_fd_sc_hd__a221o_1 \hash/CA1/_3267_  (.A1(\hash/CA1/_1595_ ),
    .A2(\hash/CA1/_0852_ ),
    .B1(\hash/CA1/_0857_ ),
    .B2(\hash/CA1/_0860_ ),
    .C1(\hash/CA1/_1594_ ),
    .X(\hash/CA1/_0861_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3268_  (.A(\hash/CA1/_1597_ ),
    .B(\hash/CA1/_0861_ ),
    .X(\hash/p5[10] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3269_  (.A1(\hash/CA1/_1595_ ),
    .A2(\hash/CA1/_1594_ ),
    .B1(\hash/CA1/_1597_ ),
    .Y(\hash/CA1/_0862_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3270_  (.A1(\hash/CA1/_1428_ ),
    .A2(\hash/CA1/_1579_ ),
    .B1(\hash/CA1/_1578_ ),
    .Y(\hash/CA1/_0863_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3271_  (.A(\hash/CA1/_1581_ ),
    .B(\hash/CA1/_1583_ ),
    .C(\hash/CA1/_1585_ ),
    .Y(\hash/CA1/_0864_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3272_  (.A(\hash/CA1/_1585_ ),
    .B(\hash/CA1/_1582_ ),
    .Y(\hash/CA1/_0865_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3273_  (.A(\hash/CA1/_1583_ ),
    .B(\hash/CA1/_1585_ ),
    .C(\hash/CA1/_1580_ ),
    .Y(\hash/CA1/_0866_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA1/_3274_  (.A1(\hash/CA1/_0863_ ),
    .A2(\hash/CA1/_0864_ ),
    .B1(\hash/CA1/_0865_ ),
    .C1(\hash/CA1/_0866_ ),
    .Y(\hash/CA1/_0867_ ));
 sky130_fd_sc_hd__o2111a_1 \hash/CA1/_3275_  (.A1(\hash/CA1/_0856_ ),
    .A2(\hash/CA1/_0867_ ),
    .B1(\hash/CA1/_0859_ ),
    .C1(\hash/CA1/_1591_ ),
    .D1(\hash/CA1/_1593_ ),
    .X(\hash/CA1/_0868_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3276_  (.A(\hash/CA1/_1594_ ),
    .B(\hash/CA1/_0852_ ),
    .C(\hash/CA1/_0868_ ),
    .Y(\hash/CA1/_0869_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3277_  (.A(\hash/CA1/_1596_ ),
    .Y(\hash/CA1/_0870_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3278_  (.A1(\hash/CA1/_0862_ ),
    .A2(\hash/CA1/_0869_ ),
    .B1(\hash/CA1/_0870_ ),
    .X(\hash/CA1/_0871_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3279_  (.A(\hash/CA1/_1599_ ),
    .B(\hash/CA1/_0871_ ),
    .Y(\hash/p5[11] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3280_  (.A(\hash/CA1/_1597_ ),
    .B(\hash/CA1/_0861_ ),
    .Y(\hash/CA1/_0872_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3281_  (.A(\hash/CA1/_0870_ ),
    .B(\hash/CA1/_0872_ ),
    .Y(\hash/CA1/_0873_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3282_  (.A1(\hash/CA1/_1599_ ),
    .A2(\hash/CA1/_0873_ ),
    .B1(\hash/CA1/_1598_ ),
    .Y(\hash/CA1/_0874_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3283_  (.A(\hash/CA1/_1601_ ),
    .B(\hash/CA1/_0874_ ),
    .Y(\hash/p5[12] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3284_  (.A(\hash/CA1/_1599_ ),
    .B(\hash/CA1/_1601_ ),
    .Y(\hash/CA1/_0875_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3285_  (.A1(\hash/CA1/_1601_ ),
    .A2(\hash/CA1/_1598_ ),
    .B1(\hash/CA1/_1600_ ),
    .Y(\hash/CA1/_0876_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3286_  (.A1(\hash/CA1/_0871_ ),
    .A2(\hash/CA1/_0875_ ),
    .B1(\hash/CA1/_0876_ ),
    .X(\hash/CA1/_0877_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3287_  (.A(\hash/CA1/_1603_ ),
    .B(\hash/CA1/_0877_ ),
    .Y(\hash/p5[13] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3288_  (.A1(\hash/CA1/_1599_ ),
    .A2(\hash/CA1/_1596_ ),
    .B1(\hash/CA1/_1598_ ),
    .X(\hash/CA1/_0878_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3289_  (.A1(\hash/CA1/_1601_ ),
    .A2(\hash/CA1/_0878_ ),
    .B1(\hash/CA1/_1600_ ),
    .Y(\hash/CA1/_0879_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3290_  (.A1(\hash/CA1/_0872_ ),
    .A2(\hash/CA1/_0875_ ),
    .B1(\hash/CA1/_0879_ ),
    .Y(\hash/CA1/_0880_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3291_  (.A1(\hash/CA1/_1603_ ),
    .A2(\hash/CA1/_0880_ ),
    .B1(\hash/CA1/_1602_ ),
    .Y(\hash/CA1/_0881_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3292_  (.A(\hash/CA1/_1605_ ),
    .B(\hash/CA1/_0881_ ),
    .Y(\hash/p5[14] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3293_  (.A(\hash/CA1/_1603_ ),
    .Y(\hash/CA1/_0882_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3294_  (.A1(\hash/CA1/_0882_ ),
    .A2(\hash/CA1/_0877_ ),
    .B1_N(\hash/CA1/_1602_ ),
    .Y(\hash/CA1/_0883_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3295_  (.A1(\hash/CA1/_1605_ ),
    .A2(\hash/CA1/_0883_ ),
    .B1(\hash/CA1/_1604_ ),
    .Y(\hash/CA1/_0884_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3296_  (.A(\hash/CA1/_1607_ ),
    .B(\hash/CA1/_0884_ ),
    .Y(\hash/p5[15] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3297_  (.A(\hash/CA1/_1603_ ),
    .B(\hash/CA1/_1605_ ),
    .Y(\hash/CA1/_0885_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3298_  (.A(\hash/CA1/_1597_ ),
    .B(\hash/CA1/_1607_ ),
    .Y(\hash/CA1/_0886_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3299_  (.A(\hash/CA1/_0875_ ),
    .B(\hash/CA1/_0885_ ),
    .C(\hash/CA1/_0886_ ),
    .Y(\hash/CA1/_0887_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3300_  (.A1(\hash/CA1/_1605_ ),
    .A2(\hash/CA1/_1602_ ),
    .B1(\hash/CA1/_1604_ ),
    .Y(\hash/CA1/_0888_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3301_  (.A1(\hash/CA1/_0879_ ),
    .A2(\hash/CA1/_0885_ ),
    .B1(\hash/CA1/_0888_ ),
    .Y(\hash/CA1/_0889_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3302_  (.A1(\hash/CA1/_1607_ ),
    .A2(\hash/CA1/_0889_ ),
    .B1(\hash/CA1/_1606_ ),
    .Y(\hash/CA1/_0890_ ));
 sky130_fd_sc_hd__a21bo_1 \hash/CA1/_3303_  (.A1(\hash/CA1/_0861_ ),
    .A2(\hash/CA1/_0887_ ),
    .B1_N(\hash/CA1/_0890_ ),
    .X(\hash/CA1/_0891_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3304_  (.A(\hash/CA1/_1609_ ),
    .B(\hash/CA1/_0891_ ),
    .X(\hash/p5[16] ));
 sky130_fd_sc_hd__or3_1 \hash/CA1/_3306_  (.A(\hash/CA1/_1594_ ),
    .B(\hash/CA1/_1596_ ),
    .C(\hash/CA1/_0852_ ),
    .X(\hash/CA1/_0893_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA1/_3307_  (.A(\hash/CA1/_1603_ ),
    .B(\hash/CA1/_1605_ ),
    .C(\hash/CA1/_1607_ ),
    .Y(\hash/CA1/_0894_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_3308_  (.A1(\hash/CA1/_0870_ ),
    .A2(\hash/CA1/_0862_ ),
    .B1(\hash/CA1/_0875_ ),
    .C1(\hash/CA1/_0894_ ),
    .Y(\hash/CA1/_0895_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3309_  (.A1(\hash/CA1/_0868_ ),
    .A2(\hash/CA1/_0893_ ),
    .B1(\hash/CA1/_0895_ ),
    .Y(\hash/CA1/_0896_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3310_  (.A(\hash/CA1/_0888_ ),
    .B_N(\hash/CA1/_1607_ ),
    .Y(\hash/CA1/_0897_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3311_  (.A(\hash/CA1/_0876_ ),
    .B(\hash/CA1/_0894_ ),
    .Y(\hash/CA1/_0898_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA1/_3312_  (.A(\hash/CA1/_1606_ ),
    .B(\hash/CA1/_0897_ ),
    .C(\hash/CA1/_0898_ ),
    .Y(\hash/CA1/_0899_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA1/_3313_  (.A1(\hash/CA1/_0896_ ),
    .A2(\hash/CA1/_0899_ ),
    .B1_N(\hash/CA1/_1609_ ),
    .Y(\hash/CA1/_0900_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3314_  (.A(\hash/CA1/_1608_ ),
    .B(\hash/CA1/_0900_ ),
    .Y(\hash/CA1/_0901_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3315_  (.A(\hash/CA1/_1611_ ),
    .B(\hash/CA1/_0901_ ),
    .Y(\hash/p5[17] ));
 sky130_fd_sc_hd__a21o_2 \hash/CA1/_3316_  (.A1(\hash/CA1/_1609_ ),
    .A2(\hash/CA1/_0891_ ),
    .B1(\hash/CA1/_1608_ ),
    .X(\hash/CA1/_0902_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3317_  (.A1(\hash/CA1/_1611_ ),
    .A2(\hash/CA1/_0902_ ),
    .B1(\hash/CA1/_1610_ ),
    .Y(\hash/CA1/_0903_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3318_  (.A(\hash/CA1/_1613_ ),
    .B(\hash/CA1/_0903_ ),
    .Y(\hash/p5[18] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3319_  (.A1(\hash/CA1/_1608_ ),
    .A2(\hash/CA1/_0900_ ),
    .B1(\hash/CA1/_1611_ ),
    .Y(\hash/CA1/_0904_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3320_  (.A_N(\hash/CA1/_1610_ ),
    .B(\hash/CA1/_0904_ ),
    .Y(\hash/CA1/_0905_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3321_  (.A1(\hash/CA1/_1613_ ),
    .A2(\hash/CA1/_0905_ ),
    .B1(\hash/CA1/_1612_ ),
    .Y(\hash/CA1/_0906_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3322_  (.A(\hash/CA1/_1615_ ),
    .B(\hash/CA1/_0906_ ),
    .Y(\hash/p5[19] ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3323_  (.A1(\hash/CA1/_1615_ ),
    .A2(\hash/CA1/_1612_ ),
    .B1(\hash/CA1/_1614_ ),
    .Y(\hash/CA1/_0907_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3324_  (.A1(\hash/CA1/_1611_ ),
    .A2(\hash/CA1/_1608_ ),
    .B1(\hash/CA1/_1610_ ),
    .Y(\hash/CA1/_0908_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3325_  (.A(\hash/CA1/_0907_ ),
    .B(\hash/CA1/_0908_ ),
    .Y(\hash/CA1/_0909_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA1/_3326_  (.A1(\hash/CA1/_1609_ ),
    .A2(\hash/CA1/_1608_ ),
    .B1(\hash/CA1/_1611_ ),
    .X(\hash/CA1/_0910_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA1/_3327_  (.A(\hash/CA1/_1613_ ),
    .B(\hash/CA1/_1615_ ),
    .X(\hash/CA1/_0911_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3328_  (.A1(\hash/CA1/_1610_ ),
    .A2(\hash/CA1/_0910_ ),
    .B1(\hash/CA1/_0911_ ),
    .Y(\hash/CA1/_0912_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3329_  (.A(\hash/CA1/_0907_ ),
    .B(\hash/CA1/_0912_ ),
    .Y(\hash/CA1/_0913_ ));
 sky130_fd_sc_hd__o211a_4 \hash/CA1/_3330_  (.A1(\hash/CA1/_0891_ ),
    .A2(\hash/CA1/_0909_ ),
    .B1(\hash/CA1/_0913_ ),
    .C1(\hash/CA1/_1617_ ),
    .X(\hash/CA1/_0914_ ));
 sky130_fd_sc_hd__and2b_2 \hash/CA1/_3331_  (.A_N(\hash/CA1/_0891_ ),
    .B(\hash/CA1/_0908_ ),
    .X(\hash/CA1/_0915_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3332_  (.A1(\hash/CA1/_0912_ ),
    .A2(\hash/CA1/_0915_ ),
    .B1(\hash/CA1/_0907_ ),
    .Y(\hash/CA1/_0916_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3333_  (.A(\hash/CA1/_1617_ ),
    .B(\hash/CA1/_0916_ ),
    .Y(\hash/CA1/_0917_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3334_  (.A(\hash/CA1/_0914_ ),
    .B(\hash/CA1/_0917_ ),
    .Y(\hash/p5[20] ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3335_  (.A1(\hash/CA1/_1613_ ),
    .A2(\hash/CA1/_1610_ ),
    .B1(\hash/CA1/_1612_ ),
    .Y(\hash/CA1/_0918_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3336_  (.A(\hash/CA1/_0918_ ),
    .B_N(\hash/CA1/_1615_ ),
    .Y(\hash/CA1/_0919_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3337_  (.A1(\hash/CA1/_1614_ ),
    .A2(\hash/CA1/_0919_ ),
    .B1(\hash/CA1/_1617_ ),
    .Y(\hash/CA1/_0920_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/CA1/_3338_  (.A1(\hash/CA1/_1611_ ),
    .A2(\hash/CA1/_1617_ ),
    .A3(\hash/CA1/_1608_ ),
    .A4(\hash/CA1/_0911_ ),
    .B1(\hash/CA1/_1616_ ),
    .Y(\hash/CA1/_0921_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3339_  (.A(\hash/CA1/_0920_ ),
    .B(\hash/CA1/_0921_ ),
    .Y(\hash/CA1/_0922_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_3340_  (.A(\hash/CA1/_1609_ ),
    .B(\hash/CA1/_1611_ ),
    .C(\hash/CA1/_1617_ ),
    .D(\hash/CA1/_0911_ ),
    .Y(\hash/CA1/_0923_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3341_  (.A1(\hash/CA1/_0896_ ),
    .A2(\hash/CA1/_0899_ ),
    .B1(\hash/CA1/_0923_ ),
    .Y(\hash/CA1/_0924_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3342_  (.A(\hash/CA1/_0922_ ),
    .B(\hash/CA1/_0924_ ),
    .Y(\hash/CA1/_0925_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3343_  (.A(\hash/CA1/_1619_ ),
    .B(\hash/CA1/_0925_ ),
    .Y(\hash/p5[21] ));
 sky130_fd_sc_hd__or2_2 \hash/CA1/_3344_  (.A(\hash/CA1/_1616_ ),
    .B(\hash/CA1/_1618_ ),
    .X(\hash/CA1/_0926_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA1/_3345_  (.A1(\hash/CA1/_1619_ ),
    .A2(\hash/CA1/_1618_ ),
    .B1(\hash/CA1/_0914_ ),
    .B2(\hash/CA1/_0926_ ),
    .Y(\hash/CA1/_0927_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3346_  (.A(\hash/CA1/_1621_ ),
    .B(\hash/CA1/_0927_ ),
    .Y(\hash/p5[22] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3347_  (.A(\hash/CA1/_1619_ ),
    .B(\hash/CA1/_1621_ ),
    .Y(\hash/CA1/_0928_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3348_  (.A1(\hash/CA1/_1621_ ),
    .A2(\hash/CA1/_1618_ ),
    .B1(\hash/CA1/_1620_ ),
    .Y(\hash/CA1/_0929_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3349_  (.A1(\hash/CA1/_0925_ ),
    .A2(\hash/CA1/_0928_ ),
    .B1(\hash/CA1/_0929_ ),
    .Y(\hash/CA1/_0930_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3350_  (.A(\hash/CA1/_1623_ ),
    .B(\hash/CA1/_0930_ ),
    .X(\hash/p5[23] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3351_  (.A(\hash/CA1/_1621_ ),
    .Y(\hash/CA1/_0931_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3352_  (.A1(\hash/CA1/_0931_ ),
    .A2(\hash/CA1/_0927_ ),
    .B1_N(\hash/CA1/_1620_ ),
    .Y(\hash/CA1/_0932_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3353_  (.A1(\hash/CA1/_1623_ ),
    .A2(\hash/CA1/_0932_ ),
    .B1(\hash/CA1/_1622_ ),
    .Y(\hash/CA1/_0933_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3354_  (.A(\hash/CA1/_1625_ ),
    .B(\hash/CA1/_0933_ ),
    .Y(\hash/p5[24] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA1/_3355_  (.A1(\hash/CA1/_1623_ ),
    .A2(\hash/CA1/_0930_ ),
    .B1(\hash/CA1/_1622_ ),
    .X(\hash/CA1/_0934_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3356_  (.A1(\hash/CA1/_1625_ ),
    .A2(\hash/CA1/_0934_ ),
    .B1(\hash/CA1/_1624_ ),
    .Y(\hash/CA1/_0935_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3357_  (.A(\hash/CA1/_1627_ ),
    .B(\hash/CA1/_0935_ ),
    .Y(\hash/p5[25] ));
 sky130_fd_sc_hd__nand4_1 \hash/CA1/_3358_  (.A(\hash/CA1/_1619_ ),
    .B(\hash/CA1/_1621_ ),
    .C(\hash/CA1/_1623_ ),
    .D(\hash/CA1/_1625_ ),
    .Y(\hash/CA1/_0936_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3359_  (.A(\hash/CA1/_1627_ ),
    .B(\hash/CA1/_1629_ ),
    .Y(\hash/CA1/_0937_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3360_  (.A(\hash/CA1/_0936_ ),
    .B(\hash/CA1/_0937_ ),
    .Y(\hash/CA1/_0938_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3361_  (.A1(\hash/CA1/_1619_ ),
    .A2(\hash/CA1/_1616_ ),
    .B1(\hash/CA1/_1618_ ),
    .Y(\hash/CA1/_0939_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3362_  (.A(\hash/CA1/_0939_ ),
    .B_N(\hash/CA1/_1621_ ),
    .Y(\hash/CA1/_0940_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3363_  (.A1(\hash/CA1/_1620_ ),
    .A2(\hash/CA1/_0940_ ),
    .B1(\hash/CA1/_1623_ ),
    .Y(\hash/CA1/_0941_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3364_  (.A_N(\hash/CA1/_1622_ ),
    .B(\hash/CA1/_0941_ ),
    .Y(\hash/CA1/_0942_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3365_  (.A1(\hash/CA1/_1625_ ),
    .A2(\hash/CA1/_0942_ ),
    .B1(\hash/CA1/_1624_ ),
    .Y(\hash/CA1/_0943_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3366_  (.A(\hash/CA1/_1629_ ),
    .B(\hash/CA1/_1626_ ),
    .Y(\hash/CA1/_0944_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3367_  (.A1(\hash/CA1/_0943_ ),
    .A2(\hash/CA1/_0937_ ),
    .B1(\hash/CA1/_0944_ ),
    .Y(\hash/CA1/_0945_ ));
 sky130_fd_sc_hd__a21o_2 \hash/CA1/_3368_  (.A1(\hash/CA1/_0914_ ),
    .A2(\hash/CA1/_0938_ ),
    .B1(\hash/CA1/_0945_ ),
    .X(\hash/CA1/_0946_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3369_  (.A(\hash/CA1/_0914_ ),
    .Y(\hash/CA1/_0947_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3370_  (.A1(\hash/CA1/_0947_ ),
    .A2(\hash/CA1/_0936_ ),
    .B1(\hash/CA1/_0943_ ),
    .Y(\hash/CA1/_0948_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_3371_  (.A1(\hash/CA1/_1627_ ),
    .A2(\hash/CA1/_0948_ ),
    .B1(\hash/CA1/_1626_ ),
    .C1(\hash/CA1/_1629_ ),
    .Y(\hash/CA1/_0949_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3372_  (.A(\hash/CA1/_0946_ ),
    .B(\hash/CA1/_0949_ ),
    .Y(\hash/p5[26] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3373_  (.A(\hash/CA1/_1623_ ),
    .B(\hash/CA1/_1625_ ),
    .Y(\hash/CA1/_0950_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3374_  (.A(\hash/CA1/_0950_ ),
    .B(\hash/CA1/_0937_ ),
    .Y(\hash/CA1/_0951_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3375_  (.A1(\hash/CA1/_1625_ ),
    .A2(\hash/CA1/_1622_ ),
    .B1(\hash/CA1/_1624_ ),
    .Y(\hash/CA1/_0952_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3376_  (.A(\hash/CA1/_0952_ ),
    .B_N(\hash/CA1/_1627_ ),
    .Y(\hash/CA1/_0953_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3377_  (.A1(\hash/CA1/_1626_ ),
    .A2(\hash/CA1/_0953_ ),
    .B1(\hash/CA1/_1629_ ),
    .Y(\hash/CA1/_0954_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3378_  (.A_N(\hash/CA1/_1628_ ),
    .B(\hash/CA1/_0954_ ),
    .Y(\hash/CA1/_0955_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3379_  (.A1(\hash/CA1/_0930_ ),
    .A2(\hash/CA1/_0951_ ),
    .B1(\hash/CA1/_0955_ ),
    .Y(\hash/CA1/_0956_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3380_  (.A(\hash/CA1/_1631_ ),
    .B(\hash/CA1/_0956_ ),
    .Y(\hash/p5[27] ));
 sky130_fd_sc_hd__a2111oi_4 \hash/CA1/_3381_  (.A1(\hash/CA1/_0914_ ),
    .A2(\hash/CA1/_0938_ ),
    .B1(\hash/CA1/_0945_ ),
    .C1(\hash/CA1/_1630_ ),
    .D1(\hash/CA1/_1628_ ),
    .Y(\hash/CA1/_0957_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3382_  (.A1(\hash/CA1/_1631_ ),
    .A2(\hash/CA1/_1630_ ),
    .B1(\hash/CA1/_1633_ ),
    .Y(\hash/CA1/_0958_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3383_  (.A(\hash/CA1/_1633_ ),
    .B(\hash/CA1/_1630_ ),
    .Y(\hash/CA1/_0959_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3384_  (.A1(\hash/CA1/_1628_ ),
    .A2(\hash/CA1/_0946_ ),
    .B1(\hash/CA1/_1631_ ),
    .Y(\hash/CA1/_0960_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \hash/CA1/_3385_  (.A1_N(\hash/CA1/_0957_ ),
    .A2_N(\hash/CA1/_0958_ ),
    .B1(\hash/CA1/_0959_ ),
    .B2(\hash/CA1/_0960_ ),
    .Y(\hash/p5[28] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3386_  (.A(\hash/CA1/_1632_ ),
    .Y(\hash/CA1/_0961_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3387_  (.A(\hash/CA1/_1631_ ),
    .B(\hash/CA1/_0951_ ),
    .Y(\hash/CA1/_0962_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3388_  (.A(\hash/CA1/_0928_ ),
    .B(\hash/CA1/_0962_ ),
    .Y(\hash/CA1/_0963_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3389_  (.A1(\hash/CA1/_0922_ ),
    .A2(\hash/CA1/_0924_ ),
    .B1(\hash/CA1/_0963_ ),
    .Y(\hash/CA1/_0964_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3390_  (.A(\hash/CA1/_0929_ ),
    .B(\hash/CA1/_0962_ ),
    .Y(\hash/CA1/_0965_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_3391_  (.A1(\hash/CA1/_1631_ ),
    .A2(\hash/CA1/_0955_ ),
    .B1(\hash/CA1/_0965_ ),
    .C1(\hash/CA1/_1630_ ),
    .Y(\hash/CA1/_0966_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3392_  (.A1(\hash/CA1/_1633_ ),
    .A2(\hash/CA1/_1632_ ),
    .B1(\hash/CA1/_1635_ ),
    .Y(\hash/CA1/_0967_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_3393_  (.A1(\hash/CA1/_0961_ ),
    .A2(\hash/CA1/_0964_ ),
    .A3(\hash/CA1/_0966_ ),
    .B1(\hash/CA1/_0967_ ),
    .Y(\hash/CA1/_0968_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3394_  (.A(\hash/CA1/_0964_ ),
    .B(\hash/CA1/_0966_ ),
    .Y(\hash/CA1/_0969_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA1/_3395_  (.A1(\hash/CA1/_1633_ ),
    .A2(\hash/CA1/_0969_ ),
    .B1(\hash/CA1/_1632_ ),
    .C1(\hash/CA1/_1635_ ),
    .Y(\hash/CA1/_0970_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3396_  (.A(\hash/CA1/_0968_ ),
    .B(\hash/CA1/_0970_ ),
    .Y(\hash/p5[29] ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3397_  (.A(\hash/CA1/_1429_ ),
    .B(\hash/CA1/_1581_ ),
    .X(\hash/p5[2] ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA1/_3398_  (.A1(\hash/CA1/_0957_ ),
    .A2(\hash/CA1/_0958_ ),
    .B1(\hash/CA1/_0961_ ),
    .Y(\hash/CA1/_0971_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3399_  (.A1(\hash/CA1/_1635_ ),
    .A2(\hash/CA1/_0971_ ),
    .B1(\hash/CA1/_1634_ ),
    .Y(\hash/CA1/_0972_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3400_  (.A(\hash/CA1/_1637_ ),
    .B(\hash/CA1/_0972_ ),
    .Y(\hash/p5[30] ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA1/_3401_  (.A_N(\hash/CA1/_1636_ ),
    .B(\hash/c[31] ),
    .Y(\hash/CA1/_0973_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA1/_3402_  (.A(\hash/c[31] ),
    .B_N(\hash/CA1/_1637_ ),
    .Y(\hash/CA1/_0974_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA1/_3403_  (.A(\hash/CA1/_0968_ ),
    .B(\hash/CA1/_0974_ ),
    .Y(\hash/CA1/_0975_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3404_  (.A(\hash/c[31] ),
    .Y(\hash/CA1/_0976_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3405_  (.A(\hash/CA1/_1637_ ),
    .B(\hash/CA1/_0973_ ),
    .Y(\hash/CA1/_0977_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA1/_3406_  (.A1(\hash/CA1/_0976_ ),
    .A2(\hash/CA1/_1636_ ),
    .B1(\hash/CA1/_1634_ ),
    .B2(\hash/CA1/_0974_ ),
    .C1(\hash/CA1/_0977_ ),
    .Y(\hash/CA1/_0978_ ));
 sky130_fd_sc_hd__o311ai_0 \hash/CA1/_3407_  (.A1(\hash/CA1/_1634_ ),
    .A2(\hash/CA1/_0968_ ),
    .A3(\hash/CA1/_0973_ ),
    .B1(\hash/CA1/_0975_ ),
    .C1(\hash/CA1/_0978_ ),
    .Y(\hash/CA1/_0979_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3408_  (.A(\hash/p4[31] ),
    .B(\hash/CA1/_0979_ ),
    .X(\hash/p5[31] ));
 sky130_fd_sc_hd__inv_1 \hash/CA1/_3409_  (.A(\hash/CA1/_1581_ ),
    .Y(\hash/CA1/_0980_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3410_  (.A1(\hash/CA1/_0980_ ),
    .A2(\hash/CA1/_0863_ ),
    .B1_N(\hash/CA1/_1580_ ),
    .Y(\hash/CA1/_0981_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA1/_3411_  (.A(\hash/CA1/_1583_ ),
    .B(\hash/CA1/_0981_ ),
    .X(\hash/p5[3] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3412_  (.A(\hash/CA1/_1585_ ),
    .B(\hash/CA1/_0855_ ),
    .Y(\hash/p5[4] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3413_  (.A(\hash/CA1/_1584_ ),
    .B(\hash/CA1/_0867_ ),
    .Y(\hash/CA1/_0982_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3414_  (.A(\hash/CA1/_1587_ ),
    .B(\hash/CA1/_0982_ ),
    .Y(\hash/p5[5] ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA1/_3415_  (.A1(\hash/CA1/_0853_ ),
    .A2(\hash/CA1/_0855_ ),
    .B1_N(\hash/CA1/_1584_ ),
    .Y(\hash/CA1/_0983_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA1/_3416_  (.A1(\hash/CA1/_1587_ ),
    .A2(\hash/CA1/_0983_ ),
    .B1(\hash/CA1/_1586_ ),
    .Y(\hash/CA1/_0984_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3417_  (.A(\hash/CA1/_1589_ ),
    .B(\hash/CA1/_0984_ ),
    .Y(\hash/p5[6] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA1/_3418_  (.A1(\hash/CA1/_0856_ ),
    .A2(\hash/CA1/_0867_ ),
    .B1(\hash/CA1/_0859_ ),
    .Y(\hash/CA1/_0985_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3419_  (.A(\hash/CA1/_1591_ ),
    .B(\hash/CA1/_0985_ ),
    .Y(\hash/p5[7] ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA1/_3420_  (.A1(\hash/CA1/_1591_ ),
    .A2(\hash/CA1/_0857_ ),
    .A3(\hash/CA1/_0859_ ),
    .B1(\hash/CA1/_1590_ ),
    .Y(\hash/CA1/_0986_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3421_  (.A(\hash/CA1/_1593_ ),
    .B(\hash/CA1/_0986_ ),
    .Y(\hash/p5[8] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA1/_3422_  (.A(\hash/CA1/_0852_ ),
    .B(\hash/CA1/_0868_ ),
    .Y(\hash/CA1/_0987_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA1/_3423_  (.A(\hash/CA1/_1595_ ),
    .B(\hash/CA1/_0987_ ),
    .Y(\hash/p5[9] ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3424_  (.A(\hash/g[0] ),
    .B(\k_value2[0] ),
    .CIN(\w_value2[0] ),
    .COUT(\hash/CA1/_0988_ ),
    .SUM(\hash/p4[0] ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3425_  (.A(\hash/g[1] ),
    .B(\k_value2[1] ),
    .CIN(\w_value2[1] ),
    .COUT(\hash/CA1/_0989_ ),
    .SUM(\hash/CA1/_0990_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3426_  (.A(\hash/g[2] ),
    .B(\k_value2[2] ),
    .CIN(\w_value2[2] ),
    .COUT(\hash/CA1/_0991_ ),
    .SUM(\hash/CA1/_0992_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3427_  (.A(\hash/CA1/_0993_ ),
    .B(\hash/CA1/_0994_ ),
    .CIN(\hash/CA1/_0995_ ),
    .COUT(\hash/CA1/_0996_ ),
    .SUM(\hash/CA1/_0997_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3428_  (.A(\hash/g[3] ),
    .B(\k_value2[3] ),
    .CIN(\w_value2[3] ),
    .COUT(\hash/CA1/_0998_ ),
    .SUM(\hash/CA1/_0999_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3429_  (.A(\hash/g[4] ),
    .B(\k_value2[4] ),
    .CIN(\w_value2[4] ),
    .COUT(\hash/CA1/_1000_ ),
    .SUM(\hash/CA1/_1001_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3430_  (.A(\hash/g[5] ),
    .B(\k_value2[5] ),
    .CIN(\w_value2[5] ),
    .COUT(\hash/CA1/_1002_ ),
    .SUM(\hash/CA1/_1003_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3431_  (.A(\hash/g[6] ),
    .B(\k_value2[6] ),
    .CIN(\w_value2[6] ),
    .COUT(\hash/CA1/_1004_ ),
    .SUM(\hash/CA1/_1005_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3432_  (.A(\hash/g[7] ),
    .B(\k_value2[7] ),
    .CIN(\w_value2[7] ),
    .COUT(\hash/CA1/_1006_ ),
    .SUM(\hash/CA1/_1007_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3433_  (.A(\hash/g[8] ),
    .B(\k_value2[8] ),
    .CIN(\w_value2[8] ),
    .COUT(\hash/CA1/_1008_ ),
    .SUM(\hash/CA1/_1009_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3434_  (.A(\hash/g[9] ),
    .B(\k_value2[9] ),
    .CIN(\w_value2[9] ),
    .COUT(\hash/CA1/_1010_ ),
    .SUM(\hash/CA1/_1011_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3435_  (.A(\hash/g[10] ),
    .B(\k_value2[10] ),
    .CIN(\w_value2[10] ),
    .COUT(\hash/CA1/_1012_ ),
    .SUM(\hash/CA1/_1013_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3436_  (.A(\hash/g[11] ),
    .B(\k_value2[11] ),
    .CIN(\w_value2[11] ),
    .COUT(\hash/CA1/_1014_ ),
    .SUM(\hash/CA1/_1015_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3437_  (.A(\hash/g[12] ),
    .B(\k_value2[12] ),
    .CIN(\w_value2[12] ),
    .COUT(\hash/CA1/_1016_ ),
    .SUM(\hash/CA1/_1017_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3438_  (.A(\hash/g[13] ),
    .B(\k_value2[13] ),
    .CIN(\w_value2[13] ),
    .COUT(\hash/CA1/_1018_ ),
    .SUM(\hash/CA1/_1019_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3439_  (.A(\hash/g[14] ),
    .B(\k_value2[14] ),
    .CIN(\w_value2[14] ),
    .COUT(\hash/CA1/_1020_ ),
    .SUM(\hash/CA1/_1021_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3440_  (.A(\hash/g[15] ),
    .B(\k_value2[15] ),
    .CIN(\w_value2[15] ),
    .COUT(\hash/CA1/_1022_ ),
    .SUM(\hash/CA1/_1023_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3441_  (.A(\hash/g[16] ),
    .B(\k_value2[16] ),
    .CIN(\w_value2[16] ),
    .COUT(\hash/CA1/_1024_ ),
    .SUM(\hash/CA1/_1025_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3442_  (.A(\hash/g[17] ),
    .B(\k_value2[17] ),
    .CIN(\w_value2[17] ),
    .COUT(\hash/CA1/_1026_ ),
    .SUM(\hash/CA1/_1027_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3443_  (.A(\hash/g[18] ),
    .B(\k_value2[18] ),
    .CIN(\w_value2[18] ),
    .COUT(\hash/CA1/_1028_ ),
    .SUM(\hash/CA1/_1029_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3444_  (.A(\hash/g[19] ),
    .B(\k_value2[19] ),
    .CIN(\w_value2[19] ),
    .COUT(\hash/CA1/_1030_ ),
    .SUM(\hash/CA1/_1031_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3445_  (.A(\hash/g[20] ),
    .B(\k_value2[20] ),
    .CIN(\w_value2[20] ),
    .COUT(\hash/CA1/_1032_ ),
    .SUM(\hash/CA1/_1033_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3446_  (.A(\hash/g[21] ),
    .B(\k_value2[21] ),
    .CIN(\w_value2[21] ),
    .COUT(\hash/CA1/_1034_ ),
    .SUM(\hash/CA1/_1035_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3447_  (.A(\hash/g[22] ),
    .B(\k_value2[22] ),
    .CIN(\w_value2[22] ),
    .COUT(\hash/CA1/_1036_ ),
    .SUM(\hash/CA1/_1037_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3448_  (.A(\hash/g[23] ),
    .B(\k_value2[23] ),
    .CIN(\w_value2[23] ),
    .COUT(\hash/CA1/_1038_ ),
    .SUM(\hash/CA1/_1039_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3449_  (.A(\hash/g[24] ),
    .B(\k_value2[24] ),
    .CIN(\w_value2[24] ),
    .COUT(\hash/CA1/_1040_ ),
    .SUM(\hash/CA1/_1041_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3450_  (.A(\hash/g[25] ),
    .B(\k_value2[25] ),
    .CIN(\w_value2[25] ),
    .COUT(\hash/CA1/_1042_ ),
    .SUM(\hash/CA1/_1043_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3451_  (.A(\hash/g[26] ),
    .B(\k_value2[26] ),
    .CIN(\w_value2[26] ),
    .COUT(\hash/CA1/_1044_ ),
    .SUM(\hash/CA1/_1045_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3452_  (.A(\hash/g[27] ),
    .B(\k_value2[27] ),
    .CIN(\w_value2[27] ),
    .COUT(\hash/CA1/_1046_ ),
    .SUM(\hash/CA1/_1047_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3453_  (.A(\hash/g[28] ),
    .B(\k_value2[28] ),
    .CIN(\w_value2[28] ),
    .COUT(\hash/CA1/_1048_ ),
    .SUM(\hash/CA1/_1049_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3454_  (.A(\hash/g[29] ),
    .B(\k_value2[29] ),
    .CIN(\w_value2[29] ),
    .COUT(\hash/CA1/_1050_ ),
    .SUM(\hash/CA1/_1051_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3455_  (.A(\hash/g[30] ),
    .B(\k_value2[30] ),
    .CIN(\w_value2[30] ),
    .COUT(\hash/CA1/_1052_ ),
    .SUM(\hash/CA1/_1053_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3456_  (.A(\hash/CA1/_1054_ ),
    .B(\hash/CA1/_1055_ ),
    .CIN(\hash/CA1/_1056_ ),
    .COUT(\hash/CA1/_1057_ ),
    .SUM(\hash/CA1/_1058_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3457_  (.A(\hash/CA1/_1059_ ),
    .B(\hash/CA1/_1060_ ),
    .CIN(\hash/CA1/_1061_ ),
    .COUT(\hash/CA1/_1062_ ),
    .SUM(\hash/CA1/_1063_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3458_  (.A(\hash/h[1] ),
    .B(\hash/CA1/_1064_ ),
    .CIN(\hash/CA1/_1065_ ),
    .COUT(\hash/CA1/_1066_ ),
    .SUM(\hash/CA1/_1067_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3459_  (.A(\hash/h[2] ),
    .B(\hash/CA1/_1068_ ),
    .CIN(\hash/CA1/_1069_ ),
    .COUT(\hash/CA1/_1070_ ),
    .SUM(\hash/CA1/_1071_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3460_  (.A(\hash/h[3] ),
    .B(\hash/CA1/_1072_ ),
    .CIN(\hash/CA1/_1073_ ),
    .COUT(\hash/CA1/_1074_ ),
    .SUM(\hash/CA1/_1075_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3461_  (.A(\hash/CA1/_1076_ ),
    .B(\hash/CA1/_1077_ ),
    .CIN(\hash/CA1/_1078_ ),
    .COUT(\hash/CA1/_1079_ ),
    .SUM(\hash/CA1/_1080_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3462_  (.A(\hash/h[5] ),
    .B(\hash/CA1/_1081_ ),
    .CIN(\hash/CA1/_1082_ ),
    .COUT(\hash/CA1/_1083_ ),
    .SUM(\hash/CA1/_1084_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3463_  (.A(\hash/h[6] ),
    .B(\hash/CA1/_1085_ ),
    .CIN(\hash/CA1/_1086_ ),
    .COUT(\hash/CA1/_1087_ ),
    .SUM(\hash/CA1/_1088_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3464_  (.A(\hash/h[7] ),
    .B(\hash/CA1/_1089_ ),
    .CIN(\hash/CA1/_1090_ ),
    .COUT(\hash/CA1/_1091_ ),
    .SUM(\hash/CA1/_1092_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3465_  (.A(\hash/h[8] ),
    .B(\hash/CA1/_1093_ ),
    .CIN(\hash/CA1/_1094_ ),
    .COUT(\hash/CA1/_1095_ ),
    .SUM(\hash/CA1/_1096_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3466_  (.A(\hash/CA1/_1099_ ),
    .B(\hash/CA1/_1100_ ),
    .CIN(\hash/CA1/_1101_ ),
    .COUT(\hash/CA1/_1102_ ),
    .SUM(\hash/CA1/_1103_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3467_  (.A(\hash/CA1/_1104_ ),
    .B(\hash/CA1/_1105_ ),
    .CIN(\hash/CA1/_1106_ ),
    .COUT(\hash/CA1/_1107_ ),
    .SUM(\hash/CA1/_1108_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3468_  (.A(\hash/CA1/_1109_ ),
    .B(\hash/CA1/_1110_ ),
    .CIN(\hash/CA1/_1111_ ),
    .COUT(\hash/CA1/_1112_ ),
    .SUM(\hash/CA1/_1113_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3469_  (.A(\hash/CA1/_1114_ ),
    .B(\hash/CA1/_1115_ ),
    .CIN(\hash/CA1/_1116_ ),
    .COUT(\hash/CA1/_1117_ ),
    .SUM(\hash/CA1/_1118_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3470_  (.A(\hash/CA1/_1119_ ),
    .B(\hash/CA1/_1120_ ),
    .CIN(\hash/CA1/_1121_ ),
    .COUT(\hash/CA1/_1122_ ),
    .SUM(\hash/CA1/_1123_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3471_  (.A(\hash/CA1/_1124_ ),
    .B(\hash/CA1/_1125_ ),
    .CIN(\hash/CA1/_1126_ ),
    .COUT(\hash/CA1/_1127_ ),
    .SUM(\hash/CA1/_1128_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3472_  (.A(\hash/h[15] ),
    .B(\hash/CA1/_1129_ ),
    .CIN(\hash/CA1/_1130_ ),
    .COUT(\hash/CA1/_1131_ ),
    .SUM(\hash/CA1/_1132_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3473_  (.A(\hash/CA1/_1135_ ),
    .B(\hash/CA1/_1136_ ),
    .CIN(\hash/CA1/_1137_ ),
    .COUT(\hash/CA1/_1138_ ),
    .SUM(\hash/CA1/_1139_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3474_  (.A(\hash/CA1/_1140_ ),
    .B(\hash/CA1/_1141_ ),
    .CIN(\hash/CA1/_1142_ ),
    .COUT(\hash/CA1/_1143_ ),
    .SUM(\hash/CA1/_1144_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3475_  (.A(\hash/CA1/_1145_ ),
    .B(\hash/CA1/_1146_ ),
    .CIN(\hash/CA1/_1147_ ),
    .COUT(\hash/CA1/_1148_ ),
    .SUM(\hash/CA1/_1149_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3476_  (.A(\hash/CA1/_1150_ ),
    .B(\hash/CA1/_1151_ ),
    .CIN(\hash/CA1/_1152_ ),
    .COUT(\hash/CA1/_1153_ ),
    .SUM(\hash/CA1/_1154_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3477_  (.A(\hash/CA1/_1155_ ),
    .B(\hash/CA1/_1156_ ),
    .CIN(\hash/CA1/_1157_ ),
    .COUT(\hash/CA1/_1158_ ),
    .SUM(\hash/CA1/_1159_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3478_  (.A(\hash/CA1/_1160_ ),
    .B(\hash/CA1/_1161_ ),
    .CIN(\hash/CA1/_1162_ ),
    .COUT(\hash/CA1/_1163_ ),
    .SUM(\hash/CA1/_1164_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3479_  (.A(\hash/CA1/_1165_ ),
    .B(\hash/CA1/_1166_ ),
    .CIN(\hash/CA1/_1167_ ),
    .COUT(\hash/CA1/_1168_ ),
    .SUM(\hash/CA1/_1169_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3480_  (.A(\hash/CA1/_1170_ ),
    .B(\hash/CA1/_1171_ ),
    .CIN(\hash/CA1/_1172_ ),
    .COUT(\hash/CA1/_1173_ ),
    .SUM(\hash/CA1/_1174_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3481_  (.A(\hash/CA1/_1175_ ),
    .B(\hash/CA1/_1176_ ),
    .CIN(\hash/CA1/_1177_ ),
    .COUT(\hash/CA1/_1178_ ),
    .SUM(\hash/CA1/_1179_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3482_  (.A(\hash/CA1/_1180_ ),
    .B(\hash/CA1/_1181_ ),
    .CIN(\hash/CA1/_1182_ ),
    .COUT(\hash/CA1/_1183_ ),
    .SUM(\hash/CA1/_1184_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3483_  (.A(\hash/CA1/_1185_ ),
    .B(\hash/CA1/_1186_ ),
    .CIN(\hash/CA1/_1187_ ),
    .COUT(\hash/CA1/_1188_ ),
    .SUM(\hash/CA1/_1189_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3484_  (.A(\hash/h[27] ),
    .B(\hash/CA1/_1190_ ),
    .CIN(\hash/CA1/_1191_ ),
    .COUT(\hash/CA1/_1192_ ),
    .SUM(\hash/CA1/_1193_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3485_  (.A(\hash/h[28] ),
    .B(\hash/CA1/_1196_ ),
    .CIN(\hash/CA1/_1197_ ),
    .COUT(\hash/CA1/_1198_ ),
    .SUM(\hash/CA1/_1199_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3486_  (.A(\hash/h[29] ),
    .B(\hash/CA1/_1202_ ),
    .CIN(\hash/CA1/_1203_ ),
    .COUT(\hash/CA1/_1204_ ),
    .SUM(\hash/CA1/_1205_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3487_  (.A(\hash/h[30] ),
    .B(\hash/CA1/_1209_ ),
    .CIN(\hash/CA1/_1210_ ),
    .COUT(\hash/CA1/_1211_ ),
    .SUM(\hash/CA1/_1212_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3488_  (.A(\hash/CA1/_1213_ ),
    .B(\hash/CA1/_1214_ ),
    .CIN(\hash/CA1/_1215_ ),
    .COUT(\hash/CA1/_1216_ ),
    .SUM(\hash/CA1/_1217_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3489_  (.A(\hash/CA1/_1218_ ),
    .B(\hash/CA1/_1219_ ),
    .CIN(\hash/CA1/_1058_ ),
    .COUT(\hash/CA1/_1220_ ),
    .SUM(\hash/CA1/_1221_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3490_  (.A(\hash/CA1/_1063_ ),
    .B(\hash/CA1/_1216_ ),
    .CIN(\hash/CA1/_1221_ ),
    .COUT(\hash/CA1/_1222_ ),
    .SUM(\hash/CA1/_1223_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3491_  (.A(\hash/CA1/_1224_ ),
    .B(\hash/CA1/_1225_ ),
    .CIN(\hash/CA1/_1226_ ),
    .COUT(\hash/CA1/_1227_ ),
    .SUM(\hash/CA1/_1228_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3492_  (.A(\hash/CA1/_1069_ ),
    .B(\hash/CA1/_1229_ ),
    .CIN(\hash/CA1/_1230_ ),
    .COUT(\hash/CA1/_1231_ ),
    .SUM(\hash/CA1/_1232_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3493_  (.A(\hash/CA1/_1233_ ),
    .B(\hash/CA1/_1234_ ),
    .CIN(\hash/CA1/_1235_ ),
    .COUT(\hash/CA1/_1236_ ),
    .SUM(\hash/CA1/_1237_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3494_  (.A(\hash/CA1/_1072_ ),
    .B(\hash/CA1/_1238_ ),
    .CIN(\hash/CA1/_1239_ ),
    .COUT(\hash/CA1/_1240_ ),
    .SUM(\hash/CA1/_1241_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3495_  (.A(\hash/d[4] ),
    .B(\hash/h[4] ),
    .CIN(\hash/CA1/_1242_ ),
    .COUT(\hash/CA1/_1243_ ),
    .SUM(\hash/CA1/_1244_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3496_  (.A(\hash/CA1/_1245_ ),
    .B(\hash/CA1/_1246_ ),
    .CIN(\hash/CA1/_1244_ ),
    .COUT(\hash/CA1/_1247_ ),
    .SUM(\hash/CA1/_1248_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3497_  (.A(\hash/d[5] ),
    .B(\hash/h[5] ),
    .CIN(\hash/CA1/_1082_ ),
    .COUT(\hash/CA1/_1249_ ),
    .SUM(\hash/CA1/_1250_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3498_  (.A(\hash/CA1/_1251_ ),
    .B(\hash/CA1/_1252_ ),
    .CIN(\hash/CA1/_1253_ ),
    .COUT(\hash/CA1/_1254_ ),
    .SUM(\hash/CA1/_1255_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3499_  (.A(\hash/d[6] ),
    .B(\hash/h[6] ),
    .CIN(\hash/CA1/_1086_ ),
    .COUT(\hash/CA1/_1256_ ),
    .SUM(\hash/CA1/_1257_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3500_  (.A(\hash/CA1/_1258_ ),
    .B(\hash/CA1/_1259_ ),
    .CIN(\hash/CA1/_1260_ ),
    .COUT(\hash/CA1/_1261_ ),
    .SUM(\hash/CA1/_1262_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3501_  (.A(\hash/d[7] ),
    .B(\hash/h[7] ),
    .CIN(\hash/CA1/_1090_ ),
    .COUT(\hash/CA1/_1263_ ),
    .SUM(\hash/CA1/_1264_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3502_  (.A(\hash/CA1/_1265_ ),
    .B(\hash/CA1/_1266_ ),
    .CIN(\hash/CA1/_1267_ ),
    .COUT(\hash/CA1/_1268_ ),
    .SUM(\hash/CA1/_1269_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3503_  (.A(\hash/CA1/_1270_ ),
    .B(\hash/CA1/_1098_ ),
    .CIN(\hash/CA1/_1097_ ),
    .COUT(\hash/CA1/_1271_ ),
    .SUM(\hash/CA1/_1272_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3504_  (.A(\hash/CA1/_1094_ ),
    .B(\hash/CA1/_1263_ ),
    .CIN(\hash/CA1/_1273_ ),
    .COUT(\hash/CA1/_1274_ ),
    .SUM(\hash/CA1/_1275_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3505_  (.A(\hash/d[9] ),
    .B(\hash/h[9] ),
    .CIN(\hash/CA1/_1276_ ),
    .COUT(\hash/CA1/_1277_ ),
    .SUM(\hash/CA1/_1278_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3506_  (.A(\hash/CA1/_1101_ ),
    .B(\hash/CA1/_1279_ ),
    .CIN(\hash/CA1/_1271_ ),
    .COUT(\hash/CA1/_1280_ ),
    .SUM(\hash/CA1/_1281_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3507_  (.A(\hash/d[10] ),
    .B(\hash/h[10] ),
    .CIN(\hash/CA1/_1282_ ),
    .COUT(\hash/CA1/_1283_ ),
    .SUM(\hash/CA1/_1284_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3508_  (.A(\hash/CA1/_1106_ ),
    .B(\hash/CA1/_1285_ ),
    .CIN(\hash/CA1/_1286_ ),
    .COUT(\hash/CA1/_1287_ ),
    .SUM(\hash/CA1/_1288_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3509_  (.A(\hash/d[11] ),
    .B(\hash/h[11] ),
    .CIN(\hash/CA1/_1289_ ),
    .COUT(\hash/CA1/_1290_ ),
    .SUM(\hash/CA1/_1291_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3510_  (.A(\hash/CA1/_1292_ ),
    .B(\hash/CA1/_1293_ ),
    .CIN(\hash/CA1/_1111_ ),
    .COUT(\hash/CA1/_1294_ ),
    .SUM(\hash/CA1/_1295_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3511_  (.A(\hash/d[12] ),
    .B(\hash/h[12] ),
    .CIN(\hash/CA1/_1296_ ),
    .COUT(\hash/CA1/_1297_ ),
    .SUM(\hash/CA1/_1298_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3512_  (.A(\hash/CA1/_1299_ ),
    .B(\hash/CA1/_1300_ ),
    .CIN(\hash/CA1/_1116_ ),
    .COUT(\hash/CA1/_1301_ ),
    .SUM(\hash/CA1/_1302_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3513_  (.A(\hash/d[13] ),
    .B(\hash/h[13] ),
    .CIN(\hash/CA1/_1303_ ),
    .COUT(\hash/CA1/_1304_ ),
    .SUM(\hash/CA1/_1305_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3514_  (.A(\hash/CA1/_1306_ ),
    .B(\hash/CA1/_1297_ ),
    .CIN(\hash/CA1/_1305_ ),
    .COUT(\hash/CA1/_1307_ ),
    .SUM(\hash/CA1/_1308_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3515_  (.A(\hash/d[14] ),
    .B(\hash/h[14] ),
    .CIN(\hash/CA1/_1309_ ),
    .COUT(\hash/CA1/_1310_ ),
    .SUM(\hash/CA1/_1311_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3516_  (.A(\hash/CA1/_1304_ ),
    .B(\hash/CA1/_1312_ ),
    .CIN(\hash/CA1/_1311_ ),
    .COUT(\hash/CA1/_1313_ ),
    .SUM(\hash/CA1/_1314_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3517_  (.A(\hash/CA1/_1315_ ),
    .B(\hash/CA1/_1134_ ),
    .CIN(\hash/CA1/_1133_ ),
    .COUT(\hash/CA1/_1316_ ),
    .SUM(\hash/CA1/_1317_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3518_  (.A(\hash/CA1/_1129_ ),
    .B(\hash/CA1/_1310_ ),
    .CIN(\hash/CA1/_1318_ ),
    .COUT(\hash/CA1/_1319_ ),
    .SUM(\hash/CA1/_1320_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3519_  (.A(\hash/d[16] ),
    .B(\hash/h[16] ),
    .CIN(\hash/CA1/_1321_ ),
    .COUT(\hash/CA1/_1322_ ),
    .SUM(\hash/CA1/_1323_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3520_  (.A(\hash/CA1/_1137_ ),
    .B(\hash/CA1/_1324_ ),
    .CIN(\hash/CA1/_1316_ ),
    .COUT(\hash/CA1/_1325_ ),
    .SUM(\hash/CA1/_1326_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3521_  (.A(\hash/d[17] ),
    .B(\hash/h[17] ),
    .CIN(\hash/CA1/_1327_ ),
    .COUT(\hash/CA1/_1328_ ),
    .SUM(\hash/CA1/_1329_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3522_  (.A(\hash/CA1/_1330_ ),
    .B(\hash/CA1/_1329_ ),
    .CIN(\hash/CA1/_1322_ ),
    .COUT(\hash/CA1/_1331_ ),
    .SUM(\hash/CA1/_1332_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3523_  (.A(\hash/d[18] ),
    .B(\hash/h[18] ),
    .CIN(\hash/CA1/_1333_ ),
    .COUT(\hash/CA1/_1334_ ),
    .SUM(\hash/CA1/_1335_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3524_  (.A(\hash/CA1/_1328_ ),
    .B(\hash/CA1/_1335_ ),
    .CIN(\hash/CA1/_1336_ ),
    .COUT(\hash/CA1/_1337_ ),
    .SUM(\hash/CA1/_1338_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3525_  (.A(\hash/d[19] ),
    .B(\hash/h[19] ),
    .CIN(\hash/CA1/_1339_ ),
    .COUT(\hash/CA1/_1340_ ),
    .SUM(\hash/CA1/_1341_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3526_  (.A(\hash/CA1/_1342_ ),
    .B(\hash/CA1/_1341_ ),
    .CIN(\hash/CA1/_1334_ ),
    .COUT(\hash/CA1/_1343_ ),
    .SUM(\hash/CA1/_1344_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3527_  (.A(\hash/d[20] ),
    .B(\hash/h[20] ),
    .CIN(\hash/CA1/_1345_ ),
    .COUT(\hash/CA1/_1346_ ),
    .SUM(\hash/CA1/_1347_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3528_  (.A(\hash/CA1/_1348_ ),
    .B(\hash/CA1/_1349_ ),
    .CIN(\hash/CA1/_1157_ ),
    .COUT(\hash/CA1/_1350_ ),
    .SUM(\hash/CA1/_1351_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3529_  (.A(\hash/d[21] ),
    .B(\hash/h[21] ),
    .CIN(\hash/CA1/_1352_ ),
    .COUT(\hash/CA1/_1353_ ),
    .SUM(\hash/CA1/_1354_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3530_  (.A(\hash/CA1/_1355_ ),
    .B(\hash/CA1/_1346_ ),
    .CIN(\hash/CA1/_1354_ ),
    .COUT(\hash/CA1/_1356_ ),
    .SUM(\hash/CA1/_1357_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3531_  (.A(\hash/d[22] ),
    .B(\hash/h[22] ),
    .CIN(\hash/CA1/_1358_ ),
    .COUT(\hash/CA1/_1359_ ),
    .SUM(\hash/CA1/_1360_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3532_  (.A(\hash/CA1/_1361_ ),
    .B(\hash/CA1/_1353_ ),
    .CIN(\hash/CA1/_1360_ ),
    .COUT(\hash/CA1/_1362_ ),
    .SUM(\hash/CA1/_1363_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3533_  (.A(\hash/d[23] ),
    .B(\hash/h[23] ),
    .CIN(\hash/CA1/_1364_ ),
    .COUT(\hash/CA1/_1365_ ),
    .SUM(\hash/CA1/_1366_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3534_  (.A(\hash/CA1/_1367_ ),
    .B(\hash/CA1/_1368_ ),
    .CIN(\hash/CA1/_1172_ ),
    .COUT(\hash/CA1/_1369_ ),
    .SUM(\hash/CA1/_1370_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3535_  (.A(\hash/d[24] ),
    .B(\hash/h[24] ),
    .CIN(\hash/CA1/_1371_ ),
    .COUT(\hash/CA1/_1372_ ),
    .SUM(\hash/CA1/_1373_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3536_  (.A(\hash/CA1/_1365_ ),
    .B(\hash/CA1/_1374_ ),
    .CIN(\hash/CA1/_1373_ ),
    .COUT(\hash/CA1/_1375_ ),
    .SUM(\hash/CA1/_1376_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3537_  (.A(\hash/d[25] ),
    .B(\hash/h[25] ),
    .CIN(\hash/CA1/_1377_ ),
    .COUT(\hash/CA1/_1378_ ),
    .SUM(\hash/CA1/_1379_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3538_  (.A(\hash/CA1/_1380_ ),
    .B(\hash/CA1/_1381_ ),
    .CIN(\hash/CA1/_1181_ ),
    .COUT(\hash/CA1/_1382_ ),
    .SUM(\hash/CA1/_1383_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3539_  (.A(\hash/d[26] ),
    .B(\hash/h[26] ),
    .CIN(\hash/CA1/_1384_ ),
    .COUT(\hash/CA1/_1385_ ),
    .SUM(\hash/CA1/_1386_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3540_  (.A(\hash/CA1/_1387_ ),
    .B(\hash/CA1/_1386_ ),
    .CIN(\hash/CA1/_1378_ ),
    .COUT(\hash/CA1/_1388_ ),
    .SUM(\hash/CA1/_1389_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3541_  (.A(\hash/CA1/_1390_ ),
    .B(\hash/CA1/_1194_ ),
    .CIN(\hash/CA1/_1195_ ),
    .COUT(\hash/CA1/_1391_ ),
    .SUM(\hash/CA1/_1392_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3542_  (.A(\hash/CA1/_1393_ ),
    .B(\hash/CA1/_1190_ ),
    .CIN(\hash/CA1/_1385_ ),
    .COUT(\hash/CA1/_1394_ ),
    .SUM(\hash/CA1/_1395_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3543_  (.A(\hash/CA1/_1396_ ),
    .B(\hash/CA1/_1201_ ),
    .CIN(\hash/CA1/_1200_ ),
    .COUT(\hash/CA1/_1397_ ),
    .SUM(\hash/CA1/_1398_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3544_  (.A(\hash/CA1/_1196_ ),
    .B(\hash/CA1/_1399_ ),
    .CIN(\hash/CA1/_1400_ ),
    .COUT(\hash/CA1/_1401_ ),
    .SUM(\hash/CA1/_1402_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3545_  (.A(\hash/CA1/_1403_ ),
    .B(\hash/CA1/_1206_ ),
    .CIN(\hash/CA1/_1207_ ),
    .COUT(\hash/CA1/_1404_ ),
    .SUM(\hash/CA1/_1405_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3546_  (.A(\hash/CA1/_1405_ ),
    .B(\hash/CA1/_1397_ ),
    .CIN(\hash/CA1/_1208_ ),
    .COUT(\hash/CA1/_1406_ ),
    .SUM(\hash/CA1/_1407_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3547_  (.A(\hash/d[30] ),
    .B(\hash/h[30] ),
    .CIN(\hash/CA1/_1209_ ),
    .COUT(\hash/CA1/_1408_ ),
    .SUM(\hash/CA1/_1409_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3548_  (.A(\hash/CA1/_1409_ ),
    .B(\hash/CA1/_1410_ ),
    .CIN(\hash/CA1/_1210_ ),
    .COUT(\hash/CA1/_1411_ ),
    .SUM(\hash/CA1/_1412_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3549_  (.A(\hash/CA1/s0[1] ),
    .B(\hash/CA1/_1413_ ),
    .CIN(\hash/CA1/_1414_ ),
    .COUT(\hash/CA1/_1415_ ),
    .SUM(\hash/p1[1] ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3550_  (.A(\hash/CA1/_1416_ ),
    .B(\hash/CA1/_1222_ ),
    .CIN(\hash/CA1/_1417_ ),
    .COUT(\hash/CA1/_1418_ ),
    .SUM(\hash/CA1/_1419_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3551_  (.A(\hash/CA1/_1214_ ),
    .B(\hash/CA1/_1420_ ),
    .CIN(\hash/CA1/_1215_ ),
    .COUT(\hash/CA1/_1421_ ),
    .SUM(\hash/CA1/_1422_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3552_  (.A(\hash/CA1/_1423_ ),
    .B(\hash/CA1/_1424_ ),
    .CIN(\hash/CA1/_1425_ ),
    .COUT(\hash/CA1/_1426_ ),
    .SUM(\hash/CA1/_1427_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA1/_3553_  (.A(\hash/c[1] ),
    .B(\hash/CA1/_1428_ ),
    .CIN(\hash/p4[1] ),
    .COUT(\hash/CA1/_1429_ ),
    .SUM(\hash/p5[1] ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3554_  (.A(\hash/CA1/s0[1] ),
    .B(\hash/CA1/_1413_ ),
    .COUT(\hash/CA1/_1430_ ),
    .SUM(\hash/CA1/_1431_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3555_  (.A(\hash/CA1/s0[2] ),
    .B(\hash/CA1/_1432_ ),
    .COUT(\hash/CA1/_1433_ ),
    .SUM(\hash/CA1/_1434_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3556_  (.A(\hash/CA1/s0[3] ),
    .B(\hash/CA1/_1435_ ),
    .COUT(\hash/CA1/_1436_ ),
    .SUM(\hash/CA1/_1437_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3557_  (.A(\hash/CA1/s0[4] ),
    .B(\hash/CA1/_1438_ ),
    .COUT(\hash/CA1/_1439_ ),
    .SUM(\hash/CA1/_1440_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3558_  (.A(\hash/CA1/s0[5] ),
    .B(\hash/CA1/_1441_ ),
    .COUT(\hash/CA1/_1442_ ),
    .SUM(\hash/CA1/_1443_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3559_  (.A(\hash/CA1/s0[6] ),
    .B(\hash/CA1/_1444_ ),
    .COUT(\hash/CA1/_1445_ ),
    .SUM(\hash/CA1/_1446_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3560_  (.A(\hash/CA1/s0[7] ),
    .B(\hash/CA1/_1447_ ),
    .COUT(\hash/CA1/_1448_ ),
    .SUM(\hash/CA1/_1449_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3561_  (.A(\hash/CA1/s0[8] ),
    .B(\hash/CA1/_1450_ ),
    .COUT(\hash/CA1/_1451_ ),
    .SUM(\hash/CA1/_1452_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3562_  (.A(\hash/CA1/s0[9] ),
    .B(\hash/CA1/_1453_ ),
    .COUT(\hash/CA1/_1454_ ),
    .SUM(\hash/CA1/_1455_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3563_  (.A(\hash/CA1/s0[10] ),
    .B(\hash/CA1/_1456_ ),
    .COUT(\hash/CA1/_1457_ ),
    .SUM(\hash/CA1/_1458_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3564_  (.A(\hash/CA1/s0[11] ),
    .B(\hash/CA1/_1459_ ),
    .COUT(\hash/CA1/_1460_ ),
    .SUM(\hash/CA1/_1461_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3565_  (.A(\hash/CA1/s0[12] ),
    .B(\hash/CA1/_1462_ ),
    .COUT(\hash/CA1/_1463_ ),
    .SUM(\hash/CA1/_1464_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3566_  (.A(\hash/CA1/s0[13] ),
    .B(\hash/CA1/_1465_ ),
    .COUT(\hash/CA1/_1466_ ),
    .SUM(\hash/CA1/_1467_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3567_  (.A(\hash/CA1/s0[14] ),
    .B(\hash/CA1/_1468_ ),
    .COUT(\hash/CA1/_1469_ ),
    .SUM(\hash/CA1/_1470_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3568_  (.A(\hash/CA1/s0[15] ),
    .B(\hash/CA1/_1471_ ),
    .COUT(\hash/CA1/_1472_ ),
    .SUM(\hash/CA1/_1473_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3569_  (.A(\hash/CA1/s0[16] ),
    .B(\hash/CA1/_1474_ ),
    .COUT(\hash/CA1/_1475_ ),
    .SUM(\hash/CA1/_1476_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3570_  (.A(\hash/CA1/s0[17] ),
    .B(\hash/CA1/_1477_ ),
    .COUT(\hash/CA1/_1478_ ),
    .SUM(\hash/CA1/_1479_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3571_  (.A(\hash/CA1/s0[18] ),
    .B(\hash/CA1/_1480_ ),
    .COUT(\hash/CA1/_1481_ ),
    .SUM(\hash/CA1/_1482_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3572_  (.A(\hash/CA1/s0[19] ),
    .B(\hash/CA1/_1483_ ),
    .COUT(\hash/CA1/_1484_ ),
    .SUM(\hash/CA1/_1485_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3573_  (.A(\hash/CA1/s0[20] ),
    .B(\hash/CA1/_1486_ ),
    .COUT(\hash/CA1/_1487_ ),
    .SUM(\hash/CA1/_1488_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3574_  (.A(\hash/CA1/s0[21] ),
    .B(\hash/CA1/_1489_ ),
    .COUT(\hash/CA1/_1490_ ),
    .SUM(\hash/CA1/_1491_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3575_  (.A(\hash/CA1/s0[22] ),
    .B(\hash/CA1/_1492_ ),
    .COUT(\hash/CA1/_1493_ ),
    .SUM(\hash/CA1/_1494_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3576_  (.A(\hash/CA1/s0[23] ),
    .B(\hash/CA1/_1495_ ),
    .COUT(\hash/CA1/_1496_ ),
    .SUM(\hash/CA1/_1497_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3577_  (.A(\hash/CA1/s0[24] ),
    .B(\hash/CA1/_1498_ ),
    .COUT(\hash/CA1/_1499_ ),
    .SUM(\hash/CA1/_1500_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3578_  (.A(\hash/CA1/s0[25] ),
    .B(\hash/CA1/_1501_ ),
    .COUT(\hash/CA1/_1502_ ),
    .SUM(\hash/CA1/_1503_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3579_  (.A(\hash/CA1/s0[26] ),
    .B(\hash/CA1/_1504_ ),
    .COUT(\hash/CA1/_1505_ ),
    .SUM(\hash/CA1/_1506_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3580_  (.A(\hash/CA1/s0[27] ),
    .B(\hash/CA1/_1507_ ),
    .COUT(\hash/CA1/_1508_ ),
    .SUM(\hash/CA1/_1509_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3581_  (.A(\hash/CA1/s0[28] ),
    .B(\hash/CA1/_1510_ ),
    .COUT(\hash/CA1/_1511_ ),
    .SUM(\hash/CA1/_1512_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3582_  (.A(\hash/CA1/s0[29] ),
    .B(\hash/CA1/_1513_ ),
    .COUT(\hash/CA1/_1514_ ),
    .SUM(\hash/CA1/_1515_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3583_  (.A(\hash/CA1/s0[30] ),
    .B(\hash/CA1/_1516_ ),
    .COUT(\hash/CA1/_1517_ ),
    .SUM(\hash/CA1/_1518_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3584_  (.A(\hash/CA1/_0988_ ),
    .B(\hash/CA1/_0990_ ),
    .COUT(\hash/CA1/_1519_ ),
    .SUM(\hash/p4[1] ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3585_  (.A(\hash/CA1/_0989_ ),
    .B(\hash/CA1/_0992_ ),
    .COUT(\hash/CA1/_1520_ ),
    .SUM(\hash/CA1/_1521_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3586_  (.A(\hash/CA1/_0999_ ),
    .B(\hash/CA1/_0991_ ),
    .COUT(\hash/CA1/_1522_ ),
    .SUM(\hash/CA1/_1523_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3587_  (.A(\hash/CA1/_0998_ ),
    .B(\hash/CA1/_1001_ ),
    .COUT(\hash/CA1/_1524_ ),
    .SUM(\hash/CA1/_1525_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3588_  (.A(\hash/CA1/_1003_ ),
    .B(\hash/CA1/_1000_ ),
    .COUT(\hash/CA1/_1526_ ),
    .SUM(\hash/CA1/_1527_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3589_  (.A(\hash/CA1/_1005_ ),
    .B(\hash/CA1/_1002_ ),
    .COUT(\hash/CA1/_1528_ ),
    .SUM(\hash/CA1/_1529_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3590_  (.A(\hash/CA1/_1004_ ),
    .B(\hash/CA1/_1007_ ),
    .COUT(\hash/CA1/_1530_ ),
    .SUM(\hash/CA1/_1531_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3591_  (.A(\hash/CA1/_1006_ ),
    .B(\hash/CA1/_1009_ ),
    .COUT(\hash/CA1/_1532_ ),
    .SUM(\hash/CA1/_1533_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3592_  (.A(\hash/CA1/_1008_ ),
    .B(\hash/CA1/_1011_ ),
    .COUT(\hash/CA1/_1534_ ),
    .SUM(\hash/CA1/_1535_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3593_  (.A(\hash/CA1/_1010_ ),
    .B(\hash/CA1/_1013_ ),
    .COUT(\hash/CA1/_1536_ ),
    .SUM(\hash/CA1/_1537_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3594_  (.A(\hash/CA1/_1012_ ),
    .B(\hash/CA1/_1015_ ),
    .COUT(\hash/CA1/_1538_ ),
    .SUM(\hash/CA1/_1539_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3595_  (.A(\hash/CA1/_1017_ ),
    .B(\hash/CA1/_1014_ ),
    .COUT(\hash/CA1/_1540_ ),
    .SUM(\hash/CA1/_1541_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3596_  (.A(\hash/CA1/_1016_ ),
    .B(\hash/CA1/_1019_ ),
    .COUT(\hash/CA1/_1542_ ),
    .SUM(\hash/CA1/_1543_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3597_  (.A(\hash/CA1/_1021_ ),
    .B(\hash/CA1/_1018_ ),
    .COUT(\hash/CA1/_1544_ ),
    .SUM(\hash/CA1/_1545_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3598_  (.A(\hash/CA1/_1023_ ),
    .B(\hash/CA1/_1020_ ),
    .COUT(\hash/CA1/_1546_ ),
    .SUM(\hash/CA1/_1547_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3599_  (.A(\hash/CA1/_1022_ ),
    .B(\hash/CA1/_1025_ ),
    .COUT(\hash/CA1/_1548_ ),
    .SUM(\hash/CA1/_1549_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3600_  (.A(\hash/CA1/_1024_ ),
    .B(\hash/CA1/_1027_ ),
    .COUT(\hash/CA1/_1550_ ),
    .SUM(\hash/CA1/_1551_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3601_  (.A(\hash/CA1/_1026_ ),
    .B(\hash/CA1/_1029_ ),
    .COUT(\hash/CA1/_1552_ ),
    .SUM(\hash/CA1/_1553_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3602_  (.A(\hash/CA1/_1028_ ),
    .B(\hash/CA1/_1031_ ),
    .COUT(\hash/CA1/_1554_ ),
    .SUM(\hash/CA1/_1555_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3603_  (.A(\hash/CA1/_1030_ ),
    .B(\hash/CA1/_1033_ ),
    .COUT(\hash/CA1/_1556_ ),
    .SUM(\hash/CA1/_1557_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3604_  (.A(\hash/CA1/_1035_ ),
    .B(\hash/CA1/_1032_ ),
    .COUT(\hash/CA1/_1558_ ),
    .SUM(\hash/CA1/_1559_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3605_  (.A(\hash/CA1/_1037_ ),
    .B(\hash/CA1/_1034_ ),
    .COUT(\hash/CA1/_1560_ ),
    .SUM(\hash/CA1/_1561_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3606_  (.A(\hash/CA1/_1039_ ),
    .B(\hash/CA1/_1036_ ),
    .COUT(\hash/CA1/_1562_ ),
    .SUM(\hash/CA1/_1563_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3607_  (.A(\hash/CA1/_1038_ ),
    .B(\hash/CA1/_1041_ ),
    .COUT(\hash/CA1/_1564_ ),
    .SUM(\hash/CA1/_1565_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3608_  (.A(\hash/CA1/_1040_ ),
    .B(\hash/CA1/_1043_ ),
    .COUT(\hash/CA1/_1566_ ),
    .SUM(\hash/CA1/_1567_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3609_  (.A(\hash/CA1/_1045_ ),
    .B(\hash/CA1/_1042_ ),
    .COUT(\hash/CA1/_1568_ ),
    .SUM(\hash/CA1/_1569_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3610_  (.A(\hash/CA1/_1044_ ),
    .B(\hash/CA1/_1047_ ),
    .COUT(\hash/CA1/_1570_ ),
    .SUM(\hash/CA1/_1571_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3611_  (.A(\hash/CA1/_1046_ ),
    .B(\hash/CA1/_1049_ ),
    .COUT(\hash/CA1/_1572_ ),
    .SUM(\hash/CA1/_1573_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3612_  (.A(\hash/CA1/_1048_ ),
    .B(\hash/CA1/_1051_ ),
    .COUT(\hash/CA1/_1574_ ),
    .SUM(\hash/CA1/_1575_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3613_  (.A(\hash/CA1/_1050_ ),
    .B(\hash/CA1/_1053_ ),
    .COUT(\hash/CA1/_1576_ ),
    .SUM(\hash/CA1/_1577_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3614_  (.A(\hash/c[1] ),
    .B(\hash/p4[1] ),
    .COUT(\hash/CA1/_1578_ ),
    .SUM(\hash/CA1/_1579_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3615_  (.A(\hash/c[2] ),
    .B(\hash/p4[2] ),
    .COUT(\hash/CA1/_1580_ ),
    .SUM(\hash/CA1/_1581_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3616_  (.A(\hash/c[3] ),
    .B(\hash/p4[3] ),
    .COUT(\hash/CA1/_1582_ ),
    .SUM(\hash/CA1/_1583_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3617_  (.A(\hash/c[4] ),
    .B(\hash/p4[4] ),
    .COUT(\hash/CA1/_1584_ ),
    .SUM(\hash/CA1/_1585_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3618_  (.A(\hash/c[5] ),
    .B(\hash/p4[5] ),
    .COUT(\hash/CA1/_1586_ ),
    .SUM(\hash/CA1/_1587_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3619_  (.A(\hash/c[6] ),
    .B(\hash/p4[6] ),
    .COUT(\hash/CA1/_1588_ ),
    .SUM(\hash/CA1/_1589_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3620_  (.A(\hash/c[7] ),
    .B(\hash/p4[7] ),
    .COUT(\hash/CA1/_1590_ ),
    .SUM(\hash/CA1/_1591_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3621_  (.A(\hash/c[8] ),
    .B(\hash/p4[8] ),
    .COUT(\hash/CA1/_1592_ ),
    .SUM(\hash/CA1/_1593_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3622_  (.A(\hash/c[9] ),
    .B(\hash/p4[9] ),
    .COUT(\hash/CA1/_1594_ ),
    .SUM(\hash/CA1/_1595_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3623_  (.A(\hash/c[10] ),
    .B(\hash/p4[10] ),
    .COUT(\hash/CA1/_1596_ ),
    .SUM(\hash/CA1/_1597_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3624_  (.A(\hash/c[11] ),
    .B(\hash/p4[11] ),
    .COUT(\hash/CA1/_1598_ ),
    .SUM(\hash/CA1/_1599_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3625_  (.A(\hash/c[12] ),
    .B(\hash/p4[12] ),
    .COUT(\hash/CA1/_1600_ ),
    .SUM(\hash/CA1/_1601_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3626_  (.A(\hash/c[13] ),
    .B(\hash/p4[13] ),
    .COUT(\hash/CA1/_1602_ ),
    .SUM(\hash/CA1/_1603_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3627_  (.A(\hash/c[14] ),
    .B(\hash/p4[14] ),
    .COUT(\hash/CA1/_1604_ ),
    .SUM(\hash/CA1/_1605_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3628_  (.A(\hash/c[15] ),
    .B(\hash/p4[15] ),
    .COUT(\hash/CA1/_1606_ ),
    .SUM(\hash/CA1/_1607_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3629_  (.A(\hash/c[16] ),
    .B(\hash/p4[16] ),
    .COUT(\hash/CA1/_1608_ ),
    .SUM(\hash/CA1/_1609_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3630_  (.A(\hash/c[17] ),
    .B(\hash/p4[17] ),
    .COUT(\hash/CA1/_1610_ ),
    .SUM(\hash/CA1/_1611_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3631_  (.A(\hash/c[18] ),
    .B(\hash/p4[18] ),
    .COUT(\hash/CA1/_1612_ ),
    .SUM(\hash/CA1/_1613_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3632_  (.A(\hash/c[19] ),
    .B(\hash/p4[19] ),
    .COUT(\hash/CA1/_1614_ ),
    .SUM(\hash/CA1/_1615_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3633_  (.A(\hash/c[20] ),
    .B(\hash/p4[20] ),
    .COUT(\hash/CA1/_1616_ ),
    .SUM(\hash/CA1/_1617_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3634_  (.A(\hash/c[21] ),
    .B(\hash/p4[21] ),
    .COUT(\hash/CA1/_1618_ ),
    .SUM(\hash/CA1/_1619_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3635_  (.A(\hash/c[22] ),
    .B(\hash/p4[22] ),
    .COUT(\hash/CA1/_1620_ ),
    .SUM(\hash/CA1/_1621_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3636_  (.A(\hash/c[23] ),
    .B(\hash/p4[23] ),
    .COUT(\hash/CA1/_1622_ ),
    .SUM(\hash/CA1/_1623_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3637_  (.A(\hash/c[24] ),
    .B(\hash/p4[24] ),
    .COUT(\hash/CA1/_1624_ ),
    .SUM(\hash/CA1/_1625_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3638_  (.A(\hash/c[25] ),
    .B(\hash/p4[25] ),
    .COUT(\hash/CA1/_1626_ ),
    .SUM(\hash/CA1/_1627_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3639_  (.A(\hash/c[26] ),
    .B(\hash/p4[26] ),
    .COUT(\hash/CA1/_1628_ ),
    .SUM(\hash/CA1/_1629_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3640_  (.A(\hash/c[27] ),
    .B(\hash/p4[27] ),
    .COUT(\hash/CA1/_1630_ ),
    .SUM(\hash/CA1/_1631_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3641_  (.A(\hash/c[28] ),
    .B(\hash/p4[28] ),
    .COUT(\hash/CA1/_1632_ ),
    .SUM(\hash/CA1/_1633_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3642_  (.A(\hash/c[29] ),
    .B(\hash/p4[29] ),
    .COUT(\hash/CA1/_1634_ ),
    .SUM(\hash/CA1/_1635_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3643_  (.A(\hash/c[30] ),
    .B(\hash/p4[30] ),
    .COUT(\hash/CA1/_1636_ ),
    .SUM(\hash/CA1/_1637_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3644_  (.A(\k_value1[0] ),
    .B(\w_value1[0] ),
    .COUT(\hash/CA1/_1638_ ),
    .SUM(\hash/CA1/_1639_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3645_  (.A(\hash/CA1/s1[0] ),
    .B(\hash/CA1/_1640_ ),
    .COUT(\hash/CA1/_1641_ ),
    .SUM(\hash/CA1/_1642_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3646_  (.A(\k_value1[1] ),
    .B(\w_value1[1] ),
    .COUT(\hash/CA1/_1643_ ),
    .SUM(\hash/CA1/_1644_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3647_  (.A(\hash/CA1/s1[1] ),
    .B(\hash/CA1/_1645_ ),
    .COUT(\hash/CA1/_1646_ ),
    .SUM(\hash/CA1/_1647_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3648_  (.A(\k_value1[2] ),
    .B(\w_value1[2] ),
    .COUT(\hash/CA1/_1648_ ),
    .SUM(\hash/CA1/_1649_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3649_  (.A(\hash/CA1/s1[2] ),
    .B(\hash/CA1/_1650_ ),
    .COUT(\hash/CA1/_1651_ ),
    .SUM(\hash/CA1/_1652_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3650_  (.A(\hash/CA1/_1071_ ),
    .B(\hash/CA1/_1066_ ),
    .COUT(\hash/CA1/_1653_ ),
    .SUM(\hash/CA1/_1654_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3651_  (.A(\k_value1[3] ),
    .B(\w_value1[3] ),
    .COUT(\hash/CA1/_1655_ ),
    .SUM(\hash/CA1/_1656_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3652_  (.A(\hash/CA1/s1[3] ),
    .B(\hash/CA1/_1657_ ),
    .COUT(\hash/CA1/_1658_ ),
    .SUM(\hash/CA1/_1659_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3653_  (.A(\hash/CA1/_1070_ ),
    .B(\hash/CA1/_1075_ ),
    .COUT(\hash/CA1/_1660_ ),
    .SUM(\hash/CA1/_1661_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3654_  (.A(\k_value1[4] ),
    .B(\w_value1[4] ),
    .COUT(\hash/CA1/_1662_ ),
    .SUM(\hash/CA1/_1663_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3655_  (.A(\hash/CA1/s1[4] ),
    .B(\hash/CA1/_1664_ ),
    .COUT(\hash/CA1/_1665_ ),
    .SUM(\hash/CA1/_1666_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3656_  (.A(\hash/CA1/_1667_ ),
    .B(\hash/CA1/_1074_ ),
    .COUT(\hash/CA1/_1668_ ),
    .SUM(\hash/CA1/_1669_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3657_  (.A(\k_value1[5] ),
    .B(\w_value1[5] ),
    .COUT(\hash/CA1/_1670_ ),
    .SUM(\hash/CA1/_1671_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3658_  (.A(\hash/CA1/s1[5] ),
    .B(\hash/CA1/_1672_ ),
    .COUT(\hash/CA1/_1673_ ),
    .SUM(\hash/CA1/_1674_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3659_  (.A(\hash/CA1/_1084_ ),
    .B(\hash/CA1/_1675_ ),
    .COUT(\hash/CA1/_1676_ ),
    .SUM(\hash/CA1/_1677_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3660_  (.A(\k_value1[6] ),
    .B(\w_value1[6] ),
    .COUT(\hash/CA1/_1678_ ),
    .SUM(\hash/CA1/_1679_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3661_  (.A(\hash/CA1/s1[6] ),
    .B(\hash/CA1/_1680_ ),
    .COUT(\hash/CA1/_1681_ ),
    .SUM(\hash/CA1/_1682_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3662_  (.A(\hash/CA1/_1083_ ),
    .B(\hash/CA1/_1088_ ),
    .COUT(\hash/CA1/_1683_ ),
    .SUM(\hash/CA1/_1684_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3663_  (.A(\k_value1[7] ),
    .B(\w_value1[7] ),
    .COUT(\hash/CA1/_1685_ ),
    .SUM(\hash/CA1/_1686_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3664_  (.A(\hash/CA1/s1[7] ),
    .B(\hash/CA1/_1687_ ),
    .COUT(\hash/CA1/_1688_ ),
    .SUM(\hash/CA1/_1689_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3665_  (.A(\hash/CA1/_1087_ ),
    .B(\hash/CA1/_1092_ ),
    .COUT(\hash/CA1/_1690_ ),
    .SUM(\hash/CA1/_1691_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3666_  (.A(\k_value1[8] ),
    .B(\w_value1[8] ),
    .COUT(\hash/CA1/_1692_ ),
    .SUM(\hash/CA1/_1693_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3667_  (.A(\hash/CA1/s1[8] ),
    .B(\hash/CA1/_1694_ ),
    .COUT(\hash/CA1/_1695_ ),
    .SUM(\hash/CA1/_1696_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3668_  (.A(\hash/CA1/_1091_ ),
    .B(\hash/CA1/_1096_ ),
    .COUT(\hash/CA1/_1697_ ),
    .SUM(\hash/CA1/_1698_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3669_  (.A(\k_value1[9] ),
    .B(\w_value1[9] ),
    .COUT(\hash/CA1/_1699_ ),
    .SUM(\hash/CA1/_1700_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3670_  (.A(\hash/CA1/s1[9] ),
    .B(\hash/CA1/_1701_ ),
    .COUT(\hash/CA1/_1702_ ),
    .SUM(\hash/CA1/_1703_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3671_  (.A(\hash/CA1/_1095_ ),
    .B(\hash/CA1/_1704_ ),
    .COUT(\hash/CA1/_1705_ ),
    .SUM(\hash/CA1/_1706_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3672_  (.A(\k_value1[10] ),
    .B(\w_value1[10] ),
    .COUT(\hash/CA1/_1707_ ),
    .SUM(\hash/CA1/_1708_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3673_  (.A(\hash/CA1/s1[10] ),
    .B(\hash/CA1/_1709_ ),
    .COUT(\hash/CA1/_1710_ ),
    .SUM(\hash/CA1/_1711_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3674_  (.A(\hash/CA1/_1712_ ),
    .B(\hash/CA1/_1713_ ),
    .COUT(\hash/CA1/_1714_ ),
    .SUM(\hash/CA1/_1715_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3675_  (.A(\k_value1[11] ),
    .B(\w_value1[11] ),
    .COUT(\hash/CA1/_1716_ ),
    .SUM(\hash/CA1/_1717_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3676_  (.A(\hash/CA1/s1[11] ),
    .B(\hash/CA1/_1718_ ),
    .COUT(\hash/CA1/_1719_ ),
    .SUM(\hash/CA1/_1720_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3677_  (.A(\hash/CA1/_1721_ ),
    .B(\hash/CA1/_1722_ ),
    .COUT(\hash/CA1/_1723_ ),
    .SUM(\hash/CA1/_1724_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3678_  (.A(\k_value1[12] ),
    .B(\w_value1[12] ),
    .COUT(\hash/CA1/_1725_ ),
    .SUM(\hash/CA1/_1726_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3679_  (.A(\hash/CA1/s1[12] ),
    .B(\hash/CA1/_1727_ ),
    .COUT(\hash/CA1/_1728_ ),
    .SUM(\hash/CA1/_1729_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3680_  (.A(\hash/CA1/_1730_ ),
    .B(\hash/CA1/_1731_ ),
    .COUT(\hash/CA1/_1732_ ),
    .SUM(\hash/CA1/_1733_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3681_  (.A(\k_value1[13] ),
    .B(\w_value1[13] ),
    .COUT(\hash/CA1/_1734_ ),
    .SUM(\hash/CA1/_1735_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3682_  (.A(\hash/CA1/s1[13] ),
    .B(\hash/CA1/_1736_ ),
    .COUT(\hash/CA1/_1737_ ),
    .SUM(\hash/CA1/_1738_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3683_  (.A(\hash/CA1/_1739_ ),
    .B(\hash/CA1/_1740_ ),
    .COUT(\hash/CA1/_1741_ ),
    .SUM(\hash/CA1/_1742_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3684_  (.A(\k_value1[14] ),
    .B(\w_value1[14] ),
    .COUT(\hash/CA1/_1743_ ),
    .SUM(\hash/CA1/_1744_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3685_  (.A(\hash/CA1/s1[14] ),
    .B(\hash/CA1/_1745_ ),
    .COUT(\hash/CA1/_1746_ ),
    .SUM(\hash/CA1/_1747_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3686_  (.A(\hash/CA1/_1748_ ),
    .B(\hash/CA1/_1749_ ),
    .COUT(\hash/CA1/_1750_ ),
    .SUM(\hash/CA1/_1751_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3687_  (.A(\k_value1[15] ),
    .B(\w_value1[15] ),
    .COUT(\hash/CA1/_1752_ ),
    .SUM(\hash/CA1/_1753_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3688_  (.A(\hash/CA1/s1[15] ),
    .B(\hash/CA1/_1754_ ),
    .COUT(\hash/CA1/_1755_ ),
    .SUM(\hash/CA1/_1756_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3689_  (.A(\hash/CA1/_1757_ ),
    .B(\hash/CA1/_1132_ ),
    .COUT(\hash/CA1/_1758_ ),
    .SUM(\hash/CA1/_1759_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3690_  (.A(\k_value1[16] ),
    .B(\w_value1[16] ),
    .COUT(\hash/CA1/_1760_ ),
    .SUM(\hash/CA1/_1761_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3691_  (.A(\hash/CA1/s1[16] ),
    .B(\hash/CA1/_1762_ ),
    .COUT(\hash/CA1/_1763_ ),
    .SUM(\hash/CA1/_1764_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3692_  (.A(\hash/CA1/_1131_ ),
    .B(\hash/CA1/_1765_ ),
    .COUT(\hash/CA1/_1766_ ),
    .SUM(\hash/CA1/_1767_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3693_  (.A(\k_value1[17] ),
    .B(\w_value1[17] ),
    .COUT(\hash/CA1/_1768_ ),
    .SUM(\hash/CA1/_1769_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3694_  (.A(\hash/CA1/s1[17] ),
    .B(\hash/CA1/_1770_ ),
    .COUT(\hash/CA1/_1771_ ),
    .SUM(\hash/CA1/_1772_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3695_  (.A(\hash/CA1/_1773_ ),
    .B(\hash/CA1/_1774_ ),
    .COUT(\hash/CA1/_1775_ ),
    .SUM(\hash/CA1/_1776_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3696_  (.A(\k_value1[18] ),
    .B(\w_value1[18] ),
    .COUT(\hash/CA1/_1777_ ),
    .SUM(\hash/CA1/_1778_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3697_  (.A(\hash/CA1/s1[18] ),
    .B(\hash/CA1/_1779_ ),
    .COUT(\hash/CA1/_1780_ ),
    .SUM(\hash/CA1/_1781_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3698_  (.A(\hash/CA1/_1782_ ),
    .B(\hash/CA1/_1783_ ),
    .COUT(\hash/CA1/_1784_ ),
    .SUM(\hash/CA1/_1785_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3699_  (.A(\k_value1[19] ),
    .B(\w_value1[19] ),
    .COUT(\hash/CA1/_1786_ ),
    .SUM(\hash/CA1/_1787_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3700_  (.A(\hash/CA1/s1[19] ),
    .B(\hash/CA1/_1788_ ),
    .COUT(\hash/CA1/_1789_ ),
    .SUM(\hash/CA1/_1790_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3701_  (.A(\hash/CA1/_1791_ ),
    .B(\hash/CA1/_1792_ ),
    .COUT(\hash/CA1/_1793_ ),
    .SUM(\hash/CA1/_1794_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3702_  (.A(\k_value1[20] ),
    .B(\w_value1[20] ),
    .COUT(\hash/CA1/_1795_ ),
    .SUM(\hash/CA1/_1796_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3703_  (.A(\hash/CA1/s1[20] ),
    .B(\hash/CA1/_1797_ ),
    .COUT(\hash/CA1/_1798_ ),
    .SUM(\hash/CA1/_1799_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3704_  (.A(\hash/CA1/_1800_ ),
    .B(\hash/CA1/_1801_ ),
    .COUT(\hash/CA1/_1802_ ),
    .SUM(\hash/CA1/_1803_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3705_  (.A(\k_value1[21] ),
    .B(\w_value1[21] ),
    .COUT(\hash/CA1/_1804_ ),
    .SUM(\hash/CA1/_1805_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3706_  (.A(\hash/CA1/s1[21] ),
    .B(\hash/CA1/_1806_ ),
    .COUT(\hash/CA1/_1807_ ),
    .SUM(\hash/CA1/_1808_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3707_  (.A(\hash/CA1/_1809_ ),
    .B(\hash/CA1/_1810_ ),
    .COUT(\hash/CA1/_1811_ ),
    .SUM(\hash/CA1/_1812_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3708_  (.A(\k_value1[22] ),
    .B(\w_value1[22] ),
    .COUT(\hash/CA1/_1813_ ),
    .SUM(\hash/CA1/_1814_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3709_  (.A(\hash/CA1/s1[22] ),
    .B(\hash/CA1/_1815_ ),
    .COUT(\hash/CA1/_1816_ ),
    .SUM(\hash/CA1/_1817_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3710_  (.A(\hash/CA1/_1818_ ),
    .B(\hash/CA1/_1819_ ),
    .COUT(\hash/CA1/_1820_ ),
    .SUM(\hash/CA1/_1821_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3711_  (.A(\k_value1[23] ),
    .B(\w_value1[23] ),
    .COUT(\hash/CA1/_1822_ ),
    .SUM(\hash/CA1/_1823_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3712_  (.A(\hash/CA1/s1[23] ),
    .B(\hash/CA1/_1824_ ),
    .COUT(\hash/CA1/_1825_ ),
    .SUM(\hash/CA1/_1826_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3713_  (.A(\hash/CA1/_1827_ ),
    .B(\hash/CA1/_1828_ ),
    .COUT(\hash/CA1/_1829_ ),
    .SUM(\hash/CA1/_1830_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3714_  (.A(\k_value1[24] ),
    .B(\w_value1[24] ),
    .COUT(\hash/CA1/_1831_ ),
    .SUM(\hash/CA1/_1832_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3715_  (.A(\hash/CA1/s1[24] ),
    .B(\hash/CA1/_1833_ ),
    .COUT(\hash/CA1/_1834_ ),
    .SUM(\hash/CA1/_1835_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3716_  (.A(\hash/CA1/_1836_ ),
    .B(\hash/CA1/_1837_ ),
    .COUT(\hash/CA1/_1838_ ),
    .SUM(\hash/CA1/_1839_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3717_  (.A(\k_value1[25] ),
    .B(\w_value1[25] ),
    .COUT(\hash/CA1/_1840_ ),
    .SUM(\hash/CA1/_1841_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3718_  (.A(\hash/CA1/s1[25] ),
    .B(\hash/CA1/_1842_ ),
    .COUT(\hash/CA1/_1843_ ),
    .SUM(\hash/CA1/_1844_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3719_  (.A(\hash/CA1/_1845_ ),
    .B(\hash/CA1/_1846_ ),
    .COUT(\hash/CA1/_1847_ ),
    .SUM(\hash/CA1/_1848_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3720_  (.A(\k_value1[26] ),
    .B(\w_value1[26] ),
    .COUT(\hash/CA1/_1849_ ),
    .SUM(\hash/CA1/_1850_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3721_  (.A(\hash/CA1/s1[26] ),
    .B(\hash/CA1/_1851_ ),
    .COUT(\hash/CA1/_1852_ ),
    .SUM(\hash/CA1/_1853_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3722_  (.A(\hash/CA1/_1854_ ),
    .B(\hash/CA1/_1855_ ),
    .COUT(\hash/CA1/_1856_ ),
    .SUM(\hash/CA1/_1857_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3723_  (.A(\k_value1[27] ),
    .B(\w_value1[27] ),
    .COUT(\hash/CA1/_1858_ ),
    .SUM(\hash/CA1/_1859_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3724_  (.A(\hash/CA1/s1[27] ),
    .B(\hash/CA1/_1860_ ),
    .COUT(\hash/CA1/_1861_ ),
    .SUM(\hash/CA1/_1862_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3725_  (.A(\hash/CA1/_1863_ ),
    .B(\hash/CA1/_1193_ ),
    .COUT(\hash/CA1/_1864_ ),
    .SUM(\hash/CA1/_1865_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3726_  (.A(\k_value1[28] ),
    .B(\w_value1[28] ),
    .COUT(\hash/CA1/_1866_ ),
    .SUM(\hash/CA1/_1867_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3727_  (.A(\hash/CA1/s1[28] ),
    .B(\hash/CA1/_1868_ ),
    .COUT(\hash/CA1/_1869_ ),
    .SUM(\hash/CA1/_1870_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3728_  (.A(\hash/CA1/_1192_ ),
    .B(\hash/CA1/_1199_ ),
    .COUT(\hash/CA1/_1871_ ),
    .SUM(\hash/CA1/_1872_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3729_  (.A(\k_value1[29] ),
    .B(\w_value1[29] ),
    .COUT(\hash/CA1/_1873_ ),
    .SUM(\hash/CA1/_1874_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3730_  (.A(\hash/CA1/s1[29] ),
    .B(\hash/CA1/_1875_ ),
    .COUT(\hash/CA1/_1876_ ),
    .SUM(\hash/CA1/_1877_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3731_  (.A(\hash/CA1/_1198_ ),
    .B(\hash/CA1/_1205_ ),
    .COUT(\hash/CA1/_1878_ ),
    .SUM(\hash/CA1/_1879_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3732_  (.A(\k_value1[30] ),
    .B(\w_value1[30] ),
    .COUT(\hash/CA1/_1880_ ),
    .SUM(\hash/CA1/_1881_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3733_  (.A(\hash/CA1/s1[30] ),
    .B(\hash/CA1/_1882_ ),
    .COUT(\hash/CA1/_1883_ ),
    .SUM(\hash/CA1/_1884_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3734_  (.A(\hash/CA1/_1212_ ),
    .B(\hash/CA1/_1204_ ),
    .COUT(\hash/CA1/_1885_ ),
    .SUM(\hash/CA1/_1886_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3735_  (.A(\hash/CA1/_1232_ ),
    .B(\hash/CA1/_1887_ ),
    .COUT(\hash/CA1/_1888_ ),
    .SUM(\hash/CA1/_1889_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3736_  (.A(\hash/CA1/_1231_ ),
    .B(\hash/CA1/_1241_ ),
    .COUT(\hash/CA1/_1890_ ),
    .SUM(\hash/CA1/_1891_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3737_  (.A(\hash/CA1/_1248_ ),
    .B(\hash/CA1/_1240_ ),
    .COUT(\hash/CA1/_1892_ ),
    .SUM(\hash/CA1/_1893_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3738_  (.A(\hash/CA1/_1247_ ),
    .B(\hash/CA1/_1894_ ),
    .COUT(\hash/CA1/_1895_ ),
    .SUM(\hash/CA1/_1896_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3739_  (.A(\hash/CA1/_1897_ ),
    .B(\hash/CA1/_1898_ ),
    .COUT(\hash/CA1/_1899_ ),
    .SUM(\hash/CA1/_1900_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3740_  (.A(\hash/CA1/_1901_ ),
    .B(\hash/CA1/_1902_ ),
    .COUT(\hash/CA1/_1903_ ),
    .SUM(\hash/CA1/_1904_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3741_  (.A(\hash/CA1/_1275_ ),
    .B(\hash/CA1/_1905_ ),
    .COUT(\hash/CA1/_1906_ ),
    .SUM(\hash/CA1/_1907_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3742_  (.A(\hash/CA1/_1274_ ),
    .B(\hash/CA1/_1908_ ),
    .COUT(\hash/CA1/_1909_ ),
    .SUM(\hash/CA1/_1910_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3743_  (.A(\hash/CA1/_1911_ ),
    .B(\hash/CA1/_1912_ ),
    .COUT(\hash/CA1/_1913_ ),
    .SUM(\hash/CA1/_1914_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3744_  (.A(\hash/CA1/_1915_ ),
    .B(\hash/CA1/_1916_ ),
    .COUT(\hash/CA1/_1917_ ),
    .SUM(\hash/CA1/_1918_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3745_  (.A(\hash/CA1/_1919_ ),
    .B(\hash/CA1/_1920_ ),
    .COUT(\hash/CA1/_1921_ ),
    .SUM(\hash/CA1/_1922_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3746_  (.A(\hash/CA1/_1923_ ),
    .B(\hash/CA1/_1308_ ),
    .COUT(\hash/CA1/_1924_ ),
    .SUM(\hash/CA1/_1925_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3747_  (.A(\hash/CA1/_1307_ ),
    .B(\hash/CA1/_1314_ ),
    .COUT(\hash/CA1/_1926_ ),
    .SUM(\hash/CA1/_1927_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3748_  (.A(\hash/CA1/_1313_ ),
    .B(\hash/CA1/_1320_ ),
    .COUT(\hash/CA1/_1928_ ),
    .SUM(\hash/CA1/_1929_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3749_  (.A(\hash/CA1/_1930_ ),
    .B(\hash/CA1/_1319_ ),
    .COUT(\hash/CA1/_1931_ ),
    .SUM(\hash/CA1/_1932_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3750_  (.A(\hash/CA1/_1332_ ),
    .B(\hash/CA1/_1933_ ),
    .COUT(\hash/CA1/_1934_ ),
    .SUM(\hash/CA1/_1935_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3751_  (.A(\hash/CA1/_1331_ ),
    .B(\hash/CA1/_1338_ ),
    .COUT(\hash/CA1/_1936_ ),
    .SUM(\hash/CA1/_1937_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3752_  (.A(\hash/CA1/_1337_ ),
    .B(\hash/CA1/_1344_ ),
    .COUT(\hash/CA1/_1938_ ),
    .SUM(\hash/CA1/_1939_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3753_  (.A(\hash/CA1/_1343_ ),
    .B(\hash/CA1/_1940_ ),
    .COUT(\hash/CA1/_1941_ ),
    .SUM(\hash/CA1/_1942_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3754_  (.A(\hash/CA1/_1943_ ),
    .B(\hash/CA1/_1357_ ),
    .COUT(\hash/CA1/_1944_ ),
    .SUM(\hash/CA1/_1945_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3755_  (.A(\hash/CA1/_1363_ ),
    .B(\hash/CA1/_1356_ ),
    .COUT(\hash/CA1/_1946_ ),
    .SUM(\hash/CA1/_1947_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3756_  (.A(\hash/CA1/_1948_ ),
    .B(\hash/CA1/_1362_ ),
    .COUT(\hash/CA1/_1949_ ),
    .SUM(\hash/CA1/_1950_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3757_  (.A(\hash/CA1/_1376_ ),
    .B(\hash/CA1/_1951_ ),
    .COUT(\hash/CA1/_1952_ ),
    .SUM(\hash/CA1/_1953_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3758_  (.A(\hash/CA1/_1375_ ),
    .B(\hash/CA1/_1954_ ),
    .COUT(\hash/CA1/_1955_ ),
    .SUM(\hash/CA1/_1956_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3759_  (.A(\hash/CA1/_1389_ ),
    .B(\hash/CA1/_1957_ ),
    .COUT(\hash/CA1/_1958_ ),
    .SUM(\hash/CA1/_1959_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3760_  (.A(\hash/CA1/_1388_ ),
    .B(\hash/CA1/_1395_ ),
    .COUT(\hash/CA1/_1960_ ),
    .SUM(\hash/CA1/_1961_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3761_  (.A(\hash/CA1/_1402_ ),
    .B(\hash/CA1/_1394_ ),
    .COUT(\hash/CA1/_1962_ ),
    .SUM(\hash/CA1/_1963_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3762_  (.A(\hash/CA1/_1964_ ),
    .B(\hash/CA1/_1401_ ),
    .COUT(\hash/CA1/_1965_ ),
    .SUM(\hash/CA1/_1966_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3763_  (.A(\hash/CA1/_1412_ ),
    .B(\hash/CA1/_1967_ ),
    .COUT(\hash/CA1/_1968_ ),
    .SUM(\hash/CA1/_1969_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3764_  (.A(\hash/CA1/s0[0] ),
    .B(\hash/CA1/_1970_ ),
    .COUT(\hash/CA1/_1414_ ),
    .SUM(\hash/p1[0] ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3765_  (.A(\hash/CA1/_1642_ ),
    .B(\hash/CA1/_1971_ ),
    .COUT(\hash/CA1/_1972_ ),
    .SUM(\hash/p2[0] ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3766_  (.A(\hash/CA1/_1973_ ),
    .B(\hash/CA1/_1972_ ),
    .COUT(\hash/CA1/_1974_ ),
    .SUM(\hash/p2[1] ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3767_  (.A(\hash/CA1/_1975_ ),
    .B(\hash/CA1/_1067_ ),
    .COUT(\hash/CA1/_1976_ ),
    .SUM(\hash/p3[1] ));
 sky130_fd_sc_hd__ha_1 \hash/CA1/_3768_  (.A(\hash/c[0] ),
    .B(\hash/p4[0] ),
    .COUT(\hash/CA1/_1428_ ),
    .SUM(\hash/p5[0] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_00_  (.A(\hash/b_new[13] ),
    .B(\hash/b_new[2] ),
    .C(\hash/b_new[22] ),
    .X(\hash/CA2/s0[0] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_01_  (.A(\hash/b_new[23] ),
    .B(\hash/b_new[12] ),
    .C(\hash/b_new[0] ),
    .X(\hash/CA2/s0[10] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_02_  (.A(\hash/b_new[13] ),
    .B(\hash/b_new[24] ),
    .C(\hash/b_new[1] ),
    .X(\hash/CA2/s0[11] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_03_  (.A(\hash/b_new[2] ),
    .B(\hash/b_new[14] ),
    .C(\hash/b_new[25] ),
    .X(\hash/CA2/s0[12] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_04_  (.A(\hash/b_new[3] ),
    .B(\hash/b_new[15] ),
    .C(\hash/b_new[26] ),
    .X(\hash/CA2/s0[13] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_05_  (.A(\hash/b_new[4] ),
    .B(\hash/b_new[16] ),
    .C(\hash/b_new[27] ),
    .X(\hash/CA2/s0[14] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_06_  (.A(\hash/b_new[5] ),
    .B(\hash/b_new[17] ),
    .C(\hash/b_new[28] ),
    .X(\hash/CA2/s0[15] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_07_  (.A(\hash/b_new[6] ),
    .B(\hash/b_new[18] ),
    .C(\hash/b_new[29] ),
    .X(\hash/CA2/s0[16] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_08_  (.A(\hash/b_new[7] ),
    .B(\hash/b_new[19] ),
    .C(\hash/b_new[30] ),
    .X(\hash/CA2/s0[17] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_09_  (.A(\hash/b_new[8] ),
    .B(\hash/b_new[20] ),
    .C(\hash/b_new[31] ),
    .X(\hash/CA2/s0[18] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_10_  (.A(\hash/b_new[9] ),
    .B(\hash/b_new[21] ),
    .C(\hash/b_new[0] ),
    .X(\hash/CA2/s0[19] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_11_  (.A(\hash/b_new[14] ),
    .B(\hash/b_new[3] ),
    .C(\hash/b_new[23] ),
    .X(\hash/CA2/s0[1] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_12_  (.A(\hash/b_new[10] ),
    .B(\hash/b_new[22] ),
    .C(\hash/b_new[1] ),
    .X(\hash/CA2/s0[20] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_13_  (.A(\hash/b_new[2] ),
    .B(\hash/b_new[11] ),
    .C(\hash/b_new[23] ),
    .X(\hash/CA2/s0[21] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_14_  (.A(\hash/b_new[3] ),
    .B(\hash/b_new[12] ),
    .C(\hash/b_new[24] ),
    .X(\hash/CA2/s0[22] ));
 sky130_fd_sc_hd__xor3_4 \hash/CA2/S0/_15_  (.A(\hash/b_new[13] ),
    .B(\hash/b_new[4] ),
    .C(\hash/b_new[25] ),
    .X(\hash/CA2/s0[23] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_16_  (.A(\hash/b_new[14] ),
    .B(\hash/b_new[5] ),
    .C(\hash/b_new[26] ),
    .X(\hash/CA2/s0[24] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_17_  (.A(\hash/b_new[15] ),
    .B(\hash/b_new[6] ),
    .C(\hash/b_new[27] ),
    .X(\hash/CA2/s0[25] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_18_  (.A(\hash/b_new[16] ),
    .B(\hash/b_new[7] ),
    .C(\hash/b_new[28] ),
    .X(\hash/CA2/s0[26] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_19_  (.A(\hash/b_new[17] ),
    .B(\hash/b_new[8] ),
    .C(\hash/b_new[29] ),
    .X(\hash/CA2/s0[27] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_20_  (.A(\hash/b_new[18] ),
    .B(\hash/b_new[9] ),
    .C(\hash/b_new[30] ),
    .X(\hash/CA2/s0[28] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_21_  (.A(\hash/b_new[19] ),
    .B(\hash/b_new[10] ),
    .C(\hash/b_new[31] ),
    .X(\hash/CA2/s0[29] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_22_  (.A(\hash/b_new[15] ),
    .B(\hash/b_new[4] ),
    .C(\hash/b_new[24] ),
    .X(\hash/CA2/s0[2] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_23_  (.A(\hash/b_new[20] ),
    .B(\hash/b_new[11] ),
    .C(\hash/b_new[0] ),
    .X(\hash/CA2/s0[30] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_24_  (.A(\hash/b_new[21] ),
    .B(\hash/b_new[12] ),
    .C(\hash/b_new[1] ),
    .X(\hash/CA2/s0[31] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_25_  (.A(\hash/b_new[16] ),
    .B(\hash/b_new[5] ),
    .C(\hash/b_new[25] ),
    .X(\hash/CA2/s0[3] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_26_  (.A(\hash/b_new[17] ),
    .B(\hash/b_new[6] ),
    .C(\hash/b_new[26] ),
    .X(\hash/CA2/s0[4] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_27_  (.A(\hash/b_new[18] ),
    .B(\hash/b_new[7] ),
    .C(\hash/b_new[27] ),
    .X(\hash/CA2/s0[5] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_28_  (.A(\hash/b_new[19] ),
    .B(\hash/b_new[8] ),
    .C(\hash/b_new[28] ),
    .X(\hash/CA2/s0[6] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_29_  (.A(\hash/b_new[20] ),
    .B(\hash/b_new[9] ),
    .C(\hash/b_new[29] ),
    .X(\hash/CA2/s0[7] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_30_  (.A(\hash/b_new[21] ),
    .B(\hash/b_new[10] ),
    .C(\hash/b_new[30] ),
    .X(\hash/CA2/s0[8] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S0/_31_  (.A(\hash/b_new[22] ),
    .B(\hash/b_new[11] ),
    .C(\hash/b_new[31] ),
    .X(\hash/CA2/s0[9] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_00_  (.A(\hash/p2_cap[11] ),
    .B(\hash/p2_cap[6] ),
    .C(\hash/p2_cap[25] ),
    .X(\hash/CA2/s1[0] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_01_  (.A(\hash/p2_cap[16] ),
    .B(\hash/p2_cap[21] ),
    .C(\hash/p2_cap[3] ),
    .X(\hash/CA2/s1[10] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_02_  (.A(\hash/p2_cap[17] ),
    .B(\hash/p2_cap[22] ),
    .C(\hash/p2_cap[4] ),
    .X(\hash/CA2/s1[11] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_03_  (.A(\hash/p2_cap[18] ),
    .B(\hash/p2_cap[23] ),
    .C(\hash/p2_cap[5] ),
    .X(\hash/CA2/s1[12] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_04_  (.A(\hash/p2_cap[6] ),
    .B(\hash/p2_cap[19] ),
    .C(\hash/p2_cap[24] ),
    .X(\hash/CA2/s1[13] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_05_  (.A(\hash/p2_cap[7] ),
    .B(\hash/p2_cap[20] ),
    .C(\hash/p2_cap[25] ),
    .X(\hash/CA2/s1[14] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_06_  (.A(\hash/p2_cap[8] ),
    .B(\hash/p2_cap[21] ),
    .C(\hash/p2_cap[26] ),
    .X(\hash/CA2/s1[15] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_07_  (.A(\hash/p2_cap[9] ),
    .B(\hash/p2_cap[22] ),
    .C(\hash/p2_cap[27] ),
    .X(\hash/CA2/s1[16] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_08_  (.A(\hash/p2_cap[10] ),
    .B(\hash/p2_cap[23] ),
    .C(\hash/p2_cap[28] ),
    .X(\hash/CA2/s1[17] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_09_  (.A(\hash/p2_cap[11] ),
    .B(\hash/p2_cap[24] ),
    .C(\hash/p2_cap[29] ),
    .X(\hash/CA2/s1[18] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_10_  (.A(\hash/p2_cap[12] ),
    .B(\hash/p2_cap[25] ),
    .C(\hash/p2_cap[30] ),
    .X(\hash/CA2/s1[19] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_11_  (.A(\hash/p2_cap[12] ),
    .B(\hash/p2_cap[7] ),
    .C(\hash/p2_cap[26] ),
    .X(\hash/CA2/s1[1] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_12_  (.A(\hash/p2_cap[13] ),
    .B(\hash/p2_cap[26] ),
    .C(\hash/p2_cap[31] ),
    .X(\hash/CA2/s1[20] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_13_  (.A(\hash/p2_cap[14] ),
    .B(\hash/p2_cap[27] ),
    .C(\hash/p2_cap[0] ),
    .X(\hash/CA2/s1[21] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_14_  (.A(\hash/p2_cap[15] ),
    .B(\hash/p2_cap[28] ),
    .C(\hash/p2_cap[1] ),
    .X(\hash/CA2/s1[22] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_15_  (.A(\hash/p2_cap[16] ),
    .B(\hash/p2_cap[29] ),
    .C(\hash/p2_cap[2] ),
    .X(\hash/CA2/s1[23] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_16_  (.A(\hash/p2_cap[17] ),
    .B(\hash/p2_cap[30] ),
    .C(\hash/p2_cap[3] ),
    .X(\hash/CA2/s1[24] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_17_  (.A(\hash/p2_cap[18] ),
    .B(\hash/p2_cap[31] ),
    .C(\hash/p2_cap[4] ),
    .X(\hash/CA2/s1[25] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_18_  (.A(\hash/p2_cap[19] ),
    .B(\hash/p2_cap[0] ),
    .C(\hash/p2_cap[5] ),
    .X(\hash/CA2/s1[26] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_19_  (.A(\hash/p2_cap[6] ),
    .B(\hash/p2_cap[20] ),
    .C(\hash/p2_cap[1] ),
    .X(\hash/CA2/s1[27] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_20_  (.A(\hash/p2_cap[7] ),
    .B(\hash/p2_cap[21] ),
    .C(\hash/p2_cap[2] ),
    .X(\hash/CA2/s1[28] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_21_  (.A(\hash/p2_cap[8] ),
    .B(\hash/p2_cap[22] ),
    .C(\hash/p2_cap[3] ),
    .X(\hash/CA2/s1[29] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_22_  (.A(\hash/p2_cap[13] ),
    .B(\hash/p2_cap[8] ),
    .C(\hash/p2_cap[27] ),
    .X(\hash/CA2/s1[2] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_23_  (.A(\hash/p2_cap[9] ),
    .B(\hash/p2_cap[23] ),
    .C(\hash/p2_cap[4] ),
    .X(\hash/CA2/s1[30] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_24_  (.A(\hash/p2_cap[10] ),
    .B(\hash/p2_cap[24] ),
    .C(\hash/p2_cap[5] ),
    .X(\hash/CA2/s1[31] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_25_  (.A(\hash/p2_cap[14] ),
    .B(\hash/p2_cap[9] ),
    .C(\hash/p2_cap[28] ),
    .X(\hash/CA2/s1[3] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_26_  (.A(\hash/p2_cap[15] ),
    .B(\hash/p2_cap[10] ),
    .C(\hash/p2_cap[29] ),
    .X(\hash/CA2/s1[4] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_27_  (.A(\hash/p2_cap[11] ),
    .B(\hash/p2_cap[16] ),
    .C(\hash/p2_cap[30] ),
    .X(\hash/CA2/s1[5] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_28_  (.A(\hash/p2_cap[12] ),
    .B(\hash/p2_cap[17] ),
    .C(\hash/p2_cap[31] ),
    .X(\hash/CA2/s1[6] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_29_  (.A(\hash/p2_cap[13] ),
    .B(\hash/p2_cap[18] ),
    .C(\hash/p2_cap[0] ),
    .X(\hash/CA2/s1[7] ));
 sky130_fd_sc_hd__xor3_4 \hash/CA2/S1/_30_  (.A(\hash/p2_cap[14] ),
    .B(\hash/p2_cap[19] ),
    .C(\hash/p2_cap[1] ),
    .X(\hash/CA2/s1[8] ));
 sky130_fd_sc_hd__xor3_1 \hash/CA2/S1/_31_  (.A(\hash/p2_cap[15] ),
    .B(\hash/p2_cap[20] ),
    .C(\hash/p2_cap[2] ),
    .X(\hash/CA2/s1[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1214_  (.A0(\hash/f_cap[0] ),
    .A1(\hash/e_cap[0] ),
    .S(\hash/p2_cap[0] ),
    .X(\hash/CA2/_0932_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1215_  (.A0(\hash/f_cap[1] ),
    .A1(\hash/e_cap[1] ),
    .S(\hash/p2_cap[1] ),
    .X(\hash/CA2/_0616_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1216_  (.A0(\hash/f_cap[2] ),
    .A1(\hash/e_cap[2] ),
    .S(\hash/p2_cap[2] ),
    .X(\hash/CA2/_0938_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1217_  (.A(\hash/CA2/_0940_ ),
    .B(\hash/CA2/_0617_ ),
    .X(\hash/CA2/_0640_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1218_  (.A(\hash/CA2/_0640_ ),
    .Y(\hash/CA2/_0637_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1219_  (.A0(\hash/f_cap[3] ),
    .A1(\hash/e_cap[3] ),
    .S(\hash/p2_cap[3] ),
    .X(\hash/CA2/_0943_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1220_  (.A1(\hash/CA2/_0615_ ),
    .A2(\hash/CA2/_0935_ ),
    .B1(\hash/CA2/_0934_ ),
    .X(\hash/CA2/_0523_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1221_  (.A1(\hash/CA2/_0940_ ),
    .A2(\hash/CA2/_0523_ ),
    .B1(\hash/CA2/_0939_ ),
    .Y(\hash/CA2/_0524_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1222_  (.A(\hash/CA2/_0945_ ),
    .B(\hash/CA2/_0524_ ),
    .Y(\hash/CA2/_0649_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1223_  (.A(\hash/CA2/_0649_ ),
    .Y(\hash/CA2/_0646_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1224_  (.A0(\hash/f_cap[4] ),
    .A1(\hash/e_cap[4] ),
    .S(\hash/p2_cap[4] ),
    .X(\hash/CA2/_0948_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1225_  (.A1(\hash/CA2/_0940_ ),
    .A2(\hash/CA2/_0617_ ),
    .B1(\hash/CA2/_0939_ ),
    .X(\hash/CA2/_0525_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1226_  (.A1(\hash/CA2/_0945_ ),
    .A2(\hash/CA2/_0525_ ),
    .B1(\hash/CA2/_0944_ ),
    .Y(\hash/CA2/_0526_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1227_  (.A(\hash/CA2/_0950_ ),
    .B(\hash/CA2/_0526_ ),
    .Y(\hash/CA2/_0658_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1228_  (.A(\hash/CA2/_0658_ ),
    .Y(\hash/CA2/_0655_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1229_  (.A0(\hash/f_cap[5] ),
    .A1(\hash/e_cap[5] ),
    .S(\hash/p2_cap[5] ),
    .X(\hash/CA2/_0953_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1230_  (.A0(\hash/f_cap[6] ),
    .A1(\hash/e_cap[6] ),
    .S(\hash/p2_cap[6] ),
    .X(\hash/CA2/_0958_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1231_  (.A0(\hash/f_cap[7] ),
    .A1(\hash/e_cap[7] ),
    .S(\hash/p2_cap[7] ),
    .X(\hash/CA2/_0963_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1232_  (.A0(\hash/f_cap[8] ),
    .A1(\hash/e_cap[8] ),
    .S(\hash/p2_cap[8] ),
    .X(\hash/CA2/_0968_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1233_  (.A(\hash/CA2/_0950_ ),
    .Y(\hash/CA2/_0527_ ));
 sky130_fd_sc_hd__nor4_1 \hash/CA2/_1234_  (.A(\hash/CA2/_0949_ ),
    .B(\hash/CA2/_0954_ ),
    .C(\hash/CA2/_0959_ ),
    .D(\hash/CA2/_0964_ ),
    .Y(\hash/CA2/_0528_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1235_  (.A1(\hash/CA2/_0527_ ),
    .A2(\hash/CA2/_0526_ ),
    .B1(\hash/CA2/_0528_ ),
    .Y(\hash/CA2/_0529_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1236_  (.A1(\hash/CA2/_0955_ ),
    .A2(\hash/CA2/_0954_ ),
    .B1(\hash/CA2/_0960_ ),
    .Y(\hash/CA2/_0530_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1237_  (.A(\hash/CA2/_0959_ ),
    .B(\hash/CA2/_0964_ ),
    .Y(\hash/CA2/_0531_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1238_  (.A(\hash/CA2/_0965_ ),
    .B(\hash/CA2/_0964_ ),
    .Y(\hash/CA2/_0532_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1239_  (.A1(\hash/CA2/_0530_ ),
    .A2(\hash/CA2/_0531_ ),
    .B1(\hash/CA2/_0532_ ),
    .Y(\hash/CA2/_0533_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_1240_  (.A(\hash/CA2/_0529_ ),
    .B(\hash/CA2/_0533_ ),
    .X(\hash/CA2/_0534_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1241_  (.A(\hash/CA2/_0970_ ),
    .B(\hash/CA2/_0534_ ),
    .X(\hash/CA2/_0687_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1242_  (.A(\hash/CA2/_0687_ ),
    .Y(\hash/CA2/_0684_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1243_  (.A0(\hash/f_cap[9] ),
    .A1(\hash/e_cap[9] ),
    .S(\hash/p2_cap[9] ),
    .X(\hash/CA2/_0973_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1244_  (.A(\hash/CA2/_0950_ ),
    .B(\hash/CA2/_0949_ ),
    .C(\hash/CA2/_0954_ ),
    .Y(\hash/CA2/_0535_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1245_  (.A(\hash/CA2/_0530_ ),
    .B(\hash/CA2/_0535_ ),
    .Y(\hash/CA2/_0536_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1246_  (.A1(\hash/CA2/_0615_ ),
    .A2(\hash/CA2/_0935_ ),
    .B1(\hash/CA2/_0934_ ),
    .C1(\hash/CA2/_0939_ ),
    .Y(\hash/CA2/_0537_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1247_  (.A1(\hash/CA2/_0940_ ),
    .A2(\hash/CA2/_0939_ ),
    .B1(\hash/CA2/_0945_ ),
    .Y(\hash/CA2/_0538_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1248_  (.A(\hash/CA2/_0944_ ),
    .B(\hash/CA2/_0949_ ),
    .C(\hash/CA2/_0954_ ),
    .Y(\hash/CA2/_0539_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA2/_1249_  (.A1(\hash/CA2/_0537_ ),
    .A2(\hash/CA2/_0538_ ),
    .B1(\hash/CA2/_0539_ ),
    .Y(\hash/CA2/_0540_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1250_  (.A1(\hash/CA2/_0536_ ),
    .A2(\hash/CA2/_0540_ ),
    .B1(\hash/CA2/_0959_ ),
    .Y(\hash/CA2/_0541_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1251_  (.A(\hash/CA2/_0541_ ),
    .B_N(\hash/CA2/_0965_ ),
    .Y(\hash/CA2/_0542_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1252_  (.A1(\hash/CA2/_0964_ ),
    .A2(\hash/CA2/_0542_ ),
    .B1(\hash/CA2/_0970_ ),
    .X(\hash/CA2/_0543_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1253_  (.A(\hash/CA2/_0969_ ),
    .B(\hash/CA2/_0543_ ),
    .Y(\hash/CA2/_0544_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1254_  (.A(\hash/CA2/_0975_ ),
    .B(\hash/CA2/_0544_ ),
    .Y(\hash/CA2/_0976_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1255_  (.A(\hash/CA2/_0976_ ),
    .Y(\hash/CA2/_0693_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1256_  (.A0(\hash/f_cap[10] ),
    .A1(\hash/e_cap[10] ),
    .S(\hash/p2_cap[10] ),
    .X(\hash/CA2/_0979_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1257_  (.A1(\hash/CA2/_0970_ ),
    .A2(\hash/CA2/_0534_ ),
    .B1(\hash/CA2/_0969_ ),
    .X(\hash/CA2/_0545_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1258_  (.A1(\hash/CA2/_0975_ ),
    .A2(\hash/CA2/_0545_ ),
    .B1(\hash/CA2/_0974_ ),
    .X(\hash/CA2/_0546_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1259_  (.A(\hash/CA2/_0981_ ),
    .B(\hash/CA2/_0546_ ),
    .X(\hash/CA2/_0982_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1260_  (.A(\hash/CA2/_0982_ ),
    .Y(\hash/CA2/_0701_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1261_  (.A0(\hash/f_cap[11] ),
    .A1(\hash/e_cap[11] ),
    .S(\hash/p2_cap[11] ),
    .X(\hash/CA2/_0985_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_1262_  (.A(\hash/CA2/_0970_ ),
    .B(\hash/CA2/_0975_ ),
    .C(\hash/CA2/_0981_ ),
    .X(\hash/CA2/_0547_ ));
 sky130_fd_sc_hd__and4_1 \hash/CA2/_1263_  (.A(\hash/CA2/_0965_ ),
    .B(\hash/CA2/_0536_ ),
    .C(\hash/CA2/_0540_ ),
    .D(\hash/CA2/_0547_ ),
    .X(\hash/CA2/_0548_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1264_  (.A1(\hash/CA2/_0975_ ),
    .A2(\hash/CA2/_0969_ ),
    .B1(\hash/CA2/_0974_ ),
    .X(\hash/CA2/_0549_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_1265_  (.A(\hash/CA2/_0970_ ),
    .B(\hash/CA2/_0975_ ),
    .C(\hash/CA2/_0964_ ),
    .X(\hash/CA2/_0550_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1266_  (.A1(\hash/CA2/_0549_ ),
    .A2(\hash/CA2/_0550_ ),
    .B1(\hash/CA2/_0981_ ),
    .Y(\hash/CA2/_0551_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA2/_1267_  (.A1(\hash/CA2/_0965_ ),
    .A2(\hash/CA2/_0959_ ),
    .A3(\hash/CA2/_0547_ ),
    .B1(\hash/CA2/_0980_ ),
    .Y(\hash/CA2/_0552_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1268_  (.A(\hash/CA2/_0551_ ),
    .B(\hash/CA2/_0552_ ),
    .Y(\hash/CA2/_0553_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA2/_1269_  (.A(\hash/CA2/_0548_ ),
    .B(\hash/CA2/_0553_ ),
    .X(\hash/CA2/_0554_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1270_  (.A(\hash/CA2/_0987_ ),
    .B(\hash/CA2/_0554_ ),
    .X(\hash/CA2/_0988_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1271_  (.A(\hash/CA2/_0988_ ),
    .Y(\hash/CA2/_0709_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1272_  (.A0(\hash/f_cap[12] ),
    .A1(\hash/e_cap[12] ),
    .S(\hash/p2_cap[12] ),
    .X(\hash/CA2/_0991_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1273_  (.A1(\hash/CA2/_0981_ ),
    .A2(\hash/CA2/_0549_ ),
    .B1(\hash/CA2/_0980_ ),
    .X(\hash/CA2/_0555_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1274_  (.A1(\hash/CA2/_0987_ ),
    .A2(\hash/CA2/_0555_ ),
    .B1(\hash/CA2/_0986_ ),
    .X(\hash/CA2/_0556_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA2/_1275_  (.A1(\hash/CA2/_0987_ ),
    .A2(\hash/CA2/_0534_ ),
    .A3(\hash/CA2/_0547_ ),
    .B1(\hash/CA2/_0556_ ),
    .Y(\hash/CA2/_0557_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1276_  (.A(\hash/CA2/_0993_ ),
    .B(\hash/CA2/_0557_ ),
    .Y(\hash/CA2/_0994_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1277_  (.A(\hash/CA2/_0994_ ),
    .Y(\hash/CA2/_0717_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1278_  (.A0(\hash/f_cap[13] ),
    .A1(\hash/e_cap[13] ),
    .S(\hash/p2_cap[13] ),
    .X(\hash/CA2/_0997_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1279_  (.A(\hash/CA2/_0993_ ),
    .Y(\hash/CA2/_0558_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1280_  (.A1(\hash/CA2/_0987_ ),
    .A2(\hash/CA2/_0554_ ),
    .B1(\hash/CA2/_0986_ ),
    .Y(\hash/CA2/_0559_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1281_  (.A1(\hash/CA2/_0558_ ),
    .A2(\hash/CA2/_0559_ ),
    .B1_N(\hash/CA2/_0992_ ),
    .Y(\hash/CA2/_0560_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1282_  (.A(\hash/CA2/_0999_ ),
    .B(\hash/CA2/_0560_ ),
    .X(\hash/CA2/_1000_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1283_  (.A(\hash/CA2/_1000_ ),
    .Y(\hash/CA2/_0725_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1284_  (.A0(\hash/f_cap[14] ),
    .A1(\hash/e_cap[14] ),
    .S(\hash/p2_cap[14] ),
    .X(\hash/CA2/_1003_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1285_  (.A1(\hash/CA2/_0558_ ),
    .A2(\hash/CA2/_0557_ ),
    .B1_N(\hash/CA2/_0992_ ),
    .Y(\hash/CA2/_0561_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1286_  (.A1(\hash/CA2/_0999_ ),
    .A2(\hash/CA2/_0561_ ),
    .B1(\hash/CA2/_0998_ ),
    .Y(\hash/CA2/_0562_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1287_  (.A(\hash/CA2/_1005_ ),
    .B(\hash/CA2/_0562_ ),
    .Y(\hash/CA2/_1006_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1288_  (.A(\hash/CA2/_1006_ ),
    .Y(\hash/CA2/_0733_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1289_  (.A0(\hash/f_cap[15] ),
    .A1(\hash/e_cap[15] ),
    .S(\hash/p2_cap[15] ),
    .X(\hash/CA2/_1009_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1290_  (.A(\hash/CA2/_0999_ ),
    .B(\hash/CA2/_1005_ ),
    .Y(\hash/CA2/_0563_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1291_  (.A(\hash/CA2/_0558_ ),
    .B(\hash/CA2/_0563_ ),
    .Y(\hash/CA2/_0564_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_1292_  (.A(\hash/CA2/_0987_ ),
    .B(\hash/CA2/_0564_ ),
    .X(\hash/CA2/_0565_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1293_  (.A1(\hash/CA2/_0993_ ),
    .A2(\hash/CA2/_0986_ ),
    .B1(\hash/CA2/_0992_ ),
    .Y(\hash/CA2/_0566_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1294_  (.A1(\hash/CA2/_1005_ ),
    .A2(\hash/CA2/_0998_ ),
    .B1(\hash/CA2/_1004_ ),
    .Y(\hash/CA2/_0567_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1295_  (.A1(\hash/CA2/_0563_ ),
    .A2(\hash/CA2/_0566_ ),
    .B1(\hash/CA2/_0567_ ),
    .Y(\hash/CA2/_0568_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1296_  (.A1(\hash/CA2/_0554_ ),
    .A2(\hash/CA2/_0565_ ),
    .B1(\hash/CA2/_0568_ ),
    .Y(\hash/CA2/_0569_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1297_  (.A(\hash/CA2/_1011_ ),
    .B(\hash/CA2/_0569_ ),
    .Y(\hash/CA2/_1012_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1298_  (.A(\hash/CA2/_1012_ ),
    .Y(\hash/CA2/_0741_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1299_  (.A0(\hash/f_cap[16] ),
    .A1(\hash/e_cap[16] ),
    .S(\hash/p2_cap[16] ),
    .X(\hash/CA2/_1015_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1300_  (.A1(\hash/CA2/_0999_ ),
    .A2(\hash/CA2/_0992_ ),
    .B1(\hash/CA2/_0998_ ),
    .X(\hash/CA2/_0570_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA2/_1301_  (.A1(\hash/CA2/_0556_ ),
    .A2(\hash/CA2/_0564_ ),
    .B1(\hash/CA2/_0570_ ),
    .B2(\hash/CA2/_1005_ ),
    .C1(\hash/CA2/_1004_ ),
    .Y(\hash/CA2/_0571_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA2/_1302_  (.A(\hash/CA2/_0529_ ),
    .B(\hash/CA2/_0533_ ),
    .C(\hash/CA2/_0547_ ),
    .D(\hash/CA2/_0565_ ),
    .Y(\hash/CA2/_0572_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1303_  (.A(\hash/CA2/_1011_ ),
    .Y(\hash/CA2/_0573_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1304_  (.A1(\hash/CA2/_0571_ ),
    .A2(\hash/CA2/_0572_ ),
    .B1(\hash/CA2/_0573_ ),
    .Y(\hash/CA2/_0574_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1305_  (.A(\hash/CA2/_1010_ ),
    .B(\hash/CA2/_0574_ ),
    .Y(\hash/CA2/_0575_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1306_  (.A(\hash/CA2/_1017_ ),
    .B(\hash/CA2/_0575_ ),
    .Y(\hash/CA2/_0752_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1307_  (.A(\hash/CA2/_0752_ ),
    .Y(\hash/CA2/_0749_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1308_  (.A0(\hash/f_cap[17] ),
    .A1(\hash/e_cap[17] ),
    .S(\hash/p2_cap[17] ),
    .X(\hash/CA2/_1020_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1309_  (.A(\hash/CA2/_1016_ ),
    .Y(\hash/CA2/_0576_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA2/_1310_  (.A1(\hash/CA2/_0548_ ),
    .A2(\hash/CA2/_0553_ ),
    .B1(\hash/CA2/_0565_ ),
    .Y(\hash/CA2/_0577_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1311_  (.A(\hash/CA2/_0568_ ),
    .Y(\hash/CA2/_0578_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1312_  (.A1(\hash/CA2/_0577_ ),
    .A2(\hash/CA2/_0578_ ),
    .B1(\hash/CA2/_0573_ ),
    .Y(\hash/CA2/_0579_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1313_  (.A1(\hash/CA2/_1010_ ),
    .A2(\hash/CA2/_0579_ ),
    .B1(\hash/CA2/_1017_ ),
    .Y(\hash/CA2/_0580_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1314_  (.A(\hash/CA2/_0576_ ),
    .B(\hash/CA2/_0580_ ),
    .Y(\hash/CA2/_0581_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1315_  (.A(\hash/CA2/_1022_ ),
    .B(\hash/CA2/_0581_ ),
    .X(\hash/CA2/_1023_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1316_  (.A(\hash/CA2/_1023_ ),
    .Y(\hash/CA2/_0758_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1317_  (.A0(\hash/f_cap[18] ),
    .A1(\hash/e_cap[18] ),
    .S(\hash/p2_cap[18] ),
    .X(\hash/CA2/_1026_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1318_  (.A(\hash/CA2/_1017_ ),
    .Y(\hash/CA2/_0582_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1319_  (.A1(\hash/CA2/_0582_ ),
    .A2(\hash/CA2/_0575_ ),
    .B1(\hash/CA2/_0576_ ),
    .Y(\hash/CA2/_0583_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1320_  (.A1(\hash/CA2/_1022_ ),
    .A2(\hash/CA2/_0583_ ),
    .B1(\hash/CA2/_1021_ ),
    .Y(\hash/CA2/_0584_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1321_  (.A(\hash/CA2/_1028_ ),
    .B(\hash/CA2/_0584_ ),
    .Y(\hash/CA2/_1029_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1322_  (.A(\hash/CA2/_1029_ ),
    .Y(\hash/CA2/_0766_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1323_  (.A0(\hash/f_cap[19] ),
    .A1(\hash/e_cap[19] ),
    .S(\hash/p2_cap[19] ),
    .X(\hash/CA2/_1032_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1324_  (.A(\hash/CA2/_1022_ ),
    .B(\hash/CA2/_1028_ ),
    .Y(\hash/CA2/_0585_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1325_  (.A1(\hash/CA2/_0576_ ),
    .A2(\hash/CA2/_0580_ ),
    .B1(\hash/CA2/_0585_ ),
    .Y(\hash/CA2/_0586_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_1326_  (.A(\hash/CA2/_1028_ ),
    .B(\hash/CA2/_1021_ ),
    .X(\hash/CA2/_0587_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1327_  (.A(\hash/CA2/_1027_ ),
    .B(\hash/CA2/_0586_ ),
    .C(\hash/CA2/_0587_ ),
    .Y(\hash/CA2/_0588_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1328_  (.A(\hash/CA2/_1034_ ),
    .B(\hash/CA2/_0588_ ),
    .Y(\hash/CA2/_1035_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1329_  (.A(\hash/CA2/_1035_ ),
    .Y(\hash/CA2/_0774_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1330_  (.A0(\hash/f_cap[20] ),
    .A1(\hash/e_cap[20] ),
    .S(\hash/p2_cap[20] ),
    .X(\hash/CA2/_1038_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1331_  (.A1(\hash/CA2/_1022_ ),
    .A2(\hash/CA2/_1016_ ),
    .B1(\hash/CA2/_1021_ ),
    .Y(\hash/CA2/_0589_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1332_  (.A(\hash/CA2/_1028_ ),
    .B(\hash/CA2/_1034_ ),
    .Y(\hash/CA2/_0590_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1333_  (.A1(\hash/CA2/_1034_ ),
    .A2(\hash/CA2/_1027_ ),
    .B1(\hash/CA2/_1033_ ),
    .Y(\hash/CA2/_0591_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1334_  (.A1(\hash/CA2/_0589_ ),
    .A2(\hash/CA2/_0590_ ),
    .B1(\hash/CA2/_0591_ ),
    .X(\hash/CA2/_0592_ ));
 sky130_fd_sc_hd__and4_4 \hash/CA2/_1335_  (.A(\hash/CA2/_1017_ ),
    .B(\hash/CA2/_1022_ ),
    .C(\hash/CA2/_1028_ ),
    .D(\hash/CA2/_1034_ ),
    .X(\hash/CA2/_0593_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1336_  (.A1(\hash/CA2/_1010_ ),
    .A2(\hash/CA2/_0574_ ),
    .B1(\hash/CA2/_0593_ ),
    .Y(\hash/CA2/_0594_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1337_  (.A(\hash/CA2/_0592_ ),
    .B(\hash/CA2/_0594_ ),
    .Y(\hash/CA2/_0595_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1338_  (.A(\hash/CA2/_1040_ ),
    .B(\hash/CA2/_0595_ ),
    .X(\hash/CA2/_1041_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1339_  (.A(\hash/CA2/_1041_ ),
    .Y(\hash/CA2/_0782_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1340_  (.A0(\hash/f_cap[21] ),
    .A1(\hash/e_cap[21] ),
    .S(\hash/p2_cap[21] ),
    .X(\hash/CA2/_1044_ ));
 sky130_fd_sc_hd__or3_1 \hash/CA2/_1341_  (.A(\hash/CA2/_1027_ ),
    .B(\hash/CA2/_1033_ ),
    .C(\hash/CA2/_1039_ ),
    .X(\hash/CA2/_0596_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1342_  (.A(\hash/CA2/_1034_ ),
    .B(\hash/CA2/_1033_ ),
    .C(\hash/CA2/_1039_ ),
    .Y(\hash/CA2/_0597_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1343_  (.A(\hash/CA2/_1040_ ),
    .B(\hash/CA2/_1039_ ),
    .Y(\hash/CA2/_0598_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1344_  (.A(\hash/CA2/_0597_ ),
    .B(\hash/CA2/_0598_ ),
    .Y(\hash/CA2/_0599_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_1345_  (.A1(\hash/CA2/_0586_ ),
    .A2(\hash/CA2/_0587_ ),
    .A3(\hash/CA2/_0596_ ),
    .B1(\hash/CA2/_0599_ ),
    .Y(\hash/CA2/_0600_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1346_  (.A(\hash/CA2/_1046_ ),
    .B(\hash/CA2/_0600_ ),
    .Y(\hash/CA2/_1047_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1347_  (.A(\hash/CA2/_1047_ ),
    .Y(\hash/CA2/_0790_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1348_  (.A0(\hash/f_cap[22] ),
    .A1(\hash/e_cap[22] ),
    .S(\hash/p2_cap[22] ),
    .X(\hash/CA2/_1050_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1349_  (.A(\hash/CA2/_1011_ ),
    .B(\hash/CA2/_1040_ ),
    .C(\hash/CA2/_0593_ ),
    .Y(\hash/CA2/_0601_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1350_  (.A1(\hash/CA2/_0571_ ),
    .A2(\hash/CA2/_0572_ ),
    .B1(\hash/CA2/_0601_ ),
    .Y(\hash/CA2/_0602_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1351_  (.A(\hash/CA2/_1010_ ),
    .B(\hash/CA2/_0593_ ),
    .Y(\hash/CA2/_0603_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1352_  (.A(\hash/CA2/_0592_ ),
    .B(\hash/CA2/_0603_ ),
    .Y(\hash/CA2/_0604_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1353_  (.A1(\hash/CA2/_1040_ ),
    .A2(\hash/CA2/_0604_ ),
    .B1(\hash/CA2/_1039_ ),
    .X(\hash/CA2/_0605_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1354_  (.A1(\hash/CA2/_0602_ ),
    .A2(\hash/CA2/_0605_ ),
    .B1(\hash/CA2/_1046_ ),
    .X(\hash/CA2/_0606_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1355_  (.A(\hash/CA2/_1045_ ),
    .B(\hash/CA2/_0606_ ),
    .Y(\hash/CA2/_0607_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1356_  (.A(\hash/CA2/_1052_ ),
    .B(\hash/CA2/_0607_ ),
    .Y(\hash/CA2/_1053_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1357_  (.A(\hash/CA2/_1053_ ),
    .Y(\hash/CA2/_0798_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1358_  (.A0(\hash/f_cap[23] ),
    .A1(\hash/e_cap[23] ),
    .S(\hash/p2_cap[23] ),
    .X(\hash/CA2/_1056_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1359_  (.A(\hash/CA2/_1039_ ),
    .B(\hash/CA2/_1045_ ),
    .Y(\hash/CA2/_0608_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1360_  (.A(\hash/CA2/_1040_ ),
    .B(\hash/CA2/_1039_ ),
    .C(\hash/CA2/_1045_ ),
    .Y(\hash/CA2/_0609_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1361_  (.A(\hash/CA2/_1046_ ),
    .B(\hash/CA2/_1045_ ),
    .Y(\hash/CA2/_0000_ ));
 sky130_fd_sc_hd__a311oi_2 \hash/CA2/_1362_  (.A1(\hash/CA2/_0592_ ),
    .A2(\hash/CA2/_0603_ ),
    .A3(\hash/CA2/_0608_ ),
    .B1(\hash/CA2/_0609_ ),
    .C1(\hash/CA2/_0000_ ),
    .Y(\hash/CA2/_0001_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1363_  (.A(\hash/CA2/_1051_ ),
    .B(\hash/CA2/_0568_ ),
    .C(\hash/CA2/_0001_ ),
    .Y(\hash/CA2/_0002_ ));
 sky130_fd_sc_hd__a41o_1 \hash/CA2/_1364_  (.A1(\hash/CA2/_1011_ ),
    .A2(\hash/CA2/_1040_ ),
    .A3(\hash/CA2/_1046_ ),
    .A4(\hash/CA2/_0593_ ),
    .B1(\hash/CA2/_1051_ ),
    .X(\hash/CA2/_0003_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA2/_1365_  (.A1(\hash/CA2/_1052_ ),
    .A2(\hash/CA2/_1051_ ),
    .B1(\hash/CA2/_0001_ ),
    .B2(\hash/CA2/_0003_ ),
    .Y(\hash/CA2/_0004_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1366_  (.A1(\hash/CA2/_0577_ ),
    .A2(\hash/CA2/_0002_ ),
    .B1(\hash/CA2/_0004_ ),
    .X(\hash/CA2/_0005_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1367_  (.A(\hash/CA2/_1058_ ),
    .B(\hash/CA2/_0005_ ),
    .Y(\hash/CA2/_1059_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1368_  (.A(\hash/CA2/_1059_ ),
    .Y(\hash/CA2/_0806_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1369_  (.A0(\hash/f_cap[24] ),
    .A1(\hash/e_cap[24] ),
    .S(\hash/p2_cap[24] ),
    .X(\hash/CA2/_1062_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1370_  (.A(\hash/CA2/_0000_ ),
    .B_N(\hash/CA2/_1052_ ),
    .Y(\hash/CA2/_0006_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_1371_  (.A1(\hash/CA2/_1045_ ),
    .A2(\hash/CA2/_0602_ ),
    .A3(\hash/CA2/_0605_ ),
    .B1(\hash/CA2/_0006_ ),
    .Y(\hash/CA2/_0007_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1372_  (.A_N(\hash/CA2/_1051_ ),
    .B(\hash/CA2/_0007_ ),
    .Y(\hash/CA2/_0008_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1373_  (.A1(\hash/CA2/_1058_ ),
    .A2(\hash/CA2/_0008_ ),
    .B1(\hash/CA2/_1057_ ),
    .X(\hash/CA2/_0009_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1374_  (.A(\hash/CA2/_1064_ ),
    .B(\hash/CA2/_0009_ ),
    .X(\hash/CA2/_1065_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1375_  (.A(\hash/CA2/_1065_ ),
    .Y(\hash/CA2/_0814_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1376_  (.A0(\hash/f_cap[25] ),
    .A1(\hash/e_cap[25] ),
    .S(\hash/p2_cap[25] ),
    .X(\hash/CA2/_1068_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1377_  (.A1(\hash/CA2/_1051_ ),
    .A2(\hash/CA2/_0006_ ),
    .B1(\hash/CA2/_1058_ ),
    .X(\hash/CA2/_0010_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1378_  (.A1(\hash/CA2/_1057_ ),
    .A2(\hash/CA2/_0010_ ),
    .B1(\hash/CA2/_1064_ ),
    .Y(\hash/CA2/_0011_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1379_  (.A(\hash/CA2/_1070_ ),
    .B(\hash/CA2/_0011_ ),
    .Y(\hash/CA2/_0012_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1380_  (.A(\hash/CA2/_1070_ ),
    .Y(\hash/CA2/_0013_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1381_  (.A1(\hash/CA2/_1052_ ),
    .A2(\hash/CA2/_1045_ ),
    .B1(\hash/CA2/_1051_ ),
    .X(\hash/CA2/_0014_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1382_  (.A1(\hash/CA2/_1058_ ),
    .A2(\hash/CA2/_0014_ ),
    .B1(\hash/CA2/_1057_ ),
    .Y(\hash/CA2/_0015_ ));
 sky130_fd_sc_hd__nor3b_1 \hash/CA2/_1383_  (.A(\hash/CA2/_0013_ ),
    .B(\hash/CA2/_1063_ ),
    .C_N(\hash/CA2/_0015_ ),
    .Y(\hash/CA2/_0016_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1384_  (.A0(\hash/CA2/_0012_ ),
    .A1(\hash/CA2/_0016_ ),
    .S(\hash/CA2/_0600_ ),
    .X(\hash/CA2/_0017_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA2/_1385_  (.A_N(\hash/CA2/_1063_ ),
    .B(\hash/CA2/_0011_ ),
    .C(\hash/CA2/_1070_ ),
    .Y(\hash/CA2/_0018_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1386_  (.A(\hash/CA2/_0013_ ),
    .B(\hash/CA2/_1063_ ),
    .Y(\hash/CA2/_0019_ ));
 sky130_fd_sc_hd__o311ai_0 \hash/CA2/_1387_  (.A1(\hash/CA2/_1070_ ),
    .A2(\hash/CA2/_0011_ ),
    .A3(\hash/CA2/_0015_ ),
    .B1(\hash/CA2/_0018_ ),
    .C1(\hash/CA2/_0019_ ),
    .Y(\hash/CA2/_0020_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1388_  (.A(\hash/CA2/_0017_ ),
    .B(\hash/CA2/_0020_ ),
    .Y(\hash/CA2/_0822_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1389_  (.A0(\hash/f_cap[26] ),
    .A1(\hash/e_cap[26] ),
    .S(\hash/p2_cap[26] ),
    .X(\hash/CA2/_1074_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1390_  (.A(\hash/CA2/_1051_ ),
    .B(\hash/CA2/_1057_ ),
    .C(\hash/CA2/_1063_ ),
    .Y(\hash/CA2/_0021_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA2/_1391_  (.A(\hash/CA2/_1058_ ),
    .B(\hash/CA2/_1057_ ),
    .X(\hash/CA2/_0022_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1392_  (.A1(\hash/CA2/_1064_ ),
    .A2(\hash/CA2/_0022_ ),
    .B1(\hash/CA2/_1063_ ),
    .Y(\hash/CA2/_0023_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1393_  (.A1(\hash/CA2/_0007_ ),
    .A2(\hash/CA2/_0021_ ),
    .B1(\hash/CA2/_0023_ ),
    .Y(\hash/CA2/_0024_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1394_  (.A1(\hash/CA2/_1070_ ),
    .A2(\hash/CA2/_0024_ ),
    .B1(\hash/CA2/_1069_ ),
    .Y(\hash/CA2/_0025_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1395_  (.A(\hash/CA2/_1076_ ),
    .B(\hash/CA2/_0025_ ),
    .Y(\hash/CA2/_1077_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1396_  (.A(\hash/CA2/_1077_ ),
    .Y(\hash/CA2/_0830_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1397_  (.A0(\hash/f_cap[27] ),
    .A1(\hash/e_cap[27] ),
    .S(\hash/p2_cap[27] ),
    .X(\hash/CA2/_1080_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1398_  (.A(\hash/CA2/_1058_ ),
    .B(\hash/CA2/_1064_ ),
    .C(\hash/CA2/_1070_ ),
    .Y(\hash/CA2/_0026_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1399_  (.A1(\hash/CA2/_1064_ ),
    .A2(\hash/CA2/_1057_ ),
    .B1(\hash/CA2/_1063_ ),
    .Y(\hash/CA2/_0027_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1400_  (.A(\hash/CA2/_0013_ ),
    .B(\hash/CA2/_0027_ ),
    .Y(\hash/CA2/_0028_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1401_  (.A(\hash/CA2/_1069_ ),
    .B(\hash/CA2/_0028_ ),
    .Y(\hash/CA2/_0029_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1402_  (.A1(\hash/CA2/_0005_ ),
    .A2(\hash/CA2/_0026_ ),
    .B1(\hash/CA2/_0029_ ),
    .Y(\hash/CA2/_0030_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1403_  (.A1(\hash/CA2/_1076_ ),
    .A2(\hash/CA2/_0030_ ),
    .B1(\hash/CA2/_1075_ ),
    .Y(\hash/CA2/_0031_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1404_  (.A(\hash/CA2/_1082_ ),
    .B(\hash/CA2/_0031_ ),
    .Y(\hash/CA2/_1083_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1405_  (.A(\hash/CA2/_1083_ ),
    .Y(\hash/CA2/_0838_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1406_  (.A0(\hash/f_cap[28] ),
    .A1(\hash/e_cap[28] ),
    .S(\hash/p2_cap[28] ),
    .X(\hash/CA2/_1086_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1407_  (.A(\hash/CA2/_1076_ ),
    .B(\hash/CA2/_1082_ ),
    .Y(\hash/CA2/_0032_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1408_  (.A1(\hash/CA2/_1082_ ),
    .A2(\hash/CA2/_1075_ ),
    .B1(\hash/CA2/_1081_ ),
    .Y(\hash/CA2/_0033_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1409_  (.A1(\hash/CA2/_0025_ ),
    .A2(\hash/CA2/_0032_ ),
    .B1(\hash/CA2/_0033_ ),
    .Y(\hash/CA2/_0034_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1410_  (.A(\hash/CA2/_1088_ ),
    .B(\hash/CA2/_0034_ ),
    .Y(\hash/CA2/_0846_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1411_  (.A0(\hash/f_cap[29] ),
    .A1(\hash/e_cap[29] ),
    .S(\hash/p2_cap[29] ),
    .X(\hash/CA2/_1091_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1412_  (.A1(\hash/CA2/_1088_ ),
    .A2(\hash/CA2/_1081_ ),
    .B1(\hash/CA2/_1087_ ),
    .Y(\hash/CA2/_0035_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1413_  (.A1(\hash/CA2/_0577_ ),
    .A2(\hash/CA2/_0002_ ),
    .B1(\hash/CA2/_0004_ ),
    .Y(\hash/CA2/_0036_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1414_  (.A(\hash/CA2/_1076_ ),
    .B(\hash/CA2/_1082_ ),
    .C(\hash/CA2/_1088_ ),
    .Y(\hash/CA2/_0037_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1415_  (.A(\hash/CA2/_0026_ ),
    .B(\hash/CA2/_0037_ ),
    .Y(\hash/CA2/_0038_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1416_  (.A(\hash/CA2/_1082_ ),
    .B(\hash/CA2/_1088_ ),
    .C(\hash/CA2/_1075_ ),
    .Y(\hash/CA2/_0039_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1417_  (.A1(\hash/CA2/_0029_ ),
    .A2(\hash/CA2/_0037_ ),
    .B1(\hash/CA2/_0039_ ),
    .Y(\hash/CA2/_0040_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1418_  (.A1(\hash/CA2/_0036_ ),
    .A2(\hash/CA2/_0038_ ),
    .B1(\hash/CA2/_0040_ ),
    .Y(\hash/CA2/_0041_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_1419_  (.A(\hash/CA2/_0035_ ),
    .B(\hash/CA2/_0041_ ),
    .X(\hash/CA2/_0042_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1420_  (.A(\hash/CA2/_1093_ ),
    .B(\hash/CA2/_0042_ ),
    .Y(\hash/CA2/_0858_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1421_  (.A(\hash/CA2/_0858_ ),
    .Y(\hash/CA2/_0855_ ));
 sky130_fd_sc_hd__mux2_2 \hash/CA2/_1422_  (.A0(\hash/f_cap[30] ),
    .A1(\hash/e_cap[30] ),
    .S(\hash/p2_cap[30] ),
    .X(\hash/CA2/_1096_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1423_  (.A1(\hash/a_cap[0] ),
    .A2(\hash/b_new[0] ),
    .B1(\hash/b_cap[0] ),
    .X(\hash/CA2/_0043_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1424_  (.A1(\hash/a_cap[0] ),
    .A2(\hash/b_new[0] ),
    .B1(\hash/CA2/_0043_ ),
    .Y(\hash/CA2/_0621_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1425_  (.A(\hash/CA2/_0614_ ),
    .Y(\hash/b_new[1] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1426_  (.A1(\hash/a_cap[1] ),
    .A2(\hash/b_new[1] ),
    .B1(\hash/b_cap[1] ),
    .X(\hash/CA2/_0044_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1427_  (.A1(\hash/a_cap[1] ),
    .A2(\hash/b_new[1] ),
    .B1(\hash/CA2/_0044_ ),
    .Y(\hash/CA2/_0626_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1428_  (.A(\hash/CA2/_0613_ ),
    .B(\hash/CA2/_0875_ ),
    .Y(\hash/b_new[2] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1429_  (.A(\hash/b_cap[2] ),
    .B(\hash/a_cap[2] ),
    .C(\hash/b_new[2] ),
    .X(\hash/CA2/_0045_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1430_  (.A(\hash/CA2/_0045_ ),
    .Y(\hash/CA2/_0634_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1431_  (.A1(\hash/CA2/_0871_ ),
    .A2(\hash/CA2/_0873_ ),
    .B1(\hash/CA2/_0872_ ),
    .C1(\hash/CA2/_0874_ ),
    .Y(\hash/CA2/_0046_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1432_  (.A1(\hash/CA2/_0875_ ),
    .A2(\hash/CA2/_0874_ ),
    .B1(\hash/CA2/_0877_ ),
    .Y(\hash/CA2/_0047_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1433_  (.A(\hash/CA2/_0046_ ),
    .B(\hash/CA2/_0047_ ),
    .Y(\hash/CA2/_0048_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1434_  (.A1(\hash/CA2/_0871_ ),
    .A2(\hash/CA2/_0873_ ),
    .B1(\hash/CA2/_0872_ ),
    .X(\hash/CA2/_0049_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1435_  (.A1(\hash/CA2/_0875_ ),
    .A2(\hash/CA2/_0049_ ),
    .B1(\hash/CA2/_0874_ ),
    .C1(\hash/CA2/_0877_ ),
    .Y(\hash/CA2/_0050_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1436_  (.A(\hash/CA2/_0048_ ),
    .B(\hash/CA2/_0050_ ),
    .Y(\hash/b_new[3] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1437_  (.A(\hash/b_cap[3] ),
    .B(\hash/a_cap[3] ),
    .C(\hash/b_new[3] ),
    .X(\hash/CA2/_0051_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1438_  (.A(\hash/CA2/_0051_ ),
    .Y(\hash/CA2/_0643_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1439_  (.A(\hash/CA2/_0613_ ),
    .B_N(\hash/CA2/_0875_ ),
    .Y(\hash/CA2/_0052_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1440_  (.A1(\hash/CA2/_0874_ ),
    .A2(\hash/CA2/_0052_ ),
    .B1(\hash/CA2/_0877_ ),
    .X(\hash/CA2/_0053_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1441_  (.A(\hash/CA2/_0876_ ),
    .B(\hash/CA2/_0053_ ),
    .Y(\hash/CA2/_0054_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1442_  (.A(\hash/CA2/_0879_ ),
    .B(\hash/CA2/_0054_ ),
    .Y(\hash/b_new[4] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1443_  (.A(\hash/b_cap[4] ),
    .B(\hash/a_cap[4] ),
    .C(\hash/b_new[4] ),
    .X(\hash/CA2/_0055_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1444_  (.A(\hash/CA2/_0055_ ),
    .Y(\hash/CA2/_0652_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1445_  (.A1(\hash/CA2/_0876_ ),
    .A2(\hash/CA2/_0053_ ),
    .B1(\hash/CA2/_0879_ ),
    .Y(\hash/CA2/_0056_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1446_  (.A(\hash/CA2/_0878_ ),
    .B(\hash/CA2/_0880_ ),
    .C(\hash/CA2/_0882_ ),
    .Y(\hash/CA2/_0057_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1447_  (.A(\hash/CA2/_0056_ ),
    .B(\hash/CA2/_0057_ ),
    .Y(\hash/CA2/_0058_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1448_  (.A1(\hash/CA2/_0881_ ),
    .A2(\hash/CA2/_0880_ ),
    .B1(\hash/CA2/_0883_ ),
    .X(\hash/CA2/_0059_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA2/_1449_  (.A(\hash/CA2/_0882_ ),
    .B(\hash/CA2/_0059_ ),
    .X(\hash/CA2/_0060_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA2/_1450_  (.A1(\hash/CA2/_0885_ ),
    .A2(\hash/CA2/_0058_ ),
    .A3(\hash/CA2/_0060_ ),
    .B1(\hash/CA2/_0884_ ),
    .Y(\hash/CA2/_0061_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1451_  (.A(\hash/CA2/_0887_ ),
    .B(\hash/CA2/_0061_ ),
    .Y(\hash/b_new[8] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1452_  (.A(\hash/b_cap[8] ),
    .B(\hash/a_cap[8] ),
    .C(\hash/b_new[8] ),
    .X(\hash/CA2/_0062_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1453_  (.A(\hash/CA2/_0062_ ),
    .Y(\hash/CA2/_0680_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1454_  (.A(\hash/CA2/_0887_ ),
    .Y(\hash/CA2/_0063_ ));
 sky130_fd_sc_hd__or4_1 \hash/CA2/_1455_  (.A(\hash/CA2/_0879_ ),
    .B(\hash/CA2/_0878_ ),
    .C(\hash/CA2/_0880_ ),
    .D(\hash/CA2/_0882_ ),
    .X(\hash/CA2/_0064_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA2/_1456_  (.A1(\hash/CA2/_0882_ ),
    .A2(\hash/CA2/_0059_ ),
    .B1(\hash/CA2/_0064_ ),
    .Y(\hash/CA2/_0065_ ));
 sky130_fd_sc_hd__nor4_1 \hash/CA2/_1457_  (.A(\hash/CA2/_0876_ ),
    .B(\hash/CA2/_0878_ ),
    .C(\hash/CA2/_0880_ ),
    .D(\hash/CA2/_0882_ ),
    .Y(\hash/CA2/_0066_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA2/_1458_  (.A1(\hash/CA2/_0046_ ),
    .A2(\hash/CA2/_0047_ ),
    .B1(\hash/CA2/_0066_ ),
    .Y(\hash/CA2/_0067_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1459_  (.A(\hash/CA2/_0065_ ),
    .B_N(\hash/CA2/_0067_ ),
    .Y(\hash/CA2/_0068_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1460_  (.A1(\hash/CA2/_0885_ ),
    .A2(\hash/CA2/_0068_ ),
    .B1(\hash/CA2/_0884_ ),
    .Y(\hash/CA2/_0069_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1461_  (.A1(\hash/CA2/_0063_ ),
    .A2(\hash/CA2/_0069_ ),
    .B1_N(\hash/CA2/_0886_ ),
    .Y(\hash/CA2/_0070_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1462_  (.A(\hash/CA2/_0889_ ),
    .B(\hash/CA2/_0070_ ),
    .X(\hash/b_new[9] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1463_  (.A(\hash/b_cap[9] ),
    .B(\hash/a_cap[9] ),
    .C(\hash/b_new[9] ),
    .X(\hash/CA2/_0071_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1464_  (.A(\hash/CA2/_0071_ ),
    .Y(\hash/CA2/_0690_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA2/_1465_  (.A(\hash/CA2/_0885_ ),
    .B(\hash/CA2/_0887_ ),
    .C(\hash/CA2/_0889_ ),
    .D(\hash/CA2/_0060_ ),
    .Y(\hash/CA2/_0072_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1466_  (.A1(\hash/CA2/_0056_ ),
    .A2(\hash/CA2/_0057_ ),
    .B1(\hash/CA2/_0072_ ),
    .X(\hash/CA2/_0073_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1467_  (.A1(\hash/CA2/_0887_ ),
    .A2(\hash/CA2/_0884_ ),
    .B1(\hash/CA2/_0886_ ),
    .X(\hash/CA2/_0074_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1468_  (.A1(\hash/CA2/_0889_ ),
    .A2(\hash/CA2/_0074_ ),
    .B1(\hash/CA2/_0888_ ),
    .Y(\hash/CA2/_0075_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1469_  (.A(\hash/CA2/_0073_ ),
    .B(\hash/CA2/_0075_ ),
    .Y(\hash/CA2/_0076_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1470_  (.A(\hash/CA2/_0891_ ),
    .B(\hash/CA2/_0076_ ),
    .X(\hash/b_new[10] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1471_  (.A(\hash/b_cap[10] ),
    .B(\hash/a_cap[10] ),
    .C(\hash/b_new[10] ),
    .X(\hash/CA2/_0077_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1472_  (.A(\hash/CA2/_0077_ ),
    .Y(\hash/CA2/_0698_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1473_  (.A1(\hash/CA2/_0891_ ),
    .A2(\hash/CA2/_0888_ ),
    .B1(\hash/CA2/_0890_ ),
    .X(\hash/CA2/_0078_ ));
 sky130_fd_sc_hd__a31o_2 \hash/CA2/_1474_  (.A1(\hash/CA2/_0889_ ),
    .A2(\hash/CA2/_0891_ ),
    .A3(\hash/CA2/_0074_ ),
    .B1(\hash/CA2/_0078_ ),
    .X(\hash/CA2/_0079_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1475_  (.A1(\hash/CA2/_0885_ ),
    .A2(\hash/CA2/_0884_ ),
    .B1(\hash/CA2/_0887_ ),
    .X(\hash/CA2/_0080_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA2/_1476_  (.A1(\hash/CA2/_0886_ ),
    .A2(\hash/CA2/_0080_ ),
    .B1(\hash/CA2/_0889_ ),
    .C1(\hash/CA2/_0891_ ),
    .Y(\hash/CA2/_0081_ ));
 sky130_fd_sc_hd__nor3b_1 \hash/CA2/_1477_  (.A(\hash/CA2/_0065_ ),
    .B(\hash/CA2/_0081_ ),
    .C_N(\hash/CA2/_0067_ ),
    .Y(\hash/CA2/_0082_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1478_  (.A(\hash/CA2/_0079_ ),
    .B(\hash/CA2/_0082_ ),
    .Y(\hash/CA2/_0083_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1479_  (.A(\hash/CA2/_0893_ ),
    .B(\hash/CA2/_0083_ ),
    .Y(\hash/b_new[11] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1480_  (.A(\hash/b_cap[11] ),
    .B(\hash/a_cap[11] ),
    .C(\hash/b_new[11] ),
    .X(\hash/CA2/_0084_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1481_  (.A(\hash/CA2/_0084_ ),
    .Y(\hash/CA2/_0706_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1482_  (.A1(\hash/CA2/_0891_ ),
    .A2(\hash/CA2/_0076_ ),
    .B1(\hash/CA2/_0890_ ),
    .X(\hash/CA2/_0085_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1483_  (.A1(\hash/CA2/_0893_ ),
    .A2(\hash/CA2/_0085_ ),
    .B1(\hash/CA2/_0892_ ),
    .Y(\hash/CA2/_0086_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1484_  (.A(\hash/CA2/_0895_ ),
    .B(\hash/CA2/_0086_ ),
    .Y(\hash/b_new[12] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1485_  (.A(\hash/b_cap[12] ),
    .B(\hash/a_cap[12] ),
    .C(\hash/b_new[12] ),
    .X(\hash/CA2/_0087_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1486_  (.A(\hash/CA2/_0087_ ),
    .Y(\hash/CA2/_0714_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1487_  (.A(\hash/CA2/_0893_ ),
    .Y(\hash/CA2/_0088_ ));
 sky130_fd_sc_hd__nor4b_1 \hash/CA2/_1488_  (.A(\hash/CA2/_0088_ ),
    .B(\hash/CA2/_0065_ ),
    .C(\hash/CA2/_0081_ ),
    .D_N(\hash/CA2/_0067_ ),
    .Y(\hash/CA2/_0089_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1489_  (.A1(\hash/CA2/_0893_ ),
    .A2(\hash/CA2/_0079_ ),
    .B1(\hash/CA2/_0892_ ),
    .X(\hash/CA2/_0090_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1490_  (.A1(\hash/CA2/_0089_ ),
    .A2(\hash/CA2/_0090_ ),
    .B1(\hash/CA2/_0895_ ),
    .X(\hash/CA2/_0091_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1491_  (.A(\hash/CA2/_0894_ ),
    .B(\hash/CA2/_0091_ ),
    .Y(\hash/CA2/_0092_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1492_  (.A(\hash/CA2/_0092_ ),
    .B_N(\hash/CA2/_0897_ ),
    .Y(\hash/CA2/_0093_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1493_  (.A(\hash/CA2/_0897_ ),
    .B(\hash/CA2/_0894_ ),
    .C(\hash/CA2/_0091_ ),
    .Y(\hash/CA2/_0094_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1494_  (.A(\hash/CA2/_0093_ ),
    .B(\hash/CA2/_0094_ ),
    .Y(\hash/b_new[13] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1495_  (.A(\hash/b_cap[13] ),
    .B(\hash/a_cap[13] ),
    .C(\hash/b_new[13] ),
    .X(\hash/CA2/_0095_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1496_  (.A(\hash/CA2/_0095_ ),
    .Y(\hash/CA2/_0722_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1497_  (.A1(\hash/CA2/_0893_ ),
    .A2(\hash/CA2/_0890_ ),
    .B1(\hash/CA2/_0892_ ),
    .X(\hash/CA2/_0096_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1498_  (.A1(\hash/CA2/_0895_ ),
    .A2(\hash/CA2/_0096_ ),
    .B1(\hash/CA2/_0894_ ),
    .X(\hash/CA2/_0097_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1499_  (.A1(\hash/CA2/_0897_ ),
    .A2(\hash/CA2/_0097_ ),
    .B1(\hash/CA2/_0896_ ),
    .Y(\hash/CA2/_0098_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_1500_  (.A(\hash/CA2/_0075_ ),
    .B(\hash/CA2/_0098_ ),
    .X(\hash/CA2/_0099_ ));
 sky130_fd_sc_hd__o211a_1 \hash/CA2/_1501_  (.A1(\hash/CA2/_0895_ ),
    .A2(\hash/CA2/_0894_ ),
    .B1(\hash/CA2/_0897_ ),
    .C1(\hash/CA2/_0893_ ),
    .X(\hash/CA2/_0100_ ));
 sky130_fd_sc_hd__a21boi_1 \hash/CA2/_1502_  (.A1(\hash/CA2/_0891_ ),
    .A2(\hash/CA2/_0100_ ),
    .B1_N(\hash/CA2/_0098_ ),
    .Y(\hash/CA2/_0101_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1503_  (.A1(\hash/CA2/_0073_ ),
    .A2(\hash/CA2/_0099_ ),
    .B1(\hash/CA2/_0101_ ),
    .X(\hash/CA2/_0102_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1504_  (.A(\hash/CA2/_0899_ ),
    .B(\hash/CA2/_0102_ ),
    .Y(\hash/b_new[14] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1505_  (.A(\hash/b_cap[14] ),
    .B(\hash/a_cap[14] ),
    .C(\hash/b_new[14] ),
    .X(\hash/CA2/_0103_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1506_  (.A(\hash/CA2/_0103_ ),
    .Y(\hash/CA2/_0730_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1507_  (.A(\hash/b_cap[15] ),
    .Y(\hash/CA2/_0104_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1508_  (.A(\hash/a_cap[15] ),
    .Y(\hash/CA2/_0105_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1509_  (.A1(\hash/CA2/_0896_ ),
    .A2(\hash/CA2/_0093_ ),
    .B1(\hash/CA2/_0899_ ),
    .Y(\hash/CA2/_0106_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1510_  (.A_N(\hash/CA2/_0898_ ),
    .B(\hash/CA2/_0106_ ),
    .Y(\hash/CA2/_0107_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1511_  (.A(\hash/CA2/_0901_ ),
    .B(\hash/CA2/_0107_ ),
    .Y(\hash/CA2/_0108_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1512_  (.A(\hash/CA2/_0104_ ),
    .B(\hash/CA2/_0105_ ),
    .C(\hash/CA2/_0108_ ),
    .X(\hash/CA2/_0738_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1513_  (.A1(\hash/CA2/_0073_ ),
    .A2(\hash/CA2/_0099_ ),
    .B1(\hash/CA2/_0101_ ),
    .Y(\hash/CA2/_0109_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1514_  (.A1(\hash/CA2/_0899_ ),
    .A2(\hash/CA2/_0109_ ),
    .B1(\hash/CA2/_0898_ ),
    .X(\hash/CA2/_0110_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1515_  (.A1(\hash/CA2/_0901_ ),
    .A2(\hash/CA2/_0110_ ),
    .B1(\hash/CA2/_0900_ ),
    .Y(\hash/CA2/_0111_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1516_  (.A(\hash/CA2/_0903_ ),
    .B(\hash/CA2/_0111_ ),
    .Y(\hash/b_new[16] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1517_  (.A(\hash/b_cap[16] ),
    .B(\hash/a_cap[16] ),
    .C(\hash/b_new[16] ),
    .X(\hash/CA2/_0112_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1518_  (.A(\hash/CA2/_0112_ ),
    .Y(\hash/CA2/_0746_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1519_  (.A1(\hash/CA2/_0901_ ),
    .A2(\hash/CA2/_0900_ ),
    .B1(\hash/CA2/_0903_ ),
    .X(\hash/CA2/_0113_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1520_  (.A(\hash/CA2/_0899_ ),
    .B(\hash/CA2/_0896_ ),
    .Y(\hash/CA2/_0114_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1521_  (.A(\hash/CA2/_0903_ ),
    .B(\hash/CA2/_0900_ ),
    .Y(\hash/CA2/_0115_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1522_  (.A(\hash/CA2/_0898_ ),
    .B(\hash/CA2/_0902_ ),
    .Y(\hash/CA2/_0116_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1523_  (.A(\hash/CA2/_0114_ ),
    .B(\hash/CA2/_0115_ ),
    .C(\hash/CA2/_0116_ ),
    .Y(\hash/CA2/_0117_ ));
 sky130_fd_sc_hd__and3b_1 \hash/CA2/_1524_  (.A_N(\hash/CA2/_0092_ ),
    .B(\hash/CA2/_0899_ ),
    .C(\hash/CA2/_0897_ ),
    .X(\hash/CA2/_0118_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA2/_1525_  (.A1(\hash/CA2/_0902_ ),
    .A2(\hash/CA2/_0113_ ),
    .B1(\hash/CA2/_0117_ ),
    .B2(\hash/CA2/_0118_ ),
    .Y(\hash/CA2/_0119_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1526_  (.A(\hash/CA2/_0905_ ),
    .B(\hash/CA2/_0119_ ),
    .Y(\hash/b_new[17] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1527_  (.A(\hash/b_cap[17] ),
    .B(\hash/a_cap[17] ),
    .C(\hash/b_new[17] ),
    .X(\hash/CA2/_0120_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1528_  (.A(\hash/CA2/_0120_ ),
    .Y(\hash/CA2/_0755_ ));
 sky130_fd_sc_hd__nand4_1 \hash/CA2/_1530_  (.A(\hash/CA2/_0899_ ),
    .B(\hash/CA2/_0901_ ),
    .C(\hash/CA2/_0903_ ),
    .D(\hash/CA2/_0905_ ),
    .Y(\hash/CA2/_0122_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1531_  (.A1(\hash/CA2/_0901_ ),
    .A2(\hash/CA2/_0898_ ),
    .B1(\hash/CA2/_0900_ ),
    .X(\hash/CA2/_0123_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1532_  (.A1(\hash/CA2/_0903_ ),
    .A2(\hash/CA2/_0123_ ),
    .B1(\hash/CA2/_0902_ ),
    .X(\hash/CA2/_0124_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1533_  (.A1(\hash/CA2/_0905_ ),
    .A2(\hash/CA2/_0124_ ),
    .B1(\hash/CA2/_0904_ ),
    .Y(\hash/CA2/_0125_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1534_  (.A1(\hash/CA2/_0102_ ),
    .A2(\hash/CA2/_0122_ ),
    .B1(\hash/CA2/_0125_ ),
    .Y(\hash/CA2/_0126_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1535_  (.A(\hash/CA2/_0907_ ),
    .B(\hash/CA2/_0126_ ),
    .X(\hash/b_new[18] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1536_  (.A(\hash/b_cap[18] ),
    .B(\hash/a_cap[18] ),
    .C(\hash/b_new[18] ),
    .X(\hash/CA2/_0127_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1537_  (.A(\hash/CA2/_0127_ ),
    .Y(\hash/CA2/_0763_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1538_  (.A(\hash/b_cap[19] ),
    .Y(\hash/CA2/_0128_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1539_  (.A(\hash/a_cap[19] ),
    .Y(\hash/CA2/_0129_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_1541_  (.A(\hash/CA2/_0114_ ),
    .B(\hash/CA2/_0115_ ),
    .C(\hash/CA2/_0116_ ),
    .X(\hash/CA2/_0131_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1542_  (.A(\hash/CA2/_0897_ ),
    .B(\hash/CA2/_0899_ ),
    .Y(\hash/CA2/_0132_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1543_  (.A1(\hash/CA2/_0902_ ),
    .A2(\hash/CA2/_0113_ ),
    .B1(\hash/CA2/_0905_ ),
    .Y(\hash/CA2/_0133_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1544_  (.A1(\hash/CA2/_0131_ ),
    .A2(\hash/CA2/_0132_ ),
    .B1(\hash/CA2/_0133_ ),
    .X(\hash/CA2/_0134_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1545_  (.A1(\hash/CA2/_0092_ ),
    .A2(\hash/CA2/_0131_ ),
    .B1(\hash/CA2/_0134_ ),
    .Y(\hash/CA2/_0135_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1546_  (.A1(\hash/CA2/_0904_ ),
    .A2(\hash/CA2/_0135_ ),
    .B1(\hash/CA2/_0907_ ),
    .Y(\hash/CA2/_0136_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1547_  (.A_N(\hash/CA2/_0906_ ),
    .B(\hash/CA2/_0136_ ),
    .Y(\hash/CA2/_0137_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1548_  (.A(\hash/CA2/_0909_ ),
    .B(\hash/CA2/_0137_ ),
    .Y(\hash/CA2/_0138_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1549_  (.A(\hash/CA2/_0128_ ),
    .B(\hash/CA2/_0129_ ),
    .C(\hash/CA2/_0138_ ),
    .X(\hash/CA2/_0771_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1550_  (.A(\hash/b_cap[20] ),
    .Y(\hash/CA2/_0139_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1551_  (.A(\hash/a_cap[20] ),
    .Y(\hash/CA2/_0140_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1552_  (.A1(\hash/CA2/_0907_ ),
    .A2(\hash/CA2/_0126_ ),
    .B1(\hash/CA2/_0906_ ),
    .X(\hash/CA2/_0141_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1553_  (.A1(\hash/CA2/_0909_ ),
    .A2(\hash/CA2/_0141_ ),
    .B1(\hash/CA2/_0908_ ),
    .X(\hash/CA2/_0142_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1554_  (.A(\hash/CA2/_0911_ ),
    .B(\hash/CA2/_0142_ ),
    .Y(\hash/CA2/_0143_ ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1555_  (.A(\hash/CA2/_0139_ ),
    .B(\hash/CA2/_0140_ ),
    .C(\hash/CA2/_0143_ ),
    .X(\hash/CA2/_0779_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1556_  (.A(\hash/CA2/_0134_ ),
    .Y(\hash/CA2/_0144_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_1557_  (.A(\hash/CA2/_0907_ ),
    .B(\hash/CA2/_0909_ ),
    .C(\hash/CA2/_0911_ ),
    .X(\hash/CA2/_0145_ ));
 sky130_fd_sc_hd__o311ai_0 \hash/CA2/_1558_  (.A1(\hash/CA2/_0894_ ),
    .A2(\hash/CA2/_0091_ ),
    .A3(\hash/CA2/_0117_ ),
    .B1(\hash/CA2/_0144_ ),
    .C1(\hash/CA2/_0145_ ),
    .Y(\hash/CA2/_0146_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1559_  (.A1(\hash/CA2/_0907_ ),
    .A2(\hash/CA2/_0904_ ),
    .B1(\hash/CA2/_0906_ ),
    .X(\hash/CA2/_0147_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1560_  (.A1(\hash/CA2/_0909_ ),
    .A2(\hash/CA2/_0147_ ),
    .B1(\hash/CA2/_0908_ ),
    .X(\hash/CA2/_0148_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1561_  (.A1(\hash/CA2/_0911_ ),
    .A2(\hash/CA2/_0148_ ),
    .B1(\hash/CA2/_0910_ ),
    .Y(\hash/CA2/_0149_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1562_  (.A(\hash/CA2/_0146_ ),
    .B(\hash/CA2/_0149_ ),
    .Y(\hash/CA2/_0150_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1563_  (.A(\hash/CA2/_0913_ ),
    .B(\hash/CA2/_0150_ ),
    .X(\hash/b_new[21] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1564_  (.A(\hash/b_cap[21] ),
    .B(\hash/a_cap[21] ),
    .C(\hash/b_new[21] ),
    .X(\hash/CA2/_0151_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1565_  (.A(\hash/CA2/_0151_ ),
    .Y(\hash/CA2/_0787_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1567_  (.A(\hash/CA2/_0907_ ),
    .B(\hash/CA2/_0909_ ),
    .Y(\hash/CA2/_0153_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1568_  (.A(\hash/CA2/_0911_ ),
    .B(\hash/CA2/_0913_ ),
    .Y(\hash/CA2/_0154_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1569_  (.A(\hash/CA2/_0122_ ),
    .B(\hash/CA2/_0153_ ),
    .C(\hash/CA2/_0154_ ),
    .Y(\hash/CA2/_0155_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_1570_  (.A(\hash/CA2/_0905_ ),
    .B(\hash/CA2/_0907_ ),
    .C(\hash/CA2/_0909_ ),
    .X(\hash/CA2/_0156_ ));
 sky130_fd_sc_hd__a32oi_1 \hash/CA2/_1571_  (.A1(\hash/CA2/_0907_ ),
    .A2(\hash/CA2/_0909_ ),
    .A3(\hash/CA2/_0904_ ),
    .B1(\hash/CA2/_0124_ ),
    .B2(\hash/CA2/_0156_ ),
    .Y(\hash/CA2/_0157_ ));
 sky130_fd_sc_hd__a2111oi_0 \hash/CA2/_1572_  (.A1(\hash/CA2/_0909_ ),
    .A2(\hash/CA2/_0906_ ),
    .B1(\hash/CA2/_0908_ ),
    .C1(\hash/CA2/_0910_ ),
    .D1(\hash/CA2/_0912_ ),
    .Y(\hash/CA2/_0158_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1573_  (.A1(\hash/CA2/_0911_ ),
    .A2(\hash/CA2/_0910_ ),
    .B1(\hash/CA2/_0913_ ),
    .X(\hash/CA2/_0159_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1574_  (.A(\hash/CA2/_0912_ ),
    .B(\hash/CA2/_0159_ ),
    .Y(\hash/CA2/_0160_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1575_  (.A1(\hash/CA2/_0157_ ),
    .A2(\hash/CA2/_0158_ ),
    .B1(\hash/CA2/_0160_ ),
    .Y(\hash/CA2/_0161_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1576_  (.A1(\hash/CA2/_0109_ ),
    .A2(\hash/CA2/_0155_ ),
    .B1(\hash/CA2/_0161_ ),
    .Y(\hash/CA2/_0162_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1577_  (.A(\hash/CA2/_0915_ ),
    .B(\hash/CA2/_0162_ ),
    .Y(\hash/b_new[22] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1578_  (.A(\hash/b_cap[22] ),
    .B(\hash/a_cap[22] ),
    .C(\hash/b_new[22] ),
    .X(\hash/CA2/_0163_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1579_  (.A(\hash/CA2/_0163_ ),
    .Y(\hash/CA2/_0795_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1580_  (.A1(\hash/CA2/_0915_ ),
    .A2(\hash/CA2/_0912_ ),
    .B1(\hash/CA2/_0914_ ),
    .Y(\hash/CA2/_0164_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1581_  (.A(\hash/CA2/_0164_ ),
    .Y(\hash/CA2/_0165_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA2/_1582_  (.A1(\hash/CA2/_0913_ ),
    .A2(\hash/CA2/_0915_ ),
    .A3(\hash/CA2/_0910_ ),
    .B1(\hash/CA2/_0165_ ),
    .Y(\hash/CA2/_0166_ ));
 sky130_fd_sc_hd__or4b_1 \hash/CA2/_1583_  (.A(\hash/CA2/_0894_ ),
    .B(\hash/CA2/_0117_ ),
    .C(\hash/CA2/_0148_ ),
    .D_N(\hash/CA2/_0166_ ),
    .X(\hash/CA2/_0167_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1584_  (.A1(\hash/CA2/_0131_ ),
    .A2(\hash/CA2/_0132_ ),
    .B1(\hash/CA2/_0133_ ),
    .C1(\hash/CA2/_0153_ ),
    .Y(\hash/CA2/_0168_ ));
 sky130_fd_sc_hd__o2111ai_1 \hash/CA2/_1585_  (.A1(\hash/CA2/_0148_ ),
    .A2(\hash/CA2/_0168_ ),
    .B1(\hash/CA2/_0911_ ),
    .C1(\hash/CA2/_0913_ ),
    .D1(\hash/CA2/_0915_ ),
    .Y(\hash/CA2/_0169_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \hash/CA2/_1586_  (.A1_N(\hash/CA2/_0091_ ),
    .A2_N(\hash/CA2/_0167_ ),
    .B1(\hash/CA2/_0169_ ),
    .B2(\hash/CA2/_0166_ ),
    .Y(\hash/CA2/_0170_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1587_  (.A(\hash/CA2/_0917_ ),
    .B(\hash/CA2/_0170_ ),
    .X(\hash/b_new[23] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1588_  (.A(\hash/b_cap[23] ),
    .B(\hash/a_cap[23] ),
    .C(\hash/b_new[23] ),
    .X(\hash/CA2/_0171_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1589_  (.A(\hash/CA2/_0171_ ),
    .Y(\hash/CA2/_0803_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1590_  (.A(\hash/CA2/_0915_ ),
    .B(\hash/CA2/_0155_ ),
    .Y(\hash/CA2/_0172_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1591_  (.A1(\hash/CA2/_0073_ ),
    .A2(\hash/CA2/_0099_ ),
    .B1(\hash/CA2/_0101_ ),
    .C1(\hash/CA2/_0172_ ),
    .Y(\hash/CA2/_0173_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1592_  (.A1(\hash/CA2/_0915_ ),
    .A2(\hash/CA2/_0161_ ),
    .B1(\hash/CA2/_0914_ ),
    .X(\hash/CA2/_0174_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1593_  (.A1(\hash/CA2/_0173_ ),
    .A2(\hash/CA2/_0174_ ),
    .B1(\hash/CA2/_0917_ ),
    .Y(\hash/CA2/_0175_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1594_  (.A_N(\hash/CA2/_0916_ ),
    .B(\hash/CA2/_0175_ ),
    .Y(\hash/CA2/_0176_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1595_  (.A(\hash/CA2/_0919_ ),
    .B(\hash/CA2/_0176_ ),
    .X(\hash/b_new[24] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1596_  (.A1(\hash/a_cap[24] ),
    .A2(\hash/b_new[24] ),
    .B1(\hash/b_cap[24] ),
    .X(\hash/CA2/_0177_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1597_  (.A1(\hash/a_cap[24] ),
    .A2(\hash/b_new[24] ),
    .B1(\hash/CA2/_0177_ ),
    .Y(\hash/CA2/_0811_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1598_  (.A1(\hash/CA2/_0919_ ),
    .A2(\hash/CA2/_0916_ ),
    .B1(\hash/CA2/_0918_ ),
    .X(\hash/CA2/_0178_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1599_  (.A1(\hash/CA2/_0917_ ),
    .A2(\hash/CA2/_0919_ ),
    .B1(\hash/CA2/_0921_ ),
    .X(\hash/CA2/_0179_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1600_  (.A(\hash/CA2/_0917_ ),
    .B(\hash/CA2/_0919_ ),
    .C(\hash/CA2/_0921_ ),
    .Y(\hash/CA2/_0180_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA2/_1601_  (.A1(\hash/CA2/_0178_ ),
    .A2(\hash/CA2/_0179_ ),
    .B1(\hash/CA2/_0180_ ),
    .B2(\hash/CA2/_0164_ ),
    .Y(\hash/CA2/_0181_ ));
 sky130_fd_sc_hd__or3_1 \hash/CA2/_1602_  (.A(\hash/CA2/_0921_ ),
    .B(\hash/CA2/_0165_ ),
    .C(\hash/CA2/_0178_ ),
    .X(\hash/CA2/_0182_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1603_  (.A(\hash/CA2/_0913_ ),
    .B(\hash/CA2/_0915_ ),
    .Y(\hash/CA2/_0183_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1604_  (.A1(\hash/CA2/_0146_ ),
    .A2(\hash/CA2/_0149_ ),
    .B1(\hash/CA2/_0183_ ),
    .Y(\hash/CA2/_0184_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA2/_1605_  (.A0(\hash/CA2/_0182_ ),
    .A1(\hash/CA2/_0180_ ),
    .S(\hash/CA2/_0184_ ),
    .Y(\hash/CA2/_0185_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1606_  (.A1(\hash/CA2/_0921_ ),
    .A2(\hash/CA2/_0178_ ),
    .B1(\hash/CA2/_0181_ ),
    .C1(\hash/CA2/_0185_ ),
    .Y(\hash/b_new[25] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1607_  (.A1(\hash/b_cap[25] ),
    .A2(\hash/a_cap[25] ),
    .B1(\hash/b_new[25] ),
    .X(\hash/CA2/_0186_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1608_  (.A1(\hash/b_cap[25] ),
    .A2(\hash/a_cap[25] ),
    .B1(\hash/CA2/_0186_ ),
    .Y(\hash/CA2/_0819_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1609_  (.A(\hash/CA2/_0923_ ),
    .Y(\hash/CA2/_0187_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1610_  (.A(\hash/CA2/_0173_ ),
    .B(\hash/CA2/_0174_ ),
    .Y(\hash/CA2/_0188_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1611_  (.A(\hash/CA2/_0916_ ),
    .B(\hash/CA2/_0918_ ),
    .C(\hash/CA2/_0920_ ),
    .Y(\hash/CA2/_0189_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1612_  (.A1(\hash/CA2/_0917_ ),
    .A2(\hash/CA2/_0916_ ),
    .B1(\hash/CA2/_0919_ ),
    .Y(\hash/CA2/_0190_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1613_  (.A_N(\hash/CA2/_0918_ ),
    .B(\hash/CA2/_0190_ ),
    .Y(\hash/CA2/_0191_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1614_  (.A1(\hash/CA2/_0921_ ),
    .A2(\hash/CA2/_0191_ ),
    .B1(\hash/CA2/_0920_ ),
    .Y(\hash/CA2/_0192_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1615_  (.A1(\hash/CA2/_0188_ ),
    .A2(\hash/CA2/_0189_ ),
    .B1(\hash/CA2/_0192_ ),
    .Y(\hash/CA2/_0193_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1616_  (.A(\hash/CA2/_0187_ ),
    .B(\hash/CA2/_0193_ ),
    .Y(\hash/b_new[26] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1617_  (.A(\hash/b_cap[26] ),
    .B(\hash/a_cap[26] ),
    .C(\hash/b_new[26] ),
    .X(\hash/CA2/_0194_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1618_  (.A(\hash/CA2/_0194_ ),
    .Y(\hash/CA2/_0827_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1619_  (.A(\hash/CA2/_0187_ ),
    .B(\hash/CA2/_0180_ ),
    .Y(\hash/CA2/_0195_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1620_  (.A1(\hash/CA2/_0921_ ),
    .A2(\hash/CA2/_0178_ ),
    .B1(\hash/CA2/_0920_ ),
    .Y(\hash/CA2/_0196_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1621_  (.A(\hash/CA2/_0187_ ),
    .B(\hash/CA2/_0196_ ),
    .Y(\hash/CA2/_0197_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1622_  (.A(\hash/CA2/_0922_ ),
    .B(\hash/CA2/_0197_ ),
    .Y(\hash/CA2/_0198_ ));
 sky130_fd_sc_hd__a21boi_1 \hash/CA2/_1623_  (.A1(\hash/CA2/_0170_ ),
    .A2(\hash/CA2/_0195_ ),
    .B1_N(\hash/CA2/_0198_ ),
    .Y(\hash/CA2/_0199_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1624_  (.A(\hash/CA2/_0925_ ),
    .B(\hash/CA2/_0199_ ),
    .Y(\hash/b_new[27] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1625_  (.A(\hash/b_cap[27] ),
    .B(\hash/a_cap[27] ),
    .C(\hash/b_new[27] ),
    .X(\hash/CA2/_0200_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1626_  (.A(\hash/CA2/_0200_ ),
    .Y(\hash/CA2/_0835_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1627_  (.A(\hash/a_cap[28] ),
    .B(\hash/CA2/_0925_ ),
    .Y(\hash/CA2/_0201_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1628_  (.A(\hash/b_cap[28] ),
    .B(\hash/CA2/_0925_ ),
    .Y(\hash/CA2/_0202_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1629_  (.A1(\hash/CA2/_0923_ ),
    .A2(\hash/CA2/_0193_ ),
    .B1(\hash/CA2/_0922_ ),
    .Y(\hash/CA2/_0203_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1630_  (.A1(\hash/CA2/_0201_ ),
    .A2(\hash/CA2/_0202_ ),
    .B1(\hash/CA2/_0927_ ),
    .C1(\hash/CA2/_0203_ ),
    .Y(\hash/CA2/_0204_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1631_  (.A(\hash/CA2/_0924_ ),
    .Y(\hash/CA2/_0205_ ));
 sky130_fd_sc_hd__o2111a_1 \hash/CA2/_1632_  (.A1(\hash/b_cap[28] ),
    .A2(\hash/a_cap[28] ),
    .B1(\hash/CA2/_0927_ ),
    .C1(\hash/CA2/_0205_ ),
    .D1(\hash/CA2/_0203_ ),
    .X(\hash/CA2/_0206_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1633_  (.A(\hash/CA2/_0925_ ),
    .Y(\hash/CA2/_0207_ ));
 sky130_fd_sc_hd__o2111ai_1 \hash/CA2/_1634_  (.A1(\hash/b_cap[28] ),
    .A2(\hash/a_cap[28] ),
    .B1(\hash/CA2/_0207_ ),
    .C1(\hash/CA2/_0927_ ),
    .D1(\hash/CA2/_0205_ ),
    .Y(\hash/CA2/_0208_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1635_  (.A(\hash/CA2/_0927_ ),
    .Y(\hash/CA2/_0209_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA2/_1636_  (.A1(\hash/b_cap[28] ),
    .A2(\hash/a_cap[28] ),
    .B1(\hash/CA2/_0209_ ),
    .C1(\hash/CA2/_0924_ ),
    .Y(\hash/CA2/_0210_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1637_  (.A(\hash/CA2/_0208_ ),
    .B(\hash/CA2/_0210_ ),
    .Y(\hash/CA2/_0211_ ));
 sky130_fd_sc_hd__a2111oi_0 \hash/CA2/_1638_  (.A1(\hash/b_cap[28] ),
    .A2(\hash/a_cap[28] ),
    .B1(\hash/CA2/_0204_ ),
    .C1(\hash/CA2/_0206_ ),
    .D1(\hash/CA2/_0211_ ),
    .Y(\hash/CA2/_0843_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1639_  (.A1(\hash/CA2/_0927_ ),
    .A2(\hash/CA2/_0924_ ),
    .B1(\hash/CA2/_0926_ ),
    .Y(\hash/CA2/_0212_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_1640_  (.A1(\hash/CA2/_0207_ ),
    .A2(\hash/CA2/_0209_ ),
    .A3(\hash/CA2/_0199_ ),
    .B1(\hash/CA2/_0212_ ),
    .Y(\hash/CA2/_0213_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1641_  (.A(\hash/CA2/_0929_ ),
    .B(\hash/CA2/_0213_ ),
    .X(\hash/b_new[29] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1642_  (.A(\hash/b_cap[29] ),
    .B(\hash/a_cap[29] ),
    .C(\hash/b_new[29] ),
    .X(\hash/CA2/_0214_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1643_  (.A(\hash/CA2/_0214_ ),
    .Y(\hash/CA2/_0852_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1644_  (.A(\hash/p1_cap[1] ),
    .Y(\hash/CA2/_0610_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1645_  (.A(\hash/p4_cap[0] ),
    .Y(\hash/CA2/_0619_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1646_  (.A(\hash/p4_cap[1] ),
    .Y(\hash/CA2/_0624_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1647_  (.A(\hash/p4_cap[2] ),
    .Y(\hash/CA2/_0632_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1648_  (.A(\hash/p4_cap[3] ),
    .Y(\hash/CA2/_0641_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1649_  (.A(\hash/p4_cap[4] ),
    .Y(\hash/CA2/_0650_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1650_  (.A(\hash/p4_cap[8] ),
    .Y(\hash/CA2/_0678_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1651_  (.A(\hash/p4_cap[9] ),
    .Y(\hash/CA2/_0688_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1652_  (.A(\hash/p4_cap[10] ),
    .Y(\hash/CA2/_0696_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1653_  (.A(\hash/p4_cap[11] ),
    .Y(\hash/CA2/_0704_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1654_  (.A(\hash/p4_cap[12] ),
    .Y(\hash/CA2/_0712_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1655_  (.A(\hash/p4_cap[13] ),
    .Y(\hash/CA2/_0720_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1656_  (.A(\hash/p4_cap[14] ),
    .Y(\hash/CA2/_0728_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1657_  (.A(\hash/p4_cap[15] ),
    .Y(\hash/CA2/_0736_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1658_  (.A(\hash/p4_cap[16] ),
    .Y(\hash/CA2/_0744_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1659_  (.A(\hash/p4_cap[17] ),
    .Y(\hash/CA2/_0753_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1660_  (.A(\hash/p4_cap[18] ),
    .Y(\hash/CA2/_0761_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1661_  (.A(\hash/p4_cap[19] ),
    .Y(\hash/CA2/_0769_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1662_  (.A(\hash/p4_cap[20] ),
    .Y(\hash/CA2/_0777_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1663_  (.A(\hash/p4_cap[21] ),
    .Y(\hash/CA2/_0785_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1664_  (.A(\hash/p4_cap[22] ),
    .Y(\hash/CA2/_0793_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1665_  (.A(\hash/p4_cap[23] ),
    .Y(\hash/CA2/_0801_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1666_  (.A(\hash/p4_cap[24] ),
    .Y(\hash/CA2/_0809_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1667_  (.A(\hash/p4_cap[25] ),
    .Y(\hash/CA2/_0817_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1668_  (.A(\hash/p4_cap[26] ),
    .Y(\hash/CA2/_0825_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1669_  (.A(\hash/p4_cap[27] ),
    .Y(\hash/CA2/_0833_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1670_  (.A(\hash/p4_cap[28] ),
    .Y(\hash/CA2/_0841_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1671_  (.A(\hash/p4_cap[29] ),
    .Y(\hash/CA2/_0850_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1672_  (.A(\hash/CA2/_1213_ ),
    .Y(\hash/CA2/_0866_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1673_  (.A(\hash/p3_cap[1] ),
    .Y(\hash/CA2/_0611_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1674_  (.A(\hash/CA2/s0[0] ),
    .Y(\hash/CA2/_0620_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1675_  (.A(\hash/CA2/s0[1] ),
    .Y(\hash/CA2/_0625_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1676_  (.A(\hash/CA2/s0[2] ),
    .Y(\hash/CA2/_0633_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1677_  (.A(\hash/CA2/s0[3] ),
    .Y(\hash/CA2/_0642_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1678_  (.A(\hash/CA2/s0[4] ),
    .Y(\hash/CA2/_0651_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1679_  (.A(\hash/CA2/s0[8] ),
    .Y(\hash/CA2/_0679_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1680_  (.A(\hash/CA2/s0[9] ),
    .Y(\hash/CA2/_0689_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1681_  (.A(\hash/CA2/s0[10] ),
    .Y(\hash/CA2/_0697_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1682_  (.A(\hash/CA2/s0[11] ),
    .Y(\hash/CA2/_0705_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1683_  (.A(\hash/CA2/s0[12] ),
    .Y(\hash/CA2/_0713_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1684_  (.A(\hash/CA2/s0[13] ),
    .Y(\hash/CA2/_0721_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1685_  (.A(\hash/CA2/s0[14] ),
    .Y(\hash/CA2/_0729_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1686_  (.A(\hash/CA2/s0[15] ),
    .Y(\hash/CA2/_0737_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1687_  (.A(\hash/CA2/s0[16] ),
    .Y(\hash/CA2/_0745_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1688_  (.A(\hash/CA2/s0[17] ),
    .Y(\hash/CA2/_0754_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1689_  (.A(\hash/CA2/s0[18] ),
    .Y(\hash/CA2/_0762_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1690_  (.A(\hash/CA2/s0[19] ),
    .Y(\hash/CA2/_0770_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1691_  (.A(\hash/CA2/s0[20] ),
    .Y(\hash/CA2/_0778_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1692_  (.A(\hash/CA2/s0[21] ),
    .Y(\hash/CA2/_0786_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1693_  (.A(\hash/CA2/s0[22] ),
    .Y(\hash/CA2/_0794_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1694_  (.A(\hash/CA2/s0[23] ),
    .Y(\hash/CA2/_0802_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1695_  (.A(\hash/CA2/s0[24] ),
    .Y(\hash/CA2/_0810_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1696_  (.A(\hash/CA2/s0[25] ),
    .Y(\hash/CA2/_0818_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1697_  (.A(\hash/CA2/s0[26] ),
    .Y(\hash/CA2/_0826_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1698_  (.A(\hash/CA2/s0[27] ),
    .Y(\hash/CA2/_0834_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1699_  (.A(\hash/CA2/s0[28] ),
    .Y(\hash/CA2/_0842_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1700_  (.A(\hash/CA2/s0[29] ),
    .Y(\hash/CA2/_0851_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1701_  (.A(\hash/CA2/_0871_ ),
    .Y(\hash/CA2/_0612_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1702_  (.A(\hash/CA2/_0868_ ),
    .Y(\hash/a_new[2] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1703_  (.A(\hash/CA2/_0618_ ),
    .Y(\hash/CA2/_0629_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1704_  (.A(\hash/CA2/_0673_ ),
    .Y(\hash/CA2/_0683_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1705_  (.A(\hash/CA2/_0630_ ),
    .Y(\hash/CA2/_1101_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1706_  (.A(\hash/CA2/_0638_ ),
    .Y(\hash/CA2/_1105_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1707_  (.A(\hash/CA2/_0647_ ),
    .Y(\hash/CA2/_1109_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1708_  (.A(\hash/CA2/_0653_ ),
    .Y(\hash/CA2/_0662_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1709_  (.A(\hash/CA2/_0656_ ),
    .Y(\hash/CA2/_1113_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1710_  (.A(\hash/CA2/_0685_ ),
    .Y(\hash/CA2/_1123_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1711_  (.A(\hash/CA2/_0694_ ),
    .Y(\hash/CA2/_1127_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1712_  (.A(\hash/CA2/_0702_ ),
    .Y(\hash/CA2/_1131_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1713_  (.A(\hash/CA2/_0710_ ),
    .Y(\hash/CA2/_1135_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1714_  (.A(\hash/CA2/_0718_ ),
    .Y(\hash/CA2/_1139_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1715_  (.A(\hash/CA2/_0726_ ),
    .Y(\hash/CA2/_1143_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1716_  (.A(\hash/CA2/_0734_ ),
    .Y(\hash/CA2/_1147_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1717_  (.A(\hash/CA2/_0742_ ),
    .Y(\hash/CA2/_1151_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1718_  (.A(\hash/CA2/_0750_ ),
    .Y(\hash/CA2/_1155_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1719_  (.A(\hash/CA2/_0759_ ),
    .Y(\hash/CA2/_1159_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1720_  (.A(\hash/CA2/_0767_ ),
    .Y(\hash/CA2/_1163_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1721_  (.A(\hash/CA2/_0775_ ),
    .Y(\hash/CA2/_1167_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1722_  (.A(\hash/CA2/_0783_ ),
    .Y(\hash/CA2/_1171_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1723_  (.A(\hash/CA2/_0791_ ),
    .Y(\hash/CA2/_1175_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1724_  (.A(\hash/CA2/_0799_ ),
    .Y(\hash/CA2/_1179_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1725_  (.A(\hash/CA2/_0807_ ),
    .Y(\hash/CA2/_1183_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1726_  (.A(\hash/CA2/_0815_ ),
    .Y(\hash/CA2/_1187_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1727_  (.A(\hash/CA2/_0823_ ),
    .Y(\hash/CA2/_1191_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1728_  (.A(\hash/CA2/_0831_ ),
    .Y(\hash/CA2/_1195_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1729_  (.A(\hash/CA2/_0839_ ),
    .Y(\hash/CA2/_1199_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1730_  (.A(\hash/CA2/_0847_ ),
    .Y(\hash/CA2/_1203_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1731_  (.A(\hash/CA2/_0853_ ),
    .Y(\hash/CA2/_0862_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1732_  (.A(\hash/CA2/_0856_ ),
    .Y(\hash/CA2/_1207_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1733_  (.A(\hash/CA2/_1070_ ),
    .B(\hash/CA2/_1076_ ),
    .Y(\hash/CA2/_0215_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1734_  (.A(\hash/CA2/_1082_ ),
    .B(\hash/CA2/_1088_ ),
    .Y(\hash/CA2/_0216_ ));
 sky130_fd_sc_hd__a2111oi_0 \hash/CA2/_1735_  (.A1(\hash/CA2/_0007_ ),
    .A2(\hash/CA2/_0021_ ),
    .B1(\hash/CA2/_0023_ ),
    .C1(\hash/CA2/_0215_ ),
    .D1(\hash/CA2/_0216_ ),
    .Y(\hash/CA2/_0217_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1736_  (.A(\hash/CA2/_1076_ ),
    .B(\hash/CA2/_1069_ ),
    .Y(\hash/CA2/_0218_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1737_  (.A(\hash/CA2/_0216_ ),
    .B(\hash/CA2/_0218_ ),
    .Y(\hash/CA2/_0219_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1738_  (.A(\hash/CA2/_1088_ ),
    .Y(\hash/CA2/_0220_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1739_  (.A1(\hash/CA2/_0220_ ),
    .A2(\hash/CA2/_0033_ ),
    .B1_N(\hash/CA2/_1087_ ),
    .Y(\hash/CA2/_0221_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_1740_  (.A1(\hash/CA2/_0217_ ),
    .A2(\hash/CA2/_0219_ ),
    .A3(\hash/CA2/_0221_ ),
    .B1(\hash/CA2/_1093_ ),
    .Y(\hash/CA2/_0222_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1741_  (.A_N(\hash/CA2/_1092_ ),
    .B(\hash/CA2/_0222_ ),
    .Y(\hash/CA2/_0223_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1742_  (.A(\hash/CA2/_1098_ ),
    .B(\hash/CA2/_0223_ ),
    .X(\hash/CA2/_0863_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1743_  (.A(\hash/CA2/_0639_ ),
    .Y(\hash/CA2/_1102_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1744_  (.A(\hash/CA2/_0648_ ),
    .Y(\hash/CA2/_1106_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1745_  (.A(\hash/CA2/_0657_ ),
    .Y(\hash/CA2/_1110_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1746_  (.A1(\hash/CA2/_0876_ ),
    .A2(\hash/CA2/_0048_ ),
    .B1(\hash/CA2/_0879_ ),
    .X(\hash/CA2/_0224_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1747_  (.A(\hash/CA2/_0878_ ),
    .B(\hash/CA2/_0224_ ),
    .Y(\hash/CA2/_0225_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1748_  (.A(\hash/CA2/_0881_ ),
    .B(\hash/CA2/_0225_ ),
    .Y(\hash/b_new[5] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1749_  (.A(\hash/b_cap[5] ),
    .B(\hash/a_cap[5] ),
    .C(\hash/b_new[5] ),
    .X(\hash/CA2/_0659_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1750_  (.A(\hash/CA2/_0537_ ),
    .B(\hash/CA2/_0538_ ),
    .Y(\hash/CA2/_0226_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1751_  (.A(\hash/CA2/_0944_ ),
    .B(\hash/CA2/_0226_ ),
    .Y(\hash/CA2/_0227_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1752_  (.A1(\hash/CA2/_0527_ ),
    .A2(\hash/CA2/_0227_ ),
    .B1_N(\hash/CA2/_0949_ ),
    .Y(\hash/CA2/_0228_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1753_  (.A(\hash/CA2/_0955_ ),
    .B(\hash/CA2/_0228_ ),
    .X(\hash/CA2/_0663_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1754_  (.A_N(\hash/CA2/_0878_ ),
    .B(\hash/CA2/_0056_ ),
    .Y(\hash/CA2/_0229_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1755_  (.A1(\hash/CA2/_0881_ ),
    .A2(\hash/CA2/_0229_ ),
    .B1(\hash/CA2/_0880_ ),
    .Y(\hash/CA2/_0230_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1756_  (.A(\hash/CA2/_0883_ ),
    .B(\hash/CA2/_0230_ ),
    .Y(\hash/b_new[6] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1757_  (.A(\hash/b_cap[6] ),
    .B(\hash/a_cap[6] ),
    .C(\hash/b_new[6] ),
    .X(\hash/CA2/_0666_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1758_  (.A1(\hash/CA2/_0527_ ),
    .A2(\hash/CA2/_0526_ ),
    .B1_N(\hash/CA2/_0949_ ),
    .Y(\hash/CA2/_0231_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1759_  (.A1(\hash/CA2/_0955_ ),
    .A2(\hash/CA2/_0231_ ),
    .B1(\hash/CA2/_0954_ ),
    .Y(\hash/CA2/_0232_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1760_  (.A(\hash/CA2/_0960_ ),
    .B(\hash/CA2/_0232_ ),
    .Y(\hash/CA2/_0669_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1761_  (.A(\hash/CA2/_0885_ ),
    .B(\hash/CA2/_0068_ ),
    .X(\hash/b_new[7] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1762_  (.A(\hash/b_cap[7] ),
    .B(\hash/a_cap[7] ),
    .C(\hash/b_new[7] ),
    .X(\hash/CA2/_0672_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1763_  (.A(\hash/CA2/_0965_ ),
    .B(\hash/CA2/_0541_ ),
    .Y(\hash/CA2/_0675_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1764_  (.A(\hash/CA2/_0686_ ),
    .Y(\hash/CA2/_1120_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1765_  (.A(\hash/CA2/_0695_ ),
    .Y(\hash/CA2/_1124_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1766_  (.A(\hash/CA2/_0703_ ),
    .Y(\hash/CA2/_1128_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1767_  (.A(\hash/CA2/_0711_ ),
    .Y(\hash/CA2/_1132_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1768_  (.A(\hash/CA2/_0719_ ),
    .Y(\hash/CA2/_1136_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1769_  (.A(\hash/CA2/_0727_ ),
    .Y(\hash/CA2/_1140_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1770_  (.A(\hash/CA2/_0735_ ),
    .Y(\hash/CA2/_1144_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1771_  (.A(\hash/CA2/_0743_ ),
    .Y(\hash/CA2/_1148_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1772_  (.A(\hash/CA2/_0751_ ),
    .Y(\hash/CA2/_1152_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1773_  (.A(\hash/CA2/_0760_ ),
    .Y(\hash/CA2/_1156_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1774_  (.A(\hash/CA2/_0768_ ),
    .Y(\hash/CA2/_1160_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1775_  (.A(\hash/CA2/_0776_ ),
    .Y(\hash/CA2/_1164_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1776_  (.A(\hash/CA2/_0784_ ),
    .Y(\hash/CA2/_1168_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1777_  (.A(\hash/CA2/_0792_ ),
    .Y(\hash/CA2/_1172_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1778_  (.A(\hash/CA2/_0800_ ),
    .Y(\hash/CA2/_1176_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1779_  (.A(\hash/CA2/_0808_ ),
    .Y(\hash/CA2/_1180_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1780_  (.A(\hash/CA2/_0816_ ),
    .Y(\hash/CA2/_1184_ ));
 sky130_fd_sc_hd__or2_2 \hash/CA2/_1781_  (.A(\hash/CA2/_0017_ ),
    .B(\hash/CA2/_0020_ ),
    .X(\hash/CA2/_1071_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1782_  (.A(\hash/CA2/_0824_ ),
    .Y(\hash/CA2/_1188_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1783_  (.A(\hash/CA2/_0832_ ),
    .Y(\hash/CA2/_1192_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1784_  (.A(\hash/CA2/_0840_ ),
    .Y(\hash/CA2/_1196_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1785_  (.A(\hash/CA2/_0220_ ),
    .B(\hash/CA2/_0034_ ),
    .Y(\hash/CA2/_0849_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1786_  (.A(\hash/CA2/_0848_ ),
    .Y(\hash/CA2/_1200_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1787_  (.A(\hash/CA2/_0857_ ),
    .Y(\hash/CA2/_1204_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1788_  (.A1(\hash/CA2/_0927_ ),
    .A2(\hash/CA2/_0926_ ),
    .B1(\hash/CA2/_0929_ ),
    .Y(\hash/CA2/_0233_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1789_  (.A(\hash/CA2/_0187_ ),
    .B(\hash/CA2/_0207_ ),
    .C(\hash/CA2/_0233_ ),
    .Y(\hash/CA2/_0234_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1790_  (.A(\hash/CA2/_0924_ ),
    .B(\hash/CA2/_0926_ ),
    .Y(\hash/CA2/_0235_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1791_  (.A(\hash/CA2/_0925_ ),
    .B(\hash/CA2/_0922_ ),
    .Y(\hash/CA2/_0236_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1792_  (.A1(\hash/CA2/_0235_ ),
    .A2(\hash/CA2/_0236_ ),
    .B1(\hash/CA2/_0233_ ),
    .Y(\hash/CA2/_0237_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1793_  (.A1(\hash/CA2/_0193_ ),
    .A2(\hash/CA2/_0234_ ),
    .B1(\hash/CA2/_0237_ ),
    .C1(\hash/CA2/_0928_ ),
    .Y(\hash/CA2/_0238_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1794_  (.A(\hash/CA2/_0931_ ),
    .B(\hash/CA2/_0238_ ),
    .Y(\hash/b_new[30] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1795_  (.A(\hash/b_cap[30] ),
    .B(\hash/a_cap[30] ),
    .C(\hash/b_new[30] ),
    .X(\hash/CA2/_0859_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1796_  (.A(\hash/CA2/_0623_ ),
    .Y(\hash/CA2/_1210_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1797_  (.A(\hash/CA2/_0631_ ),
    .Y(\hash/CA2/_1212_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1798_  (.A(\hash/CA2/_1112_ ),
    .Y(\hash/CA2/_0239_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1799_  (.A1(\hash/CA2/_1213_ ),
    .A2(\hash/CA2/_1104_ ),
    .B1(\hash/CA2/_1103_ ),
    .X(\hash/CA2/_0240_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1800_  (.A1(\hash/CA2/_1108_ ),
    .A2(\hash/CA2/_0240_ ),
    .B1(\hash/CA2/_1107_ ),
    .Y(\hash/CA2/_0241_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1801_  (.A(\hash/CA2/_1111_ ),
    .B(\hash/CA2/_1114_ ),
    .Y(\hash/CA2/_0242_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/CA2/_1802_  (.A1(\hash/CA2/_0239_ ),
    .A2(\hash/CA2/_0241_ ),
    .B1(\hash/CA2/_0242_ ),
    .Y(\hash/CA2/_0243_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1803_  (.A1(\hash/CA2/_1115_ ),
    .A2(\hash/CA2/_1114_ ),
    .B1(\hash/CA2/_1117_ ),
    .X(\hash/CA2/_0244_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1804_  (.A1(\hash/CA2/_0243_ ),
    .A2(\hash/CA2/_0244_ ),
    .B1(\hash/CA2/_1116_ ),
    .Y(\hash/CA2/_0245_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1805_  (.A(\hash/CA2/_0245_ ),
    .B_N(\hash/CA2/_1119_ ),
    .Y(\hash/CA2/_0246_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1806_  (.A1(\hash/CA2/_1118_ ),
    .A2(\hash/CA2/_0246_ ),
    .B1(\hash/CA2/_1122_ ),
    .Y(\hash/CA2/_0247_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1807_  (.A_N(\hash/CA2/_1121_ ),
    .B(\hash/CA2/_0247_ ),
    .Y(\hash/CA2/_0248_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1808_  (.A1(\hash/CA2/_1126_ ),
    .A2(\hash/CA2/_0248_ ),
    .B1(\hash/CA2/_1125_ ),
    .Y(\hash/CA2/_0249_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1809_  (.A(\hash/CA2/_1130_ ),
    .B(\hash/CA2/_0249_ ),
    .Y(\hash/a_new[10] ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1810_  (.A(\hash/CA2/_0867_ ),
    .B_N(\hash/CA2/_1108_ ),
    .Y(\hash/CA2/_0250_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1811_  (.A1(\hash/CA2/_1107_ ),
    .A2(\hash/CA2/_0250_ ),
    .B1(\hash/CA2/_1112_ ),
    .X(\hash/CA2/_0251_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1812_  (.A1(\hash/CA2/_1111_ ),
    .A2(\hash/CA2/_0251_ ),
    .B1(\hash/CA2/_1115_ ),
    .Y(\hash/CA2/_0252_ ));
 sky130_fd_sc_hd__nor4_1 \hash/CA2/_1813_  (.A(\hash/CA2/_1114_ ),
    .B(\hash/CA2/_1116_ ),
    .C(\hash/CA2/_1118_ ),
    .D(\hash/CA2/_1121_ ),
    .Y(\hash/CA2/_0253_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1814_  (.A1(\hash/CA2/_1117_ ),
    .A2(\hash/CA2/_1116_ ),
    .B1(\hash/CA2/_1119_ ),
    .Y(\hash/CA2/_0254_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1815_  (.A_N(\hash/CA2/_1118_ ),
    .B(\hash/CA2/_0254_ ),
    .Y(\hash/CA2/_0255_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1816_  (.A1(\hash/CA2/_1122_ ),
    .A2(\hash/CA2/_0255_ ),
    .B1(\hash/CA2/_1121_ ),
    .Y(\hash/CA2/_0256_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1817_  (.A1(\hash/CA2/_0252_ ),
    .A2(\hash/CA2/_0253_ ),
    .B1(\hash/CA2/_0256_ ),
    .Y(\hash/CA2/_0257_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1818_  (.A1(\hash/CA2/_1126_ ),
    .A2(\hash/CA2/_0257_ ),
    .B1(\hash/CA2/_1125_ ),
    .X(\hash/CA2/_0258_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1819_  (.A1(\hash/CA2/_1130_ ),
    .A2(\hash/CA2/_0258_ ),
    .B1(\hash/CA2/_1129_ ),
    .X(\hash/CA2/_0259_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1820_  (.A(\hash/CA2/_1134_ ),
    .B(\hash/CA2/_0259_ ),
    .X(\hash/a_new[11] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1821_  (.A(\hash/CA2/_1138_ ),
    .Y(\hash/CA2/_0260_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1822_  (.A(\hash/CA2/_1134_ ),
    .B(\hash/CA2/_1130_ ),
    .Y(\hash/CA2/_0261_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1823_  (.A1(\hash/CA2/_1134_ ),
    .A2(\hash/CA2/_1129_ ),
    .B1(\hash/CA2/_1133_ ),
    .X(\hash/CA2/_0262_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1824_  (.A1(\hash/CA2/_0249_ ),
    .A2(\hash/CA2/_0261_ ),
    .B1_N(\hash/CA2/_0262_ ),
    .Y(\hash/CA2/_0263_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1825_  (.A(\hash/CA2/_0260_ ),
    .B(\hash/CA2/_0263_ ),
    .Y(\hash/a_new[12] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1826_  (.A(\hash/CA2/_1142_ ),
    .Y(\hash/CA2/_0264_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1827_  (.A1(\hash/CA2/_1134_ ),
    .A2(\hash/CA2/_0259_ ),
    .B1(\hash/CA2/_1133_ ),
    .Y(\hash/CA2/_0265_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1828_  (.A1(\hash/CA2/_0260_ ),
    .A2(\hash/CA2/_0265_ ),
    .B1_N(\hash/CA2/_1137_ ),
    .Y(\hash/CA2/_0266_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1829_  (.A(\hash/CA2/_0264_ ),
    .B(\hash/CA2/_0266_ ),
    .Y(\hash/a_new[13] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1830_  (.A(\hash/CA2/_1146_ ),
    .Y(\hash/CA2/_0267_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1831_  (.A(\hash/CA2/_1119_ ),
    .B(\hash/CA2/_1122_ ),
    .C(\hash/CA2/_1126_ ),
    .Y(\hash/CA2/_0268_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1832_  (.A1(\hash/CA2/_1138_ ),
    .A2(\hash/CA2/_0262_ ),
    .B1(\hash/CA2/_1137_ ),
    .Y(\hash/CA2/_0269_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1833_  (.A1(\hash/CA2/_1122_ ),
    .A2(\hash/CA2/_1118_ ),
    .B1(\hash/CA2/_1121_ ),
    .X(\hash/CA2/_0270_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1834_  (.A1(\hash/CA2/_1126_ ),
    .A2(\hash/CA2/_0270_ ),
    .B1(\hash/CA2/_1141_ ),
    .C1(\hash/CA2/_1125_ ),
    .Y(\hash/CA2/_0271_ ));
 sky130_fd_sc_hd__o221a_2 \hash/CA2/_1835_  (.A1(\hash/CA2/_0245_ ),
    .A2(\hash/CA2/_0268_ ),
    .B1(\hash/CA2/_0269_ ),
    .B2(\hash/CA2/_0264_ ),
    .C1(\hash/CA2/_0271_ ),
    .X(\hash/CA2/_0272_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1836_  (.A(\hash/CA2/_1134_ ),
    .B(\hash/CA2/_1130_ ),
    .C(\hash/CA2/_1138_ ),
    .Y(\hash/CA2/_0273_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1837_  (.A(\hash/CA2/_0269_ ),
    .B(\hash/CA2/_0273_ ),
    .Y(\hash/CA2/_0274_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1838_  (.A1(\hash/CA2/_1142_ ),
    .A2(\hash/CA2/_0274_ ),
    .B1(\hash/CA2/_1141_ ),
    .Y(\hash/CA2/_0275_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1839_  (.A(\hash/CA2/_0272_ ),
    .B(\hash/CA2/_0275_ ),
    .Y(\hash/CA2/_0276_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1840_  (.A(\hash/CA2/_0267_ ),
    .B(\hash/CA2/_0276_ ),
    .Y(\hash/a_new[14] ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1841_  (.A(\hash/CA2/_1134_ ),
    .B(\hash/CA2/_1138_ ),
    .C(\hash/CA2/_1142_ ),
    .Y(\hash/CA2/_0277_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1842_  (.A1(\hash/CA2/_1130_ ),
    .A2(\hash/CA2/_1125_ ),
    .B1(\hash/CA2/_1129_ ),
    .Y(\hash/CA2/_0278_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1843_  (.A(\hash/CA2/_1142_ ),
    .B(\hash/CA2/_1126_ ),
    .Y(\hash/CA2/_0279_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1844_  (.A(\hash/CA2/_0273_ ),
    .B(\hash/CA2/_0279_ ),
    .Y(\hash/CA2/_0280_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1845_  (.A(\hash/CA2/_0257_ ),
    .B(\hash/CA2/_0280_ ),
    .Y(\hash/CA2/_0281_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1846_  (.A1(\hash/CA2/_1138_ ),
    .A2(\hash/CA2/_1133_ ),
    .B1(\hash/CA2/_1137_ ),
    .X(\hash/CA2/_0282_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1847_  (.A1(\hash/CA2/_1142_ ),
    .A2(\hash/CA2/_0282_ ),
    .B1(\hash/CA2/_1141_ ),
    .Y(\hash/CA2/_0283_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA2/_1848_  (.A1(\hash/CA2/_0277_ ),
    .A2(\hash/CA2/_0278_ ),
    .B1(\hash/CA2/_0281_ ),
    .C1(\hash/CA2/_0283_ ),
    .Y(\hash/CA2/_0284_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1849_  (.A1(\hash/CA2/_1146_ ),
    .A2(\hash/CA2/_0284_ ),
    .B1(\hash/CA2/_1145_ ),
    .Y(\hash/CA2/_0285_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1850_  (.A(\hash/CA2/_1150_ ),
    .B(\hash/CA2/_0285_ ),
    .Y(\hash/a_new[15] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1851_  (.A1(\hash/CA2/_1146_ ),
    .A2(\hash/CA2/_0276_ ),
    .B1(\hash/CA2/_1145_ ),
    .X(\hash/CA2/_0286_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1852_  (.A1(\hash/CA2/_1150_ ),
    .A2(\hash/CA2/_0286_ ),
    .B1(\hash/CA2/_1149_ ),
    .Y(\hash/CA2/_0287_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1853_  (.A(\hash/CA2/_1154_ ),
    .B(\hash/CA2/_0287_ ),
    .Y(\hash/a_new[16] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1854_  (.A1(\hash/CA2/_1146_ ),
    .A2(\hash/CA2/_1145_ ),
    .B1(\hash/CA2/_1150_ ),
    .Y(\hash/CA2/_0288_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1855_  (.A_N(\hash/CA2/_1149_ ),
    .B(\hash/CA2/_0288_ ),
    .Y(\hash/CA2/_0289_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1856_  (.A1(\hash/CA2/_1154_ ),
    .A2(\hash/CA2/_0289_ ),
    .B1(\hash/CA2/_1153_ ),
    .Y(\hash/CA2/_0290_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1857_  (.A1(\hash/CA2/_1154_ ),
    .A2(\hash/CA2/_1149_ ),
    .B1(\hash/CA2/_1153_ ),
    .C1(\hash/CA2/_1145_ ),
    .Y(\hash/CA2/_0291_ ));
 sky130_fd_sc_hd__o311ai_0 \hash/CA2/_1858_  (.A1(\hash/CA2/_0267_ ),
    .A2(\hash/CA2/_0277_ ),
    .A3(\hash/CA2/_0278_ ),
    .B1(\hash/CA2/_0283_ ),
    .C1(\hash/CA2/_0291_ ),
    .Y(\hash/CA2/_0292_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1859_  (.A1(\hash/CA2/_0257_ ),
    .A2(\hash/CA2/_0280_ ),
    .B1(\hash/CA2/_0292_ ),
    .Y(\hash/CA2/_0293_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1860_  (.A(\hash/CA2/_0290_ ),
    .B(\hash/CA2/_0293_ ),
    .Y(\hash/CA2/_0294_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1861_  (.A(\hash/CA2/_1158_ ),
    .B(\hash/CA2/_0294_ ),
    .X(\hash/a_new[17] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1862_  (.A(\hash/CA2/_1162_ ),
    .Y(\hash/CA2/_0295_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1863_  (.A1(\hash/CA2/_1150_ ),
    .A2(\hash/CA2/_1145_ ),
    .B1(\hash/CA2/_1149_ ),
    .X(\hash/CA2/_0296_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1864_  (.A1(\hash/CA2/_1154_ ),
    .A2(\hash/CA2/_0296_ ),
    .B1(\hash/CA2/_1153_ ),
    .X(\hash/CA2/_0297_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1865_  (.A1(\hash/CA2/_1158_ ),
    .A2(\hash/CA2/_0297_ ),
    .B1(\hash/CA2/_1157_ ),
    .Y(\hash/CA2/_0298_ ));
 sky130_fd_sc_hd__and4_1 \hash/CA2/_1866_  (.A(\hash/CA2/_1146_ ),
    .B(\hash/CA2/_1150_ ),
    .C(\hash/CA2/_1154_ ),
    .D(\hash/CA2/_1158_ ),
    .X(\hash/CA2/_0299_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1867_  (.A(\hash/CA2/_0276_ ),
    .B(\hash/CA2/_0299_ ),
    .Y(\hash/CA2/_0300_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1868_  (.A(\hash/CA2/_0298_ ),
    .B(\hash/CA2/_0300_ ),
    .Y(\hash/CA2/_0301_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1869_  (.A(\hash/CA2/_0295_ ),
    .B(\hash/CA2/_0301_ ),
    .Y(\hash/a_new[18] ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1870_  (.A1(\hash/CA2/_1158_ ),
    .A2(\hash/CA2/_0294_ ),
    .B1(\hash/CA2/_1157_ ),
    .Y(\hash/CA2/_0302_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1871_  (.A1(\hash/CA2/_0295_ ),
    .A2(\hash/CA2/_0302_ ),
    .B1_N(\hash/CA2/_1161_ ),
    .Y(\hash/CA2/_0303_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1872_  (.A(\hash/CA2/_1166_ ),
    .B(\hash/CA2/_0303_ ),
    .X(\hash/a_new[19] ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1873_  (.A(\hash/CA2/_1162_ ),
    .B(\hash/CA2/_1166_ ),
    .C(\hash/CA2/_0299_ ),
    .Y(\hash/CA2/_0304_ ));
 sky130_fd_sc_hd__or3_1 \hash/CA2/_1874_  (.A(\hash/CA2/_0272_ ),
    .B(\hash/CA2/_0275_ ),
    .C(\hash/CA2/_0304_ ),
    .X(\hash/CA2/_0305_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1875_  (.A1(\hash/CA2/_0295_ ),
    .A2(\hash/CA2/_0298_ ),
    .B1_N(\hash/CA2/_1161_ ),
    .Y(\hash/CA2/_0306_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1876_  (.A1(\hash/CA2/_1166_ ),
    .A2(\hash/CA2/_0306_ ),
    .B1(\hash/CA2/_1165_ ),
    .Y(\hash/CA2/_0307_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1877_  (.A(\hash/CA2/_0305_ ),
    .B(\hash/CA2/_0307_ ),
    .Y(\hash/CA2/_0308_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1878_  (.A(\hash/CA2/_1170_ ),
    .B(\hash/CA2/_0308_ ),
    .X(\hash/a_new[20] ));
 sky130_fd_sc_hd__nand4_1 \hash/CA2/_1879_  (.A(\hash/CA2/_1158_ ),
    .B(\hash/CA2/_1162_ ),
    .C(\hash/CA2/_1166_ ),
    .D(\hash/CA2/_1170_ ),
    .Y(\hash/CA2/_0309_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_1880_  (.A(\hash/CA2/_1162_ ),
    .B(\hash/CA2/_1157_ ),
    .X(\hash/CA2/_0310_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA2/_1881_  (.A1(\hash/CA2/_1161_ ),
    .A2(\hash/CA2/_0310_ ),
    .B1(\hash/CA2/_1166_ ),
    .C1(\hash/CA2/_1170_ ),
    .Y(\hash/CA2/_0311_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1882_  (.A1(\hash/CA2/_0290_ ),
    .A2(\hash/CA2/_0309_ ),
    .B1(\hash/CA2/_0311_ ),
    .Y(\hash/CA2/_0312_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1883_  (.A(\hash/CA2/_1161_ ),
    .B(\hash/CA2/_0310_ ),
    .Y(\hash/CA2/_0313_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1884_  (.A(\hash/CA2/_0293_ ),
    .B(\hash/CA2/_0313_ ),
    .Y(\hash/CA2/_0314_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1885_  (.A1(\hash/CA2/_1170_ ),
    .A2(\hash/CA2/_1165_ ),
    .B1(\hash/CA2/_1169_ ),
    .X(\hash/CA2/_0315_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1886_  (.A1(\hash/CA2/_0312_ ),
    .A2(\hash/CA2/_0314_ ),
    .B1(\hash/CA2/_0315_ ),
    .Y(\hash/CA2/_0316_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1887_  (.A(\hash/CA2/_1174_ ),
    .B(\hash/CA2/_0316_ ),
    .Y(\hash/a_new[21] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1888_  (.A1(\hash/CA2/_1170_ ),
    .A2(\hash/CA2/_0308_ ),
    .B1(\hash/CA2/_1169_ ),
    .X(\hash/CA2/_0317_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1889_  (.A(\hash/CA2/_1174_ ),
    .B(\hash/CA2/_0317_ ),
    .Y(\hash/CA2/_0318_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1890_  (.A(\hash/CA2/_1178_ ),
    .B(\hash/CA2/_1173_ ),
    .Y(\hash/CA2/_0319_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1891_  (.A(\hash/CA2/_1178_ ),
    .B(\hash/CA2/_1173_ ),
    .Y(\hash/CA2/_0320_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1892_  (.A(\hash/CA2/_1174_ ),
    .B(\hash/CA2/_1178_ ),
    .C(\hash/CA2/_1169_ ),
    .Y(\hash/CA2/_0321_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1893_  (.A(\hash/CA2/_0320_ ),
    .B(\hash/CA2/_0321_ ),
    .Y(\hash/CA2/_0322_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1894_  (.A(\hash/CA2/_1170_ ),
    .B(\hash/CA2/_1174_ ),
    .C(\hash/CA2/_1178_ ),
    .Y(\hash/CA2/_0323_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1895_  (.A1(\hash/CA2/_0305_ ),
    .A2(\hash/CA2/_0307_ ),
    .B1(\hash/CA2/_0323_ ),
    .Y(\hash/CA2/_0324_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_1896_  (.A1(\hash/CA2/_0318_ ),
    .A2(\hash/CA2/_0319_ ),
    .B1(\hash/CA2/_0322_ ),
    .C1(\hash/CA2/_0324_ ),
    .Y(\hash/a_new[22] ));
 sky130_fd_sc_hd__nor4_1 \hash/CA2/_1897_  (.A(\hash/CA2/_1161_ ),
    .B(\hash/CA2/_0292_ ),
    .C(\hash/CA2/_0315_ ),
    .D(\hash/CA2/_0310_ ),
    .Y(\hash/CA2/_0325_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA2/_1898_  (.A1(\hash/CA2/_0257_ ),
    .A2(\hash/CA2/_0280_ ),
    .B1_N(\hash/CA2/_0325_ ),
    .Y(\hash/CA2/_0326_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1899_  (.A1(\hash/CA2/_0315_ ),
    .A2(\hash/CA2/_0312_ ),
    .B1(\hash/CA2/_1174_ ),
    .Y(\hash/CA2/_0327_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1900_  (.A1(\hash/CA2/_0326_ ),
    .A2(\hash/CA2/_0327_ ),
    .B1_N(\hash/CA2/_1173_ ),
    .Y(\hash/CA2/_0328_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1901_  (.A1(\hash/CA2/_1178_ ),
    .A2(\hash/CA2/_0328_ ),
    .B1(\hash/CA2/_1177_ ),
    .Y(\hash/CA2/_0329_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1902_  (.A(\hash/CA2/_1182_ ),
    .B(\hash/CA2/_0329_ ),
    .Y(\hash/a_new[23] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1903_  (.A(\hash/CA2/_1182_ ),
    .Y(\hash/CA2/_0330_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1904_  (.A(\hash/CA2/_1177_ ),
    .B(\hash/CA2/_0324_ ),
    .C(\hash/CA2/_0322_ ),
    .Y(\hash/CA2/_0331_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1905_  (.A1(\hash/CA2/_0330_ ),
    .A2(\hash/CA2/_0331_ ),
    .B1_N(\hash/CA2/_1181_ ),
    .Y(\hash/CA2/_0332_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1906_  (.A(\hash/CA2/_1186_ ),
    .B(\hash/CA2/_0332_ ),
    .X(\hash/a_new[24] ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1907_  (.A1(\hash/CA2/_0330_ ),
    .A2(\hash/CA2/_0329_ ),
    .B1_N(\hash/CA2/_1181_ ),
    .Y(\hash/CA2/_0333_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1908_  (.A1(\hash/CA2/_1186_ ),
    .A2(\hash/CA2/_0333_ ),
    .B1(\hash/CA2/_1185_ ),
    .Y(\hash/CA2/_0334_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1909_  (.A(\hash/CA2/_1190_ ),
    .B(\hash/CA2/_0334_ ),
    .Y(\hash/a_new[25] ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1910_  (.A(\hash/CA2/_1182_ ),
    .B(\hash/CA2/_1186_ ),
    .C(\hash/CA2/_1190_ ),
    .Y(\hash/CA2/_0335_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1911_  (.A1(\hash/CA2/_1186_ ),
    .A2(\hash/CA2/_1181_ ),
    .B1(\hash/CA2/_1185_ ),
    .X(\hash/CA2/_0336_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1912_  (.A1(\hash/CA2/_1190_ ),
    .A2(\hash/CA2/_0336_ ),
    .B1(\hash/CA2/_1189_ ),
    .Y(\hash/CA2/_0337_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1913_  (.A1(\hash/CA2/_0331_ ),
    .A2(\hash/CA2/_0335_ ),
    .B1(\hash/CA2/_0337_ ),
    .Y(\hash/CA2/_0338_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1914_  (.A(\hash/CA2/_1194_ ),
    .B(\hash/CA2/_0338_ ),
    .X(\hash/a_new[26] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1915_  (.A(\hash/CA2/_1173_ ),
    .B(\hash/CA2/_1177_ ),
    .Y(\hash/CA2/_0339_ ));
 sky130_fd_sc_hd__o211a_1 \hash/CA2/_1916_  (.A1(\hash/CA2/_0326_ ),
    .A2(\hash/CA2/_0327_ ),
    .B1(\hash/CA2/_0337_ ),
    .C1(\hash/CA2/_0339_ ),
    .X(\hash/CA2/_0340_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1917_  (.A(\hash/CA2/_1178_ ),
    .B(\hash/CA2/_1177_ ),
    .Y(\hash/CA2/_0341_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1918_  (.A1(\hash/CA2/_0335_ ),
    .A2(\hash/CA2/_0341_ ),
    .B1(\hash/CA2/_0337_ ),
    .X(\hash/CA2/_0342_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1919_  (.A(\hash/CA2/_0340_ ),
    .B(\hash/CA2/_0342_ ),
    .Y(\hash/CA2/_0343_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1920_  (.A1(\hash/CA2/_1194_ ),
    .A2(\hash/CA2/_0343_ ),
    .B1(\hash/CA2/_1193_ ),
    .Y(\hash/CA2/_0344_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1921_  (.A(\hash/CA2/_1198_ ),
    .B(\hash/CA2/_0344_ ),
    .Y(\hash/a_new[27] ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_1922_  (.A(\hash/CA2/_1202_ ),
    .B_N(\hash/CA2/_1198_ ),
    .Y(\hash/CA2/_0345_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1923_  (.A(\hash/CA2/_1202_ ),
    .Y(\hash/CA2/_0346_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1924_  (.A(\hash/CA2/_0346_ ),
    .B(\hash/CA2/_1193_ ),
    .C(\hash/CA2/_1197_ ),
    .Y(\hash/CA2/_0347_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1925_  (.A_N(\hash/CA2/_1177_ ),
    .B(\hash/CA2/_0337_ ),
    .Y(\hash/CA2/_0348_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA2/_1926_  (.A1(\hash/CA2/_0337_ ),
    .A2(\hash/CA2/_0335_ ),
    .B1_N(\hash/CA2/_1194_ ),
    .Y(\hash/CA2/_0349_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_1927_  (.A1(\hash/CA2/_0324_ ),
    .A2(\hash/CA2/_0322_ ),
    .A3(\hash/CA2/_0348_ ),
    .B1(\hash/CA2/_0349_ ),
    .Y(\hash/CA2/_0350_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA2/_1928_  (.A0(\hash/CA2/_0345_ ),
    .A1(\hash/CA2/_0347_ ),
    .S(\hash/CA2/_0350_ ),
    .Y(\hash/CA2/_0351_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1929_  (.A(\hash/CA2/_1198_ ),
    .B(\hash/CA2/_0346_ ),
    .C(\hash/CA2/_1197_ ),
    .Y(\hash/CA2/_0352_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA2/_1930_  (.A1(\hash/CA2/_0346_ ),
    .A2(\hash/CA2/_1197_ ),
    .B1(\hash/CA2/_0345_ ),
    .B2(\hash/CA2/_1193_ ),
    .C1(\hash/CA2/_0352_ ),
    .Y(\hash/CA2/_0353_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1931_  (.A(\hash/CA2/_0351_ ),
    .B(\hash/CA2/_0353_ ),
    .Y(\hash/a_new[28] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1932_  (.A(\hash/CA2/_1198_ ),
    .B(\hash/CA2/_1202_ ),
    .Y(\hash/CA2/_0354_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1933_  (.A1(\hash/CA2/_1202_ ),
    .A2(\hash/CA2/_1197_ ),
    .B1(\hash/CA2/_1201_ ),
    .Y(\hash/CA2/_0355_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1934_  (.A1(\hash/CA2/_0344_ ),
    .A2(\hash/CA2/_0354_ ),
    .B1(\hash/CA2/_0355_ ),
    .Y(\hash/CA2/_0356_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1935_  (.A(\hash/CA2/_1206_ ),
    .B(\hash/CA2/_0356_ ),
    .X(\hash/a_new[29] ));
 sky130_fd_sc_hd__nand4_1 \hash/CA2/_1936_  (.A(\hash/CA2/_1194_ ),
    .B(\hash/CA2/_1198_ ),
    .C(\hash/CA2/_1202_ ),
    .D(\hash/CA2/_1206_ ),
    .Y(\hash/CA2/_0357_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1937_  (.A1(\hash/CA2/_1198_ ),
    .A2(\hash/CA2/_1193_ ),
    .B1(\hash/CA2/_1197_ ),
    .Y(\hash/CA2/_0358_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1938_  (.A1(\hash/CA2/_0346_ ),
    .A2(\hash/CA2/_0358_ ),
    .B1_N(\hash/CA2/_1201_ ),
    .Y(\hash/CA2/_0359_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1939_  (.A1(\hash/CA2/_1206_ ),
    .A2(\hash/CA2/_0359_ ),
    .B1(\hash/CA2/_1205_ ),
    .Y(\hash/CA2/_0360_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1940_  (.A1(\hash/CA2/_0337_ ),
    .A2(\hash/CA2/_0357_ ),
    .B1(\hash/CA2/_0360_ ),
    .X(\hash/CA2/_0361_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_1941_  (.A1(\hash/CA2/_0331_ ),
    .A2(\hash/CA2/_0335_ ),
    .A3(\hash/CA2/_0357_ ),
    .B1(\hash/CA2/_0361_ ),
    .Y(\hash/CA2/_0362_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1942_  (.A(\hash/CA2/_1209_ ),
    .B(\hash/CA2/_0362_ ),
    .X(\hash/a_new[30] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1943_  (.A(\hash/CA2/_1092_ ),
    .B(\hash/CA2/_1097_ ),
    .Y(\hash/CA2/_0363_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_1944_  (.A(\hash/CA2/_1093_ ),
    .B(\hash/CA2/_1092_ ),
    .C(\hash/CA2/_1097_ ),
    .Y(\hash/CA2/_0364_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1945_  (.A(\hash/CA2/_1098_ ),
    .B(\hash/CA2/_1097_ ),
    .Y(\hash/CA2/_0365_ ));
 sky130_fd_sc_hd__a311oi_2 \hash/CA2/_1946_  (.A1(\hash/CA2/_0035_ ),
    .A2(\hash/CA2/_0041_ ),
    .A3(\hash/CA2/_0363_ ),
    .B1(\hash/CA2/_0364_ ),
    .C1(\hash/CA2/_0365_ ),
    .Y(\hash/CA2/_0366_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/CA2/_1947_  (.A0(\hash/f_cap[31] ),
    .A1(\hash/e_cap[31] ),
    .S(\hash/p2_cap[31] ),
    .Y(\hash/CA2/_0367_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1948_  (.A(\hash/CA2/s1[31] ),
    .B(\hash/CA2/_0367_ ),
    .X(\hash/CA2/_0368_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1949_  (.A(\hash/CA2/_0366_ ),
    .B(\hash/CA2/_0368_ ),
    .Y(\hash/CA2/_0369_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1950_  (.A(\hash/CA2/_0860_ ),
    .B(\hash/CA2/_0864_ ),
    .X(\hash/CA2/_0370_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1951_  (.A(\hash/p4_cap[31] ),
    .B(\hash/CA2/s0[31] ),
    .Y(\hash/CA2/_0371_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1952_  (.A(\hash/CA2/_0370_ ),
    .B(\hash/CA2/_0371_ ),
    .Y(\hash/CA2/_0372_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_1953_  (.A1(\hash/CA2/_0340_ ),
    .A2(\hash/CA2/_0342_ ),
    .A3(\hash/CA2/_0357_ ),
    .B1(\hash/CA2/_0360_ ),
    .Y(\hash/CA2/_0373_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1954_  (.A1(\hash/CA2/_1209_ ),
    .A2(\hash/CA2/_0373_ ),
    .B1(\hash/CA2/_1208_ ),
    .Y(\hash/CA2/_0374_ ));
 sky130_fd_sc_hd__xnor3_1 \hash/CA2/_1955_  (.A(\hash/CA2/_0369_ ),
    .B(\hash/CA2/_0372_ ),
    .C(\hash/CA2/_0374_ ),
    .X(\hash/CA2/_0375_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1956_  (.A(\hash/p1_cap[31] ),
    .B(\hash/p3_cap[31] ),
    .Y(\hash/CA2/_0376_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1957_  (.A(\hash/CA2/_0931_ ),
    .Y(\hash/CA2/_0377_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_1958_  (.A(\hash/CA2/_0925_ ),
    .B(\hash/CA2/_0927_ ),
    .C(\hash/CA2/_0929_ ),
    .X(\hash/CA2/_0378_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_1959_  (.A(\hash/CA2/_0925_ ),
    .B(\hash/CA2/_0927_ ),
    .C(\hash/CA2/_0929_ ),
    .Y(\hash/CA2/_0379_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/CA2/_1960_  (.A1(\hash/CA2/_0235_ ),
    .A2(\hash/CA2/_0233_ ),
    .B1(\hash/CA2/_0379_ ),
    .B2(\hash/CA2/_0198_ ),
    .Y(\hash/CA2/_0380_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/CA2/_1961_  (.A1(\hash/CA2/_0170_ ),
    .A2(\hash/CA2/_0195_ ),
    .A3(\hash/CA2/_0378_ ),
    .B1(\hash/CA2/_0380_ ),
    .C1(\hash/CA2/_0928_ ),
    .Y(\hash/CA2/_0381_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1962_  (.A1(\hash/CA2/_0377_ ),
    .A2(\hash/CA2/_0381_ ),
    .B1_N(\hash/CA2/_0930_ ),
    .Y(\hash/CA2/_0382_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1963_  (.A(\hash/CA2/_0376_ ),
    .B(\hash/CA2/_0382_ ),
    .Y(\hash/b_new[31] ));
 sky130_fd_sc_hd__maj3_1 \hash/CA2/_1964_  (.A(\hash/b_cap[31] ),
    .B(\hash/a_cap[31] ),
    .C(\hash/b_new[31] ),
    .X(\hash/CA2/_0383_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1965_  (.A(\hash/CA2/_0375_ ),
    .B(\hash/CA2/_0383_ ),
    .X(\hash/a_new[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1966_  (.A(\hash/CA2/_0867_ ),
    .B(\hash/CA2/_1108_ ),
    .Y(\hash/a_new[3] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1967_  (.A(\hash/CA2/_1112_ ),
    .B(\hash/CA2/_0241_ ),
    .Y(\hash/a_new[4] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1968_  (.A(\hash/CA2/_1111_ ),
    .B(\hash/CA2/_0251_ ),
    .Y(\hash/CA2/_0384_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1969_  (.A(\hash/CA2/_1115_ ),
    .B(\hash/CA2/_0384_ ),
    .Y(\hash/a_new[5] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1970_  (.A(\hash/CA2/_1117_ ),
    .B(\hash/CA2/_1114_ ),
    .Y(\hash/CA2/_0385_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1971_  (.A(\hash/CA2/_0239_ ),
    .B(\hash/CA2/_0241_ ),
    .Y(\hash/CA2/_0386_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1972_  (.A1(\hash/CA2/_1111_ ),
    .A2(\hash/CA2/_0386_ ),
    .B1(\hash/CA2/_1115_ ),
    .Y(\hash/CA2/_0387_ ));
 sky130_fd_sc_hd__a22oi_1 \hash/CA2/_1973_  (.A1(\hash/CA2/_0243_ ),
    .A2(\hash/CA2/_0244_ ),
    .B1(\hash/CA2/_0385_ ),
    .B2(\hash/CA2/_0387_ ),
    .Y(\hash/a_new[6] ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_1974_  (.A_N(\hash/CA2/_1114_ ),
    .B(\hash/CA2/_0252_ ),
    .Y(\hash/CA2/_0388_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1975_  (.A1(\hash/CA2/_1117_ ),
    .A2(\hash/CA2/_0388_ ),
    .B1(\hash/CA2/_1116_ ),
    .Y(\hash/CA2/_0389_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1976_  (.A(\hash/CA2/_1119_ ),
    .B(\hash/CA2/_0389_ ),
    .Y(\hash/a_new[7] ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1977_  (.A(\hash/CA2/_1118_ ),
    .B(\hash/CA2/_0246_ ),
    .Y(\hash/CA2/_0390_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1978_  (.A(\hash/CA2/_1122_ ),
    .B(\hash/CA2/_0390_ ),
    .Y(\hash/a_new[8] ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_1979_  (.A(\hash/CA2/_1126_ ),
    .B(\hash/CA2/_0257_ ),
    .X(\hash/a_new[9] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1980_  (.A(\hash/CA2/_0108_ ),
    .Y(\hash/b_new[15] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1981_  (.A(\hash/CA2/_0138_ ),
    .Y(\hash/b_new[19] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1982_  (.A(\hash/CA2/_0143_ ),
    .Y(\hash/b_new[20] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1983_  (.A1(\hash/CA2/_0207_ ),
    .A2(\hash/CA2/_0203_ ),
    .B1(\hash/CA2/_0205_ ),
    .Y(\hash/CA2/_0391_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1984_  (.A(\hash/CA2/_0209_ ),
    .B(\hash/CA2/_0391_ ),
    .Y(\hash/b_new[28] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_1985_  (.A1(\hash/CA2/_0967_ ),
    .A2(\hash/CA2/_0966_ ),
    .B1(\hash/CA2/_0972_ ),
    .Y(\hash/CA2/_0392_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1986_  (.A(\hash/CA2/_0971_ ),
    .B(\hash/CA2/_0977_ ),
    .Y(\hash/CA2/_0393_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1987_  (.A(\hash/CA2/_0978_ ),
    .B(\hash/CA2/_0977_ ),
    .Y(\hash/CA2/_0394_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1988_  (.A1(\hash/CA2/_0392_ ),
    .A2(\hash/CA2/_0393_ ),
    .B1(\hash/CA2/_0394_ ),
    .Y(\hash/CA2/_0395_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1989_  (.A(\hash/CA2/_0962_ ),
    .Y(\hash/CA2/_0396_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_1990_  (.A(\hash/CA2/_0952_ ),
    .Y(\hash/CA2/_0397_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_1991_  (.A1(\hash/CA2/_0870_ ),
    .A2(\hash/CA2/_0942_ ),
    .B1(\hash/CA2/_0941_ ),
    .X(\hash/CA2/_0398_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1992_  (.A1(\hash/CA2/_0947_ ),
    .A2(\hash/CA2/_0398_ ),
    .B1(\hash/CA2/_0946_ ),
    .Y(\hash/CA2/_0399_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_1993_  (.A1(\hash/CA2/_0397_ ),
    .A2(\hash/CA2/_0399_ ),
    .B1_N(\hash/CA2/_0951_ ),
    .Y(\hash/CA2/_0400_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_1994_  (.A1(\hash/CA2/_0957_ ),
    .A2(\hash/CA2/_0400_ ),
    .B1(\hash/CA2/_0956_ ),
    .Y(\hash/CA2/_0401_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_1995_  (.A(\hash/CA2/_0961_ ),
    .B(\hash/CA2/_0966_ ),
    .Y(\hash/CA2/_0402_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA2/_1996_  (.A1(\hash/CA2/_0396_ ),
    .A2(\hash/CA2/_0401_ ),
    .B1(\hash/CA2/_0402_ ),
    .C1(\hash/CA2/_0393_ ),
    .Y(\hash/CA2/_0403_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_1997_  (.A(\hash/CA2/_0395_ ),
    .B(\hash/CA2/_0403_ ),
    .Y(\hash/CA2/_0404_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_1998_  (.A(\hash/CA2/_0984_ ),
    .B(\hash/CA2/_0404_ ),
    .Y(\hash/e_new[10] ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_1999_  (.A1(\hash/CA2/_0952_ ),
    .A2(\hash/CA2/_0951_ ),
    .B1(\hash/CA2/_0957_ ),
    .X(\hash/CA2/_0405_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2000_  (.A1(\hash/CA2/_0956_ ),
    .A2(\hash/CA2/_0405_ ),
    .B1(\hash/CA2/_0962_ ),
    .Y(\hash/CA2/_0406_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2001_  (.A1(\hash/CA2/_0869_ ),
    .A2(\hash/CA2/_0937_ ),
    .B1(\hash/CA2/_0936_ ),
    .X(\hash/CA2/_0407_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2002_  (.A1(\hash/CA2/_0947_ ),
    .A2(\hash/CA2/_0941_ ),
    .B1(\hash/CA2/_0946_ ),
    .X(\hash/CA2/_0408_ ));
 sky130_fd_sc_hd__or4_1 \hash/CA2/_2003_  (.A(\hash/CA2/_0951_ ),
    .B(\hash/CA2/_0956_ ),
    .C(\hash/CA2/_0961_ ),
    .D(\hash/CA2/_0966_ ),
    .X(\hash/CA2/_0409_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/CA2/_2004_  (.A1(\hash/CA2/_0942_ ),
    .A2(\hash/CA2/_0947_ ),
    .A3(\hash/CA2/_0407_ ),
    .B1(\hash/CA2/_0408_ ),
    .C1(\hash/CA2/_0409_ ),
    .Y(\hash/CA2/_0410_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/CA2/_2005_  (.A1(\hash/CA2/_0402_ ),
    .A2(\hash/CA2/_0406_ ),
    .B1(\hash/CA2/_0410_ ),
    .C1(\hash/CA2/_0392_ ),
    .Y(\hash/CA2/_0411_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_2006_  (.A1(\hash/CA2/_0971_ ),
    .A2(\hash/CA2/_0411_ ),
    .B1(\hash/CA2/_0978_ ),
    .X(\hash/CA2/_0412_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2007_  (.A1(\hash/CA2/_0977_ ),
    .A2(\hash/CA2/_0412_ ),
    .B1(\hash/CA2/_0984_ ),
    .Y(\hash/CA2/_0413_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_2008_  (.A(\hash/CA2/_0983_ ),
    .B_N(\hash/CA2/_0413_ ),
    .Y(\hash/CA2/_0414_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2009_  (.A(\hash/CA2/_0990_ ),
    .B(\hash/CA2/_0414_ ),
    .Y(\hash/e_new[11] ));
 sky130_fd_sc_hd__a31o_2 \hash/CA2/_2010_  (.A1(\hash/CA2/_0984_ ),
    .A2(\hash/CA2/_0395_ ),
    .A3(\hash/CA2/_0403_ ),
    .B1(\hash/CA2/_0983_ ),
    .X(\hash/CA2/_0415_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2011_  (.A1(\hash/CA2/_0990_ ),
    .A2(\hash/CA2/_0415_ ),
    .B1(\hash/CA2/_0989_ ),
    .Y(\hash/CA2/_0416_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2012_  (.A(\hash/CA2/_0996_ ),
    .B(\hash/CA2/_0416_ ),
    .Y(\hash/e_new[12] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_2013_  (.A(\hash/CA2/_0990_ ),
    .Y(\hash/CA2/_0417_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_2014_  (.A1(\hash/CA2/_0417_ ),
    .A2(\hash/CA2/_0414_ ),
    .B1_N(\hash/CA2/_0989_ ),
    .Y(\hash/CA2/_0418_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2015_  (.A1(\hash/CA2/_0996_ ),
    .A2(\hash/CA2/_0418_ ),
    .B1(\hash/CA2/_0995_ ),
    .Y(\hash/CA2/_0419_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2016_  (.A(\hash/CA2/_1002_ ),
    .B(\hash/CA2/_0419_ ),
    .Y(\hash/e_new[13] ));
 sky130_fd_sc_hd__and4_1 \hash/CA2/_2017_  (.A(\hash/CA2/_0984_ ),
    .B(\hash/CA2/_0990_ ),
    .C(\hash/CA2/_0996_ ),
    .D(\hash/CA2/_1002_ ),
    .X(\hash/CA2/_0420_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_2018_  (.A(\hash/CA2/_0996_ ),
    .Y(\hash/CA2/_0421_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2019_  (.A1(\hash/CA2/_0990_ ),
    .A2(\hash/CA2/_0983_ ),
    .B1(\hash/CA2/_0989_ ),
    .Y(\hash/CA2/_0422_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/CA2/_2020_  (.A1(\hash/CA2/_0421_ ),
    .A2(\hash/CA2/_0422_ ),
    .B1_N(\hash/CA2/_0995_ ),
    .Y(\hash/CA2/_0423_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2021_  (.A1(\hash/CA2/_1002_ ),
    .A2(\hash/CA2/_0423_ ),
    .B1(\hash/CA2/_1001_ ),
    .Y(\hash/CA2/_0424_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_2022_  (.A(\hash/CA2/_0424_ ),
    .Y(\hash/CA2/_0425_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA2/_2023_  (.A1(\hash/CA2/_0395_ ),
    .A2(\hash/CA2/_0403_ ),
    .A3(\hash/CA2/_0420_ ),
    .B1(\hash/CA2/_0425_ ),
    .Y(\hash/CA2/_0426_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2024_  (.A(\hash/CA2/_1008_ ),
    .B(\hash/CA2/_0426_ ),
    .Y(\hash/e_new[14] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2025_  (.A1(\hash/CA2/_0984_ ),
    .A2(\hash/CA2/_0977_ ),
    .B1(\hash/CA2/_0983_ ),
    .X(\hash/CA2/_0427_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2026_  (.A1(\hash/CA2/_0990_ ),
    .A2(\hash/CA2/_0427_ ),
    .B1(\hash/CA2/_0989_ ),
    .Y(\hash/CA2/_0428_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_2027_  (.A(\hash/CA2/_0995_ ),
    .B(\hash/CA2/_1001_ ),
    .C(\hash/CA2/_1007_ ),
    .Y(\hash/CA2/_0429_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2028_  (.A1(\hash/CA2/_0421_ ),
    .A2(\hash/CA2/_0428_ ),
    .B1(\hash/CA2/_0429_ ),
    .Y(\hash/CA2/_0430_ ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_2029_  (.A(\hash/CA2/_1002_ ),
    .B(\hash/CA2/_1001_ ),
    .C(\hash/CA2/_1007_ ),
    .Y(\hash/CA2/_0431_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_2030_  (.A(\hash/CA2/_1008_ ),
    .B(\hash/CA2/_1007_ ),
    .Y(\hash/CA2/_0432_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_2031_  (.A(\hash/CA2/_0431_ ),
    .B(\hash/CA2/_0432_ ),
    .Y(\hash/CA2/_0433_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_2032_  (.A(\hash/CA2/_1008_ ),
    .B(\hash/CA2/_0420_ ),
    .X(\hash/CA2/_0434_ ));
 sky130_fd_sc_hd__a22o_1 \hash/CA2/_2033_  (.A1(\hash/CA2/_0430_ ),
    .A2(\hash/CA2/_0433_ ),
    .B1(\hash/CA2/_0434_ ),
    .B2(\hash/CA2/_0412_ ),
    .X(\hash/CA2/_0435_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_2034_  (.A(\hash/CA2/_1014_ ),
    .B(\hash/CA2/_0435_ ),
    .X(\hash/e_new[15] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2035_  (.A(\hash/CA2/_1008_ ),
    .B(\hash/CA2/_1014_ ),
    .Y(\hash/CA2/_0436_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2036_  (.A1(\hash/CA2/_1014_ ),
    .A2(\hash/CA2/_1007_ ),
    .B1(\hash/CA2/_1013_ ),
    .Y(\hash/CA2/_0437_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2037_  (.A1(\hash/CA2/_0426_ ),
    .A2(\hash/CA2/_0436_ ),
    .B1(\hash/CA2/_0437_ ),
    .Y(\hash/CA2/_0438_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_2038_  (.A(\hash/CA2/_1019_ ),
    .B(\hash/CA2/_0438_ ),
    .X(\hash/e_new[16] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2039_  (.A1(\hash/CA2/_1014_ ),
    .A2(\hash/CA2/_0435_ ),
    .B1(\hash/CA2/_1013_ ),
    .X(\hash/CA2/_0439_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2040_  (.A1(\hash/CA2/_1019_ ),
    .A2(\hash/CA2/_0439_ ),
    .B1(\hash/CA2/_1018_ ),
    .Y(\hash/CA2/_0440_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2041_  (.A(\hash/CA2/_1025_ ),
    .B(\hash/CA2/_0440_ ),
    .Y(\hash/e_new[17] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2042_  (.A1(\hash/CA2/_1019_ ),
    .A2(\hash/CA2/_0438_ ),
    .B1(\hash/CA2/_1018_ ),
    .X(\hash/CA2/_0441_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2043_  (.A1(\hash/CA2/_1025_ ),
    .A2(\hash/CA2/_0441_ ),
    .B1(\hash/CA2/_1024_ ),
    .Y(\hash/CA2/_0442_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2044_  (.A(\hash/CA2/_1031_ ),
    .B(\hash/CA2/_0442_ ),
    .Y(\hash/e_new[18] ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_2045_  (.A(\hash/CA2/_1014_ ),
    .B(\hash/CA2/_1019_ ),
    .C(\hash/CA2/_1025_ ),
    .X(\hash/CA2/_0443_ ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_2046_  (.A(\hash/CA2/_1008_ ),
    .B(\hash/CA2/_0420_ ),
    .C(\hash/CA2/_0443_ ),
    .X(\hash/CA2/_0444_ ));
 sky130_fd_sc_hd__o211ai_2 \hash/CA2/_2047_  (.A1(\hash/CA2/_0971_ ),
    .A2(\hash/CA2/_0411_ ),
    .B1(\hash/CA2/_0444_ ),
    .C1(\hash/CA2/_0978_ ),
    .Y(\hash/CA2/_0445_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2048_  (.A1(\hash/CA2/_1019_ ),
    .A2(\hash/CA2/_1013_ ),
    .B1(\hash/CA2/_1018_ ),
    .X(\hash/CA2/_0446_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2049_  (.A1(\hash/CA2/_1025_ ),
    .A2(\hash/CA2/_0446_ ),
    .B1(\hash/CA2/_1024_ ),
    .X(\hash/CA2/_0447_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/CA2/_2050_  (.A1(\hash/CA2/_0430_ ),
    .A2(\hash/CA2/_0433_ ),
    .A3(\hash/CA2/_0443_ ),
    .B1(\hash/CA2/_0447_ ),
    .Y(\hash/CA2/_0448_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2051_  (.A(\hash/CA2/_0445_ ),
    .B(\hash/CA2/_0448_ ),
    .Y(\hash/CA2/_0449_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2052_  (.A1(\hash/CA2/_1031_ ),
    .A2(\hash/CA2/_0449_ ),
    .B1(\hash/CA2/_1030_ ),
    .Y(\hash/CA2/_0450_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2053_  (.A(\hash/CA2/_1037_ ),
    .B(\hash/CA2/_0450_ ),
    .Y(\hash/e_new[19] ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2054_  (.A1(\hash/CA2/_1031_ ),
    .A2(\hash/CA2/_0447_ ),
    .B1(\hash/CA2/_1030_ ),
    .Y(\hash/CA2/_0451_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2055_  (.A(\hash/CA2/_0424_ ),
    .B(\hash/CA2/_0451_ ),
    .Y(\hash/CA2/_0452_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/CA2/_2056_  (.A1(\hash/CA2/_0395_ ),
    .A2(\hash/CA2/_0403_ ),
    .A3(\hash/CA2/_0420_ ),
    .B1(\hash/CA2/_0452_ ),
    .C1(\hash/CA2/_1007_ ),
    .Y(\hash/CA2/_0453_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2057_  (.A(\hash/CA2/_1031_ ),
    .B(\hash/CA2/_0443_ ),
    .Y(\hash/CA2/_0454_ ));
 sky130_fd_sc_hd__o21a_1 \hash/CA2/_2058_  (.A1(\hash/CA2/_0432_ ),
    .A2(\hash/CA2/_0454_ ),
    .B1(\hash/CA2/_0451_ ),
    .X(\hash/CA2/_0455_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_2059_  (.A(\hash/CA2/_0453_ ),
    .B(\hash/CA2/_0455_ ),
    .Y(\hash/CA2/_0456_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2060_  (.A1(\hash/CA2/_1037_ ),
    .A2(\hash/CA2/_0456_ ),
    .B1(\hash/CA2/_1036_ ),
    .X(\hash/CA2/_0457_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_2061_  (.A(\hash/CA2/_1043_ ),
    .B(\hash/CA2/_0457_ ),
    .X(\hash/e_new[20] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2062_  (.A(\hash/CA2/_1031_ ),
    .B(\hash/CA2/_1037_ ),
    .Y(\hash/CA2/_0458_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2063_  (.A1(\hash/CA2/_0445_ ),
    .A2(\hash/CA2/_0448_ ),
    .B1(\hash/CA2/_0458_ ),
    .Y(\hash/CA2/_0459_ ));
 sky130_fd_sc_hd__a211o_1 \hash/CA2/_2064_  (.A1(\hash/CA2/_1037_ ),
    .A2(\hash/CA2/_1030_ ),
    .B1(\hash/CA2/_1036_ ),
    .C1(\hash/CA2/_0459_ ),
    .X(\hash/CA2/_0460_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2065_  (.A1(\hash/CA2/_1043_ ),
    .A2(\hash/CA2/_0460_ ),
    .B1(\hash/CA2/_1042_ ),
    .Y(\hash/CA2/_0461_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2066_  (.A(\hash/CA2/_1049_ ),
    .B(\hash/CA2/_0461_ ),
    .Y(\hash/e_new[21] ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_2067_  (.A(\hash/CA2/_1037_ ),
    .B(\hash/CA2/_1043_ ),
    .C(\hash/CA2/_1049_ ),
    .X(\hash/CA2/_0462_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2068_  (.A1(\hash/CA2/_1049_ ),
    .A2(\hash/CA2/_1042_ ),
    .B1(\hash/CA2/_1048_ ),
    .Y(\hash/CA2/_0463_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_2069_  (.A(\hash/CA2/_1043_ ),
    .B(\hash/CA2/_1049_ ),
    .X(\hash/CA2/_0464_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2070_  (.A(\hash/CA2/_1036_ ),
    .B(\hash/CA2/_0464_ ),
    .Y(\hash/CA2/_0465_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2071_  (.A(\hash/CA2/_0463_ ),
    .B(\hash/CA2/_0465_ ),
    .Y(\hash/CA2/_0466_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2072_  (.A1(\hash/CA2/_0456_ ),
    .A2(\hash/CA2/_0462_ ),
    .B1(\hash/CA2/_0466_ ),
    .Y(\hash/CA2/_0467_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2073_  (.A(\hash/CA2/_1055_ ),
    .B(\hash/CA2/_0467_ ),
    .Y(\hash/e_new[22] ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2074_  (.A(\hash/CA2/_0460_ ),
    .B(\hash/CA2/_0464_ ),
    .Y(\hash/CA2/_0468_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2075_  (.A(\hash/CA2/_0463_ ),
    .B(\hash/CA2/_0468_ ),
    .Y(\hash/CA2/_0469_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2076_  (.A1(\hash/CA2/_1055_ ),
    .A2(\hash/CA2/_0469_ ),
    .B1(\hash/CA2/_1054_ ),
    .Y(\hash/CA2/_0470_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2077_  (.A(\hash/CA2/_1061_ ),
    .B(\hash/CA2/_0470_ ),
    .Y(\hash/e_new[23] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_2078_  (.A(\hash/CA2/_1067_ ),
    .Y(\hash/CA2/_0471_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2079_  (.A(\hash/CA2/_1055_ ),
    .B(\hash/CA2/_1061_ ),
    .Y(\hash/CA2/_0472_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2080_  (.A1(\hash/CA2/_1061_ ),
    .A2(\hash/CA2/_1054_ ),
    .B1(\hash/CA2/_1060_ ),
    .Y(\hash/CA2/_0473_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2081_  (.A1(\hash/CA2/_0467_ ),
    .A2(\hash/CA2/_0472_ ),
    .B1(\hash/CA2/_0473_ ),
    .Y(\hash/CA2/_0474_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2082_  (.A(\hash/CA2/_0471_ ),
    .B(\hash/CA2/_0474_ ),
    .Y(\hash/e_new[24] ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_2083_  (.A(\hash/CA2/_1055_ ),
    .B(\hash/CA2/_1061_ ),
    .X(\hash/CA2/_0475_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2084_  (.A(\hash/CA2/_1061_ ),
    .B(\hash/CA2/_1054_ ),
    .Y(\hash/CA2/_0476_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2085_  (.A1(\hash/CA2/_0463_ ),
    .A2(\hash/CA2/_0472_ ),
    .B1(\hash/CA2/_0476_ ),
    .Y(\hash/CA2/_0477_ ));
 sky130_fd_sc_hd__a311o_1 \hash/CA2/_2086_  (.A1(\hash/CA2/_0460_ ),
    .A2(\hash/CA2/_0464_ ),
    .A3(\hash/CA2/_0475_ ),
    .B1(\hash/CA2/_0477_ ),
    .C1(\hash/CA2/_1060_ ),
    .X(\hash/CA2/_0478_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2087_  (.A1(\hash/CA2/_1067_ ),
    .A2(\hash/CA2/_0478_ ),
    .B1(\hash/CA2/_1066_ ),
    .Y(\hash/CA2/_0479_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2088_  (.A(\hash/CA2/_1073_ ),
    .B(\hash/CA2/_0479_ ),
    .Y(\hash/e_new[25] ));
 sky130_fd_sc_hd__and3_1 \hash/CA2/_2089_  (.A(\hash/CA2/_1067_ ),
    .B(\hash/CA2/_1073_ ),
    .C(\hash/CA2/_0475_ ),
    .X(\hash/CA2/_0480_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA2/_2090_  (.A1(\hash/CA2/_0463_ ),
    .A2(\hash/CA2/_0465_ ),
    .B1_N(\hash/CA2/_0480_ ),
    .Y(\hash/CA2/_0481_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_2091_  (.A(\hash/CA2/_0471_ ),
    .B(\hash/CA2/_0473_ ),
    .Y(\hash/CA2/_0482_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2092_  (.A1(\hash/CA2/_1066_ ),
    .A2(\hash/CA2/_0482_ ),
    .B1(\hash/CA2/_1073_ ),
    .Y(\hash/CA2/_0483_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/CA2/_2093_  (.A_N(\hash/CA2/_1072_ ),
    .B(\hash/CA2/_0483_ ),
    .Y(\hash/CA2/_0484_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/CA2/_2094_  (.A1(\hash/CA2/_0456_ ),
    .A2(\hash/CA2/_0462_ ),
    .A3(\hash/CA2/_0480_ ),
    .B1(\hash/CA2/_0481_ ),
    .C1(\hash/CA2/_0484_ ),
    .Y(\hash/CA2/_0485_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2095_  (.A(\hash/CA2/_1079_ ),
    .B(\hash/CA2/_0485_ ),
    .Y(\hash/e_new[26] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2097_  (.A1(\hash/CA2/_0463_ ),
    .A2(\hash/CA2/_0472_ ),
    .B1(\hash/CA2/_0473_ ),
    .Y(\hash/CA2/_0487_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2098_  (.A1(\hash/CA2/_1067_ ),
    .A2(\hash/CA2/_0487_ ),
    .B1(\hash/CA2/_1066_ ),
    .X(\hash/CA2/_0488_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2099_  (.A1(\hash/CA2/_1073_ ),
    .A2(\hash/CA2/_0488_ ),
    .B1(\hash/CA2/_1072_ ),
    .X(\hash/CA2/_0489_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2100_  (.A1(\hash/CA2/_1079_ ),
    .A2(\hash/CA2/_0489_ ),
    .B1(\hash/CA2/_1078_ ),
    .Y(\hash/CA2/_0490_ ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_2101_  (.A(\hash/CA2/_0490_ ),
    .Y(\hash/CA2/_0491_ ));
 sky130_fd_sc_hd__a41o_1 \hash/CA2/_2102_  (.A1(\hash/CA2/_1079_ ),
    .A2(\hash/CA2/_0460_ ),
    .A3(\hash/CA2/_0464_ ),
    .A4(\hash/CA2/_0480_ ),
    .B1(\hash/CA2/_0491_ ),
    .X(\hash/CA2/_0492_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_2103_  (.A(\hash/CA2/_1085_ ),
    .B(\hash/CA2/_0492_ ),
    .X(\hash/e_new[27] ));
 sky130_fd_sc_hd__o2111a_1 \hash/CA2/_2104_  (.A1(\hash/CA2/_1079_ ),
    .A2(\hash/CA2/_1078_ ),
    .B1(\hash/CA2/_0464_ ),
    .C1(\hash/CA2/_0480_ ),
    .D1(\hash/CA2/_1085_ ),
    .X(\hash/CA2/_0493_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/CA2/_2105_  (.A1(\hash/CA2/_1085_ ),
    .A2(\hash/CA2/_0491_ ),
    .B1(\hash/CA2/_0493_ ),
    .B2(\hash/CA2/_0457_ ),
    .C1(\hash/CA2/_1084_ ),
    .Y(\hash/CA2/_0494_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2106_  (.A(\hash/CA2/_1090_ ),
    .B(\hash/CA2/_0494_ ),
    .Y(\hash/e_new[28] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2107_  (.A1(\hash/CA2/_1085_ ),
    .A2(\hash/CA2/_0492_ ),
    .B1(\hash/CA2/_1084_ ),
    .X(\hash/CA2/_0495_ ));
 sky130_fd_sc_hd__a21oi_2 \hash/CA2/_2108_  (.A1(\hash/CA2/_1090_ ),
    .A2(\hash/CA2/_0495_ ),
    .B1(\hash/CA2/_1089_ ),
    .Y(\hash/CA2/_0496_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2109_  (.A(\hash/CA2/_1095_ ),
    .B(\hash/CA2/_0496_ ),
    .Y(\hash/e_new[29] ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_2110_  (.A(\hash/CA2/_0870_ ),
    .B(\hash/CA2/_0942_ ),
    .X(\hash/e_new[2] ));
 sky130_fd_sc_hd__nand4_1 \hash/CA2/_2111_  (.A(\hash/CA2/_1079_ ),
    .B(\hash/CA2/_1085_ ),
    .C(\hash/CA2/_1090_ ),
    .D(\hash/CA2/_1095_ ),
    .Y(\hash/CA2/_0497_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2112_  (.A1(\hash/CA2/_1085_ ),
    .A2(\hash/CA2/_1078_ ),
    .B1(\hash/CA2/_1084_ ),
    .X(\hash/CA2/_0498_ ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2113_  (.A1(\hash/CA2/_1090_ ),
    .A2(\hash/CA2/_0498_ ),
    .B1(\hash/CA2/_1089_ ),
    .X(\hash/CA2/_0499_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2114_  (.A1(\hash/CA2/_1095_ ),
    .A2(\hash/CA2/_0499_ ),
    .B1(\hash/CA2/_1094_ ),
    .Y(\hash/CA2/_0500_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2115_  (.A1(\hash/CA2/_0485_ ),
    .A2(\hash/CA2/_0497_ ),
    .B1(\hash/CA2/_0500_ ),
    .Y(\hash/CA2/_0501_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_2116_  (.A(\hash/CA2/_1100_ ),
    .B(\hash/CA2/_0501_ ),
    .X(\hash/e_new[30] ));
 sky130_fd_sc_hd__a21o_1 \hash/CA2/_2117_  (.A1(\hash/CA2/_1090_ ),
    .A2(\hash/CA2/_1084_ ),
    .B1(\hash/CA2/_1089_ ),
    .X(\hash/CA2/_0502_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2118_  (.A1(\hash/CA2/_1095_ ),
    .A2(\hash/CA2/_0502_ ),
    .B1(\hash/CA2/_1094_ ),
    .Y(\hash/CA2/_0503_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/CA2/_2119_  (.A_N(\hash/CA2/_1099_ ),
    .B(\hash/CA2/_0503_ ),
    .C(\hash/p5_cap[31] ),
    .Y(\hash/CA2/_0504_ ));
 sky130_fd_sc_hd__nand3_1 \hash/CA2/_2120_  (.A(\hash/CA2/_1085_ ),
    .B(\hash/CA2/_1090_ ),
    .C(\hash/CA2/_1095_ ),
    .Y(\hash/CA2/_0505_ ));
 sky130_fd_sc_hd__nor3b_1 \hash/CA2/_2121_  (.A(\hash/CA2/_0505_ ),
    .B(\hash/p5_cap[31] ),
    .C_N(\hash/CA2/_1100_ ),
    .Y(\hash/CA2/_0506_ ));
 sky130_fd_sc_hd__nand2_1 \hash/CA2/_2122_  (.A(\hash/CA2/_0492_ ),
    .B(\hash/CA2/_0506_ ),
    .Y(\hash/CA2/_0507_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_2123_  (.A(\hash/CA2/_0503_ ),
    .B_N(\hash/CA2/_1100_ ),
    .Y(\hash/CA2/_0508_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/CA2/_2124_  (.A1(\hash/CA2/_0505_ ),
    .A2(\hash/CA2/_0503_ ),
    .B1_N(\hash/CA2/_1100_ ),
    .Y(\hash/CA2/_0509_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2125_  (.A1(\hash/CA2/_1099_ ),
    .A2(\hash/CA2/_0509_ ),
    .B1(\hash/p5_cap[31] ),
    .Y(\hash/CA2/_0510_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/CA2/_2126_  (.A1(\hash/p5_cap[31] ),
    .A2(\hash/CA2/_1099_ ),
    .A3(\hash/CA2/_0508_ ),
    .B1(\hash/CA2/_0510_ ),
    .Y(\hash/CA2/_0511_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/CA2/_2127_  (.A1(\hash/CA2/_0492_ ),
    .A2(\hash/CA2/_0504_ ),
    .B1(\hash/CA2/_0507_ ),
    .C1(\hash/CA2/_0511_ ),
    .Y(\hash/CA2/_0512_ ));
 sky130_fd_sc_hd__xor2_1 \hash/CA2/_2128_  (.A(\hash/CA2/_0369_ ),
    .B(\hash/CA2/_0512_ ),
    .X(\hash/e_new[31] ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2129_  (.A1(\hash/CA2/_0942_ ),
    .A2(\hash/CA2/_0407_ ),
    .B1(\hash/CA2/_0941_ ),
    .Y(\hash/CA2/_0513_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2130_  (.A(\hash/CA2/_0947_ ),
    .B(\hash/CA2/_0513_ ),
    .Y(\hash/e_new[3] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2131_  (.A(\hash/CA2/_0952_ ),
    .B(\hash/CA2/_0399_ ),
    .Y(\hash/e_new[4] ));
 sky130_fd_sc_hd__a31o_2 \hash/CA2/_2132_  (.A1(\hash/CA2/_0942_ ),
    .A2(\hash/CA2/_0947_ ),
    .A3(\hash/CA2/_0407_ ),
    .B1(\hash/CA2/_0408_ ),
    .X(\hash/CA2/_0514_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2133_  (.A1(\hash/CA2/_0952_ ),
    .A2(\hash/CA2/_0514_ ),
    .B1(\hash/CA2/_0951_ ),
    .Y(\hash/CA2/_0515_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2134_  (.A(\hash/CA2/_0957_ ),
    .B(\hash/CA2/_0515_ ),
    .Y(\hash/e_new[5] ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2135_  (.A(\hash/CA2/_0962_ ),
    .B(\hash/CA2/_0401_ ),
    .Y(\hash/e_new[6] ));
 sky130_fd_sc_hd__inv_1 \hash/CA2/_2136_  (.A(\hash/CA2/_0961_ ),
    .Y(\hash/CA2/_0516_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/CA2/_2137_  (.A(\hash/CA2/_0515_ ),
    .B_N(\hash/CA2/_0957_ ),
    .Y(\hash/CA2/_0517_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2138_  (.A1(\hash/CA2/_0956_ ),
    .A2(\hash/CA2/_0517_ ),
    .B1(\hash/CA2/_0962_ ),
    .Y(\hash/CA2/_0518_ ));
 sky130_fd_sc_hd__and2_1 \hash/CA2/_2139_  (.A(\hash/CA2/_0516_ ),
    .B(\hash/CA2/_0518_ ),
    .X(\hash/CA2/_0519_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2140_  (.A(\hash/CA2/_0967_ ),
    .B(\hash/CA2/_0519_ ),
    .Y(\hash/e_new[7] ));
 sky130_fd_sc_hd__o21ai_0 \hash/CA2/_2141_  (.A1(\hash/CA2/_0396_ ),
    .A2(\hash/CA2/_0401_ ),
    .B1(\hash/CA2/_0516_ ),
    .Y(\hash/CA2/_0520_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/CA2/_2142_  (.A1(\hash/CA2/_0967_ ),
    .A2(\hash/CA2/_0520_ ),
    .B1(\hash/CA2/_0966_ ),
    .Y(\hash/CA2/_0521_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/CA2/_2143_  (.A(\hash/CA2/_0972_ ),
    .B(\hash/CA2/_0521_ ),
    .Y(\hash/e_new[8] ));
 sky130_fd_sc_hd__nor3_1 \hash/CA2/_2144_  (.A(\hash/CA2/_0978_ ),
    .B(\hash/CA2/_0971_ ),
    .C(\hash/CA2/_0411_ ),
    .Y(\hash/CA2/_0522_ ));
 sky130_fd_sc_hd__nor2_1 \hash/CA2/_2145_  (.A(\hash/CA2/_0412_ ),
    .B(\hash/CA2/_0522_ ),
    .Y(\hash/e_new[9] ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2146_  (.A(\hash/CA2/_0610_ ),
    .B(\hash/CA2/_0611_ ),
    .CIN(\hash/CA2/_0612_ ),
    .COUT(\hash/CA2/_0613_ ),
    .SUM(\hash/CA2/_0614_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2147_  (.A(\hash/CA2/s1[1] ),
    .B(\hash/CA2/_0615_ ),
    .CIN(\hash/CA2/_0616_ ),
    .COUT(\hash/CA2/_0617_ ),
    .SUM(\hash/CA2/_0618_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2148_  (.A(\hash/CA2/_0619_ ),
    .B(\hash/CA2/_0620_ ),
    .CIN(\hash/CA2/_0621_ ),
    .COUT(\hash/CA2/_0622_ ),
    .SUM(\hash/CA2/_0623_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2149_  (.A(\hash/CA2/_0624_ ),
    .B(\hash/CA2/_0625_ ),
    .CIN(\hash/CA2/_0626_ ),
    .COUT(\hash/CA2/_0627_ ),
    .SUM(\hash/CA2/_0628_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2150_  (.A(\hash/CA2/_0629_ ),
    .B(\hash/CA2/_0622_ ),
    .CIN(\hash/CA2/_0628_ ),
    .COUT(\hash/CA2/_0630_ ),
    .SUM(\hash/CA2/_0631_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2151_  (.A(\hash/CA2/_0632_ ),
    .B(\hash/CA2/_0633_ ),
    .CIN(\hash/CA2/_0634_ ),
    .COUT(\hash/CA2/_0635_ ),
    .SUM(\hash/CA2/_0636_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2152_  (.A(\hash/CA2/_0627_ ),
    .B(\hash/CA2/_0636_ ),
    .CIN(\hash/CA2/_0637_ ),
    .COUT(\hash/CA2/_0638_ ),
    .SUM(\hash/CA2/_0639_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2153_  (.A(\hash/CA2/_0641_ ),
    .B(\hash/CA2/_0642_ ),
    .CIN(\hash/CA2/_0643_ ),
    .COUT(\hash/CA2/_0644_ ),
    .SUM(\hash/CA2/_0645_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2154_  (.A(\hash/CA2/_0635_ ),
    .B(\hash/CA2/_0645_ ),
    .CIN(\hash/CA2/_0646_ ),
    .COUT(\hash/CA2/_0647_ ),
    .SUM(\hash/CA2/_0648_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2155_  (.A(\hash/CA2/_0650_ ),
    .B(\hash/CA2/_0651_ ),
    .CIN(\hash/CA2/_0652_ ),
    .COUT(\hash/CA2/_0653_ ),
    .SUM(\hash/CA2/_0654_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2156_  (.A(\hash/CA2/_0644_ ),
    .B(\hash/CA2/_0654_ ),
    .CIN(\hash/CA2/_0655_ ),
    .COUT(\hash/CA2/_0656_ ),
    .SUM(\hash/CA2/_0657_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2157_  (.A(\hash/p4_cap[5] ),
    .B(\hash/CA2/s0[5] ),
    .CIN(\hash/CA2/_0659_ ),
    .COUT(\hash/CA2/_0660_ ),
    .SUM(\hash/CA2/_0661_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2158_  (.A(\hash/CA2/_0662_ ),
    .B(\hash/CA2/_0661_ ),
    .CIN(\hash/CA2/_0663_ ),
    .COUT(\hash/CA2/_0664_ ),
    .SUM(\hash/CA2/_0665_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2159_  (.A(\hash/p4_cap[6] ),
    .B(\hash/CA2/s0[6] ),
    .CIN(\hash/CA2/_0666_ ),
    .COUT(\hash/CA2/_0667_ ),
    .SUM(\hash/CA2/_0668_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2160_  (.A(\hash/CA2/_0668_ ),
    .B(\hash/CA2/_0660_ ),
    .CIN(\hash/CA2/_0669_ ),
    .COUT(\hash/CA2/_0670_ ),
    .SUM(\hash/CA2/_0671_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2161_  (.A(\hash/p4_cap[7] ),
    .B(\hash/CA2/s0[7] ),
    .CIN(\hash/CA2/_0672_ ),
    .COUT(\hash/CA2/_0673_ ),
    .SUM(\hash/CA2/_0674_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2162_  (.A(\hash/CA2/_0667_ ),
    .B(\hash/CA2/_0674_ ),
    .CIN(\hash/CA2/_0675_ ),
    .COUT(\hash/CA2/_0676_ ),
    .SUM(\hash/CA2/_0677_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2163_  (.A(\hash/CA2/_0678_ ),
    .B(\hash/CA2/_0679_ ),
    .CIN(\hash/CA2/_0680_ ),
    .COUT(\hash/CA2/_0681_ ),
    .SUM(\hash/CA2/_0682_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2164_  (.A(\hash/CA2/_0683_ ),
    .B(\hash/CA2/_0682_ ),
    .CIN(\hash/CA2/_0684_ ),
    .COUT(\hash/CA2/_0685_ ),
    .SUM(\hash/CA2/_0686_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2165_  (.A(\hash/CA2/_0688_ ),
    .B(\hash/CA2/_0689_ ),
    .CIN(\hash/CA2/_0690_ ),
    .COUT(\hash/CA2/_0691_ ),
    .SUM(\hash/CA2/_0692_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2166_  (.A(\hash/CA2/_0681_ ),
    .B(\hash/CA2/_0692_ ),
    .CIN(\hash/CA2/_0693_ ),
    .COUT(\hash/CA2/_0694_ ),
    .SUM(\hash/CA2/_0695_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2167_  (.A(\hash/CA2/_0696_ ),
    .B(\hash/CA2/_0697_ ),
    .CIN(\hash/CA2/_0698_ ),
    .COUT(\hash/CA2/_0699_ ),
    .SUM(\hash/CA2/_0700_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2168_  (.A(\hash/CA2/_0691_ ),
    .B(\hash/CA2/_0700_ ),
    .CIN(\hash/CA2/_0701_ ),
    .COUT(\hash/CA2/_0702_ ),
    .SUM(\hash/CA2/_0703_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2169_  (.A(\hash/CA2/_0704_ ),
    .B(\hash/CA2/_0705_ ),
    .CIN(\hash/CA2/_0706_ ),
    .COUT(\hash/CA2/_0707_ ),
    .SUM(\hash/CA2/_0708_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2170_  (.A(\hash/CA2/_0699_ ),
    .B(\hash/CA2/_0708_ ),
    .CIN(\hash/CA2/_0709_ ),
    .COUT(\hash/CA2/_0710_ ),
    .SUM(\hash/CA2/_0711_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2171_  (.A(\hash/CA2/_0712_ ),
    .B(\hash/CA2/_0713_ ),
    .CIN(\hash/CA2/_0714_ ),
    .COUT(\hash/CA2/_0715_ ),
    .SUM(\hash/CA2/_0716_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2172_  (.A(\hash/CA2/_0707_ ),
    .B(\hash/CA2/_0716_ ),
    .CIN(\hash/CA2/_0717_ ),
    .COUT(\hash/CA2/_0718_ ),
    .SUM(\hash/CA2/_0719_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2173_  (.A(\hash/CA2/_0720_ ),
    .B(\hash/CA2/_0721_ ),
    .CIN(\hash/CA2/_0722_ ),
    .COUT(\hash/CA2/_0723_ ),
    .SUM(\hash/CA2/_0724_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2174_  (.A(\hash/CA2/_0715_ ),
    .B(\hash/CA2/_0724_ ),
    .CIN(\hash/CA2/_0725_ ),
    .COUT(\hash/CA2/_0726_ ),
    .SUM(\hash/CA2/_0727_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2175_  (.A(\hash/CA2/_0728_ ),
    .B(\hash/CA2/_0729_ ),
    .CIN(\hash/CA2/_0730_ ),
    .COUT(\hash/CA2/_0731_ ),
    .SUM(\hash/CA2/_0732_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2176_  (.A(\hash/CA2/_0723_ ),
    .B(\hash/CA2/_0732_ ),
    .CIN(\hash/CA2/_0733_ ),
    .COUT(\hash/CA2/_0734_ ),
    .SUM(\hash/CA2/_0735_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2177_  (.A(\hash/CA2/_0736_ ),
    .B(\hash/CA2/_0737_ ),
    .CIN(\hash/CA2/_0738_ ),
    .COUT(\hash/CA2/_0739_ ),
    .SUM(\hash/CA2/_0740_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2178_  (.A(\hash/CA2/_0731_ ),
    .B(\hash/CA2/_0740_ ),
    .CIN(\hash/CA2/_0741_ ),
    .COUT(\hash/CA2/_0742_ ),
    .SUM(\hash/CA2/_0743_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2179_  (.A(\hash/CA2/_0744_ ),
    .B(\hash/CA2/_0745_ ),
    .CIN(\hash/CA2/_0746_ ),
    .COUT(\hash/CA2/_0747_ ),
    .SUM(\hash/CA2/_0748_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2180_  (.A(\hash/CA2/_0739_ ),
    .B(\hash/CA2/_0748_ ),
    .CIN(\hash/CA2/_0749_ ),
    .COUT(\hash/CA2/_0750_ ),
    .SUM(\hash/CA2/_0751_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2181_  (.A(\hash/CA2/_0753_ ),
    .B(\hash/CA2/_0754_ ),
    .CIN(\hash/CA2/_0755_ ),
    .COUT(\hash/CA2/_0756_ ),
    .SUM(\hash/CA2/_0757_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2182_  (.A(\hash/CA2/_0747_ ),
    .B(\hash/CA2/_0757_ ),
    .CIN(\hash/CA2/_0758_ ),
    .COUT(\hash/CA2/_0759_ ),
    .SUM(\hash/CA2/_0760_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2183_  (.A(\hash/CA2/_0761_ ),
    .B(\hash/CA2/_0762_ ),
    .CIN(\hash/CA2/_0763_ ),
    .COUT(\hash/CA2/_0764_ ),
    .SUM(\hash/CA2/_0765_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2184_  (.A(\hash/CA2/_0765_ ),
    .B(\hash/CA2/_0756_ ),
    .CIN(\hash/CA2/_0766_ ),
    .COUT(\hash/CA2/_0767_ ),
    .SUM(\hash/CA2/_0768_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2185_  (.A(\hash/CA2/_0769_ ),
    .B(\hash/CA2/_0770_ ),
    .CIN(\hash/CA2/_0771_ ),
    .COUT(\hash/CA2/_0772_ ),
    .SUM(\hash/CA2/_0773_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2186_  (.A(\hash/CA2/_0764_ ),
    .B(\hash/CA2/_0773_ ),
    .CIN(\hash/CA2/_0774_ ),
    .COUT(\hash/CA2/_0775_ ),
    .SUM(\hash/CA2/_0776_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2187_  (.A(\hash/CA2/_0777_ ),
    .B(\hash/CA2/_0778_ ),
    .CIN(\hash/CA2/_0779_ ),
    .COUT(\hash/CA2/_0780_ ),
    .SUM(\hash/CA2/_0781_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2188_  (.A(\hash/CA2/_0772_ ),
    .B(\hash/CA2/_0781_ ),
    .CIN(\hash/CA2/_0782_ ),
    .COUT(\hash/CA2/_0783_ ),
    .SUM(\hash/CA2/_0784_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2189_  (.A(\hash/CA2/_0785_ ),
    .B(\hash/CA2/_0786_ ),
    .CIN(\hash/CA2/_0787_ ),
    .COUT(\hash/CA2/_0788_ ),
    .SUM(\hash/CA2/_0789_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2190_  (.A(\hash/CA2/_0789_ ),
    .B(\hash/CA2/_0780_ ),
    .CIN(\hash/CA2/_0790_ ),
    .COUT(\hash/CA2/_0791_ ),
    .SUM(\hash/CA2/_0792_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2191_  (.A(\hash/CA2/_0793_ ),
    .B(\hash/CA2/_0794_ ),
    .CIN(\hash/CA2/_0795_ ),
    .COUT(\hash/CA2/_0796_ ),
    .SUM(\hash/CA2/_0797_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2192_  (.A(\hash/CA2/_0788_ ),
    .B(\hash/CA2/_0797_ ),
    .CIN(\hash/CA2/_0798_ ),
    .COUT(\hash/CA2/_0799_ ),
    .SUM(\hash/CA2/_0800_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2193_  (.A(\hash/CA2/_0801_ ),
    .B(\hash/CA2/_0802_ ),
    .CIN(\hash/CA2/_0803_ ),
    .COUT(\hash/CA2/_0804_ ),
    .SUM(\hash/CA2/_0805_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2194_  (.A(\hash/CA2/_0796_ ),
    .B(\hash/CA2/_0805_ ),
    .CIN(\hash/CA2/_0806_ ),
    .COUT(\hash/CA2/_0807_ ),
    .SUM(\hash/CA2/_0808_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2195_  (.A(\hash/CA2/_0809_ ),
    .B(\hash/CA2/_0810_ ),
    .CIN(\hash/CA2/_0811_ ),
    .COUT(\hash/CA2/_0812_ ),
    .SUM(\hash/CA2/_0813_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2196_  (.A(\hash/CA2/_0804_ ),
    .B(\hash/CA2/_0813_ ),
    .CIN(\hash/CA2/_0814_ ),
    .COUT(\hash/CA2/_0815_ ),
    .SUM(\hash/CA2/_0816_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2197_  (.A(\hash/CA2/_0817_ ),
    .B(\hash/CA2/_0818_ ),
    .CIN(\hash/CA2/_0819_ ),
    .COUT(\hash/CA2/_0820_ ),
    .SUM(\hash/CA2/_0821_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2198_  (.A(\hash/CA2/_0812_ ),
    .B(\hash/CA2/_0821_ ),
    .CIN(\hash/CA2/_0822_ ),
    .COUT(\hash/CA2/_0823_ ),
    .SUM(\hash/CA2/_0824_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2199_  (.A(\hash/CA2/_0825_ ),
    .B(\hash/CA2/_0826_ ),
    .CIN(\hash/CA2/_0827_ ),
    .COUT(\hash/CA2/_0828_ ),
    .SUM(\hash/CA2/_0829_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2200_  (.A(\hash/CA2/_0820_ ),
    .B(\hash/CA2/_0829_ ),
    .CIN(\hash/CA2/_0830_ ),
    .COUT(\hash/CA2/_0831_ ),
    .SUM(\hash/CA2/_0832_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2201_  (.A(\hash/CA2/_0833_ ),
    .B(\hash/CA2/_0834_ ),
    .CIN(\hash/CA2/_0835_ ),
    .COUT(\hash/CA2/_0836_ ),
    .SUM(\hash/CA2/_0837_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2202_  (.A(\hash/CA2/_0828_ ),
    .B(\hash/CA2/_0837_ ),
    .CIN(\hash/CA2/_0838_ ),
    .COUT(\hash/CA2/_0839_ ),
    .SUM(\hash/CA2/_0840_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2203_  (.A(\hash/CA2/_0841_ ),
    .B(\hash/CA2/_0842_ ),
    .CIN(\hash/CA2/_0843_ ),
    .COUT(\hash/CA2/_0844_ ),
    .SUM(\hash/CA2/_0845_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2204_  (.A(\hash/CA2/_0836_ ),
    .B(\hash/CA2/_0845_ ),
    .CIN(\hash/CA2/_0846_ ),
    .COUT(\hash/CA2/_0847_ ),
    .SUM(\hash/CA2/_0848_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2205_  (.A(\hash/CA2/_0850_ ),
    .B(\hash/CA2/_0851_ ),
    .CIN(\hash/CA2/_0852_ ),
    .COUT(\hash/CA2/_0853_ ),
    .SUM(\hash/CA2/_0854_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2206_  (.A(\hash/CA2/_0844_ ),
    .B(\hash/CA2/_0854_ ),
    .CIN(\hash/CA2/_0855_ ),
    .COUT(\hash/CA2/_0856_ ),
    .SUM(\hash/CA2/_0857_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2207_  (.A(\hash/p4_cap[30] ),
    .B(\hash/CA2/s0[30] ),
    .CIN(\hash/CA2/_0859_ ),
    .COUT(\hash/CA2/_0860_ ),
    .SUM(\hash/CA2/_0861_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2208_  (.A(\hash/CA2/_0862_ ),
    .B(\hash/CA2/_0861_ ),
    .CIN(\hash/CA2/_0863_ ),
    .COUT(\hash/CA2/_0864_ ),
    .SUM(\hash/CA2/_0865_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2209_  (.A(\hash/CA2/_0866_ ),
    .B(\hash/CA2/_0630_ ),
    .CIN(\hash/CA2/_0639_ ),
    .COUT(\hash/CA2/_0867_ ),
    .SUM(\hash/CA2/_0868_ ));
 sky130_fd_sc_hd__fa_1 \hash/CA2/_2210_  (.A(\hash/p5_cap[1] ),
    .B(\hash/CA2/_0869_ ),
    .CIN(\hash/CA2/_0618_ ),
    .COUT(\hash/CA2/_0870_ ),
    .SUM(\hash/e_new[1] ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2211_  (.A(\hash/p1_cap[0] ),
    .B(\hash/p3_cap[0] ),
    .COUT(\hash/CA2/_0871_ ),
    .SUM(\hash/b_new[0] ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2212_  (.A(\hash/p1_cap[1] ),
    .B(\hash/p3_cap[1] ),
    .COUT(\hash/CA2/_0872_ ),
    .SUM(\hash/CA2/_0873_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2213_  (.A(\hash/p1_cap[2] ),
    .B(\hash/p3_cap[2] ),
    .COUT(\hash/CA2/_0874_ ),
    .SUM(\hash/CA2/_0875_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2214_  (.A(\hash/p1_cap[3] ),
    .B(\hash/p3_cap[3] ),
    .COUT(\hash/CA2/_0876_ ),
    .SUM(\hash/CA2/_0877_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2215_  (.A(\hash/p1_cap[4] ),
    .B(\hash/p3_cap[4] ),
    .COUT(\hash/CA2/_0878_ ),
    .SUM(\hash/CA2/_0879_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2216_  (.A(\hash/p1_cap[5] ),
    .B(\hash/p3_cap[5] ),
    .COUT(\hash/CA2/_0880_ ),
    .SUM(\hash/CA2/_0881_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2217_  (.A(\hash/p1_cap[6] ),
    .B(\hash/p3_cap[6] ),
    .COUT(\hash/CA2/_0882_ ),
    .SUM(\hash/CA2/_0883_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2218_  (.A(\hash/p1_cap[7] ),
    .B(\hash/p3_cap[7] ),
    .COUT(\hash/CA2/_0884_ ),
    .SUM(\hash/CA2/_0885_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2219_  (.A(\hash/p1_cap[8] ),
    .B(\hash/p3_cap[8] ),
    .COUT(\hash/CA2/_0886_ ),
    .SUM(\hash/CA2/_0887_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2220_  (.A(\hash/p1_cap[9] ),
    .B(\hash/p3_cap[9] ),
    .COUT(\hash/CA2/_0888_ ),
    .SUM(\hash/CA2/_0889_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2221_  (.A(\hash/p1_cap[10] ),
    .B(\hash/p3_cap[10] ),
    .COUT(\hash/CA2/_0890_ ),
    .SUM(\hash/CA2/_0891_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2222_  (.A(\hash/p1_cap[11] ),
    .B(\hash/p3_cap[11] ),
    .COUT(\hash/CA2/_0892_ ),
    .SUM(\hash/CA2/_0893_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2223_  (.A(\hash/p1_cap[12] ),
    .B(\hash/p3_cap[12] ),
    .COUT(\hash/CA2/_0894_ ),
    .SUM(\hash/CA2/_0895_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2224_  (.A(\hash/p1_cap[13] ),
    .B(\hash/p3_cap[13] ),
    .COUT(\hash/CA2/_0896_ ),
    .SUM(\hash/CA2/_0897_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2225_  (.A(\hash/p1_cap[14] ),
    .B(\hash/p3_cap[14] ),
    .COUT(\hash/CA2/_0898_ ),
    .SUM(\hash/CA2/_0899_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2226_  (.A(\hash/p1_cap[15] ),
    .B(\hash/p3_cap[15] ),
    .COUT(\hash/CA2/_0900_ ),
    .SUM(\hash/CA2/_0901_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2227_  (.A(\hash/p1_cap[16] ),
    .B(\hash/p3_cap[16] ),
    .COUT(\hash/CA2/_0902_ ),
    .SUM(\hash/CA2/_0903_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2228_  (.A(\hash/p1_cap[17] ),
    .B(\hash/p3_cap[17] ),
    .COUT(\hash/CA2/_0904_ ),
    .SUM(\hash/CA2/_0905_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2229_  (.A(\hash/p1_cap[18] ),
    .B(\hash/p3_cap[18] ),
    .COUT(\hash/CA2/_0906_ ),
    .SUM(\hash/CA2/_0907_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2230_  (.A(\hash/p1_cap[19] ),
    .B(\hash/p3_cap[19] ),
    .COUT(\hash/CA2/_0908_ ),
    .SUM(\hash/CA2/_0909_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2231_  (.A(\hash/p1_cap[20] ),
    .B(\hash/p3_cap[20] ),
    .COUT(\hash/CA2/_0910_ ),
    .SUM(\hash/CA2/_0911_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2232_  (.A(\hash/p1_cap[21] ),
    .B(\hash/p3_cap[21] ),
    .COUT(\hash/CA2/_0912_ ),
    .SUM(\hash/CA2/_0913_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2233_  (.A(\hash/p1_cap[22] ),
    .B(\hash/p3_cap[22] ),
    .COUT(\hash/CA2/_0914_ ),
    .SUM(\hash/CA2/_0915_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2234_  (.A(\hash/p1_cap[23] ),
    .B(\hash/p3_cap[23] ),
    .COUT(\hash/CA2/_0916_ ),
    .SUM(\hash/CA2/_0917_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2235_  (.A(\hash/p1_cap[24] ),
    .B(\hash/p3_cap[24] ),
    .COUT(\hash/CA2/_0918_ ),
    .SUM(\hash/CA2/_0919_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2236_  (.A(\hash/p1_cap[25] ),
    .B(\hash/p3_cap[25] ),
    .COUT(\hash/CA2/_0920_ ),
    .SUM(\hash/CA2/_0921_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2237_  (.A(\hash/p1_cap[26] ),
    .B(\hash/p3_cap[26] ),
    .COUT(\hash/CA2/_0922_ ),
    .SUM(\hash/CA2/_0923_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2238_  (.A(\hash/p1_cap[27] ),
    .B(\hash/p3_cap[27] ),
    .COUT(\hash/CA2/_0924_ ),
    .SUM(\hash/CA2/_0925_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2239_  (.A(\hash/p1_cap[28] ),
    .B(\hash/p3_cap[28] ),
    .COUT(\hash/CA2/_0926_ ),
    .SUM(\hash/CA2/_0927_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2240_  (.A(\hash/p1_cap[29] ),
    .B(\hash/p3_cap[29] ),
    .COUT(\hash/CA2/_0928_ ),
    .SUM(\hash/CA2/_0929_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2241_  (.A(\hash/p1_cap[30] ),
    .B(\hash/p3_cap[30] ),
    .COUT(\hash/CA2/_0930_ ),
    .SUM(\hash/CA2/_0931_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2242_  (.A(\hash/CA2/s1[0] ),
    .B(\hash/CA2/_0932_ ),
    .COUT(\hash/CA2/_0615_ ),
    .SUM(\hash/CA2/_0933_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2243_  (.A(\hash/CA2/s1[1] ),
    .B(\hash/CA2/_0616_ ),
    .COUT(\hash/CA2/_0934_ ),
    .SUM(\hash/CA2/_0935_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2244_  (.A(\hash/p5_cap[1] ),
    .B(\hash/CA2/_0618_ ),
    .COUT(\hash/CA2/_0936_ ),
    .SUM(\hash/CA2/_0937_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2245_  (.A(\hash/CA2/s1[2] ),
    .B(\hash/CA2/_0938_ ),
    .COUT(\hash/CA2/_0939_ ),
    .SUM(\hash/CA2/_0940_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2246_  (.A(\hash/p5_cap[2] ),
    .B(\hash/CA2/_0640_ ),
    .COUT(\hash/CA2/_0941_ ),
    .SUM(\hash/CA2/_0942_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2247_  (.A(\hash/CA2/s1[3] ),
    .B(\hash/CA2/_0943_ ),
    .COUT(\hash/CA2/_0944_ ),
    .SUM(\hash/CA2/_0945_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2248_  (.A(\hash/p5_cap[3] ),
    .B(\hash/CA2/_0649_ ),
    .COUT(\hash/CA2/_0946_ ),
    .SUM(\hash/CA2/_0947_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2249_  (.A(\hash/CA2/s1[4] ),
    .B(\hash/CA2/_0948_ ),
    .COUT(\hash/CA2/_0949_ ),
    .SUM(\hash/CA2/_0950_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2250_  (.A(\hash/p5_cap[4] ),
    .B(\hash/CA2/_0658_ ),
    .COUT(\hash/CA2/_0951_ ),
    .SUM(\hash/CA2/_0952_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2251_  (.A(\hash/CA2/s1[5] ),
    .B(\hash/CA2/_0953_ ),
    .COUT(\hash/CA2/_0954_ ),
    .SUM(\hash/CA2/_0955_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2252_  (.A(\hash/p5_cap[5] ),
    .B(\hash/CA2/_0663_ ),
    .COUT(\hash/CA2/_0956_ ),
    .SUM(\hash/CA2/_0957_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2253_  (.A(\hash/CA2/s1[6] ),
    .B(\hash/CA2/_0958_ ),
    .COUT(\hash/CA2/_0959_ ),
    .SUM(\hash/CA2/_0960_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2254_  (.A(\hash/p5_cap[6] ),
    .B(\hash/CA2/_0669_ ),
    .COUT(\hash/CA2/_0961_ ),
    .SUM(\hash/CA2/_0962_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2255_  (.A(\hash/CA2/s1[7] ),
    .B(\hash/CA2/_0963_ ),
    .COUT(\hash/CA2/_0964_ ),
    .SUM(\hash/CA2/_0965_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2256_  (.A(\hash/p5_cap[7] ),
    .B(\hash/CA2/_0675_ ),
    .COUT(\hash/CA2/_0966_ ),
    .SUM(\hash/CA2/_0967_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2257_  (.A(\hash/CA2/s1[8] ),
    .B(\hash/CA2/_0968_ ),
    .COUT(\hash/CA2/_0969_ ),
    .SUM(\hash/CA2/_0970_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2258_  (.A(\hash/p5_cap[8] ),
    .B(\hash/CA2/_0687_ ),
    .COUT(\hash/CA2/_0971_ ),
    .SUM(\hash/CA2/_0972_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2259_  (.A(\hash/CA2/s1[9] ),
    .B(\hash/CA2/_0973_ ),
    .COUT(\hash/CA2/_0974_ ),
    .SUM(\hash/CA2/_0975_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2260_  (.A(\hash/p5_cap[9] ),
    .B(\hash/CA2/_0976_ ),
    .COUT(\hash/CA2/_0977_ ),
    .SUM(\hash/CA2/_0978_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2261_  (.A(\hash/CA2/s1[10] ),
    .B(\hash/CA2/_0979_ ),
    .COUT(\hash/CA2/_0980_ ),
    .SUM(\hash/CA2/_0981_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2262_  (.A(\hash/p5_cap[10] ),
    .B(\hash/CA2/_0982_ ),
    .COUT(\hash/CA2/_0983_ ),
    .SUM(\hash/CA2/_0984_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2263_  (.A(\hash/CA2/s1[11] ),
    .B(\hash/CA2/_0985_ ),
    .COUT(\hash/CA2/_0986_ ),
    .SUM(\hash/CA2/_0987_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2264_  (.A(\hash/p5_cap[11] ),
    .B(\hash/CA2/_0988_ ),
    .COUT(\hash/CA2/_0989_ ),
    .SUM(\hash/CA2/_0990_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2265_  (.A(\hash/CA2/s1[12] ),
    .B(\hash/CA2/_0991_ ),
    .COUT(\hash/CA2/_0992_ ),
    .SUM(\hash/CA2/_0993_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2266_  (.A(\hash/p5_cap[12] ),
    .B(\hash/CA2/_0994_ ),
    .COUT(\hash/CA2/_0995_ ),
    .SUM(\hash/CA2/_0996_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2267_  (.A(\hash/CA2/s1[13] ),
    .B(\hash/CA2/_0997_ ),
    .COUT(\hash/CA2/_0998_ ),
    .SUM(\hash/CA2/_0999_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2268_  (.A(\hash/p5_cap[13] ),
    .B(\hash/CA2/_1000_ ),
    .COUT(\hash/CA2/_1001_ ),
    .SUM(\hash/CA2/_1002_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2269_  (.A(\hash/CA2/s1[14] ),
    .B(\hash/CA2/_1003_ ),
    .COUT(\hash/CA2/_1004_ ),
    .SUM(\hash/CA2/_1005_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2270_  (.A(\hash/p5_cap[14] ),
    .B(\hash/CA2/_1006_ ),
    .COUT(\hash/CA2/_1007_ ),
    .SUM(\hash/CA2/_1008_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2271_  (.A(\hash/CA2/s1[15] ),
    .B(\hash/CA2/_1009_ ),
    .COUT(\hash/CA2/_1010_ ),
    .SUM(\hash/CA2/_1011_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2272_  (.A(\hash/p5_cap[15] ),
    .B(\hash/CA2/_1012_ ),
    .COUT(\hash/CA2/_1013_ ),
    .SUM(\hash/CA2/_1014_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2273_  (.A(\hash/CA2/s1[16] ),
    .B(\hash/CA2/_1015_ ),
    .COUT(\hash/CA2/_1016_ ),
    .SUM(\hash/CA2/_1017_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2274_  (.A(\hash/p5_cap[16] ),
    .B(\hash/CA2/_0752_ ),
    .COUT(\hash/CA2/_1018_ ),
    .SUM(\hash/CA2/_1019_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2275_  (.A(\hash/CA2/s1[17] ),
    .B(\hash/CA2/_1020_ ),
    .COUT(\hash/CA2/_1021_ ),
    .SUM(\hash/CA2/_1022_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2276_  (.A(\hash/p5_cap[17] ),
    .B(\hash/CA2/_1023_ ),
    .COUT(\hash/CA2/_1024_ ),
    .SUM(\hash/CA2/_1025_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2277_  (.A(\hash/CA2/s1[18] ),
    .B(\hash/CA2/_1026_ ),
    .COUT(\hash/CA2/_1027_ ),
    .SUM(\hash/CA2/_1028_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2278_  (.A(\hash/p5_cap[18] ),
    .B(\hash/CA2/_1029_ ),
    .COUT(\hash/CA2/_1030_ ),
    .SUM(\hash/CA2/_1031_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2279_  (.A(\hash/CA2/s1[19] ),
    .B(\hash/CA2/_1032_ ),
    .COUT(\hash/CA2/_1033_ ),
    .SUM(\hash/CA2/_1034_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2280_  (.A(\hash/p5_cap[19] ),
    .B(\hash/CA2/_1035_ ),
    .COUT(\hash/CA2/_1036_ ),
    .SUM(\hash/CA2/_1037_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2281_  (.A(\hash/CA2/s1[20] ),
    .B(\hash/CA2/_1038_ ),
    .COUT(\hash/CA2/_1039_ ),
    .SUM(\hash/CA2/_1040_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2282_  (.A(\hash/p5_cap[20] ),
    .B(\hash/CA2/_1041_ ),
    .COUT(\hash/CA2/_1042_ ),
    .SUM(\hash/CA2/_1043_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2283_  (.A(\hash/CA2/s1[21] ),
    .B(\hash/CA2/_1044_ ),
    .COUT(\hash/CA2/_1045_ ),
    .SUM(\hash/CA2/_1046_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2284_  (.A(\hash/p5_cap[21] ),
    .B(\hash/CA2/_1047_ ),
    .COUT(\hash/CA2/_1048_ ),
    .SUM(\hash/CA2/_1049_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2285_  (.A(\hash/CA2/s1[22] ),
    .B(\hash/CA2/_1050_ ),
    .COUT(\hash/CA2/_1051_ ),
    .SUM(\hash/CA2/_1052_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2286_  (.A(\hash/p5_cap[22] ),
    .B(\hash/CA2/_1053_ ),
    .COUT(\hash/CA2/_1054_ ),
    .SUM(\hash/CA2/_1055_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2287_  (.A(\hash/CA2/s1[23] ),
    .B(\hash/CA2/_1056_ ),
    .COUT(\hash/CA2/_1057_ ),
    .SUM(\hash/CA2/_1058_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2288_  (.A(\hash/p5_cap[23] ),
    .B(\hash/CA2/_1059_ ),
    .COUT(\hash/CA2/_1060_ ),
    .SUM(\hash/CA2/_1061_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2289_  (.A(\hash/CA2/s1[24] ),
    .B(\hash/CA2/_1062_ ),
    .COUT(\hash/CA2/_1063_ ),
    .SUM(\hash/CA2/_1064_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2290_  (.A(\hash/p5_cap[24] ),
    .B(\hash/CA2/_1065_ ),
    .COUT(\hash/CA2/_1066_ ),
    .SUM(\hash/CA2/_1067_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2291_  (.A(\hash/CA2/s1[25] ),
    .B(\hash/CA2/_1068_ ),
    .COUT(\hash/CA2/_1069_ ),
    .SUM(\hash/CA2/_1070_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2292_  (.A(\hash/p5_cap[25] ),
    .B(\hash/CA2/_1071_ ),
    .COUT(\hash/CA2/_1072_ ),
    .SUM(\hash/CA2/_1073_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2293_  (.A(\hash/CA2/s1[26] ),
    .B(\hash/CA2/_1074_ ),
    .COUT(\hash/CA2/_1075_ ),
    .SUM(\hash/CA2/_1076_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2294_  (.A(\hash/p5_cap[26] ),
    .B(\hash/CA2/_1077_ ),
    .COUT(\hash/CA2/_1078_ ),
    .SUM(\hash/CA2/_1079_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2295_  (.A(\hash/CA2/s1[27] ),
    .B(\hash/CA2/_1080_ ),
    .COUT(\hash/CA2/_1081_ ),
    .SUM(\hash/CA2/_1082_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2296_  (.A(\hash/p5_cap[27] ),
    .B(\hash/CA2/_1083_ ),
    .COUT(\hash/CA2/_1084_ ),
    .SUM(\hash/CA2/_1085_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2297_  (.A(\hash/CA2/s1[28] ),
    .B(\hash/CA2/_1086_ ),
    .COUT(\hash/CA2/_1087_ ),
    .SUM(\hash/CA2/_1088_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2298_  (.A(\hash/p5_cap[28] ),
    .B(\hash/CA2/_0849_ ),
    .COUT(\hash/CA2/_1089_ ),
    .SUM(\hash/CA2/_1090_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2299_  (.A(\hash/CA2/s1[29] ),
    .B(\hash/CA2/_1091_ ),
    .COUT(\hash/CA2/_1092_ ),
    .SUM(\hash/CA2/_1093_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2300_  (.A(\hash/p5_cap[29] ),
    .B(\hash/CA2/_0858_ ),
    .COUT(\hash/CA2/_1094_ ),
    .SUM(\hash/CA2/_1095_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2301_  (.A(\hash/CA2/s1[30] ),
    .B(\hash/CA2/_1096_ ),
    .COUT(\hash/CA2/_1097_ ),
    .SUM(\hash/CA2/_1098_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2302_  (.A(\hash/p5_cap[30] ),
    .B(\hash/CA2/_0863_ ),
    .COUT(\hash/CA2/_1099_ ),
    .SUM(\hash/CA2/_1100_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2303_  (.A(\hash/CA2/_1101_ ),
    .B(\hash/CA2/_1102_ ),
    .COUT(\hash/CA2/_1103_ ),
    .SUM(\hash/CA2/_1104_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2304_  (.A(\hash/CA2/_1105_ ),
    .B(\hash/CA2/_1106_ ),
    .COUT(\hash/CA2/_1107_ ),
    .SUM(\hash/CA2/_1108_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2305_  (.A(\hash/CA2/_1109_ ),
    .B(\hash/CA2/_1110_ ),
    .COUT(\hash/CA2/_1111_ ),
    .SUM(\hash/CA2/_1112_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2306_  (.A(\hash/CA2/_1113_ ),
    .B(\hash/CA2/_0665_ ),
    .COUT(\hash/CA2/_1114_ ),
    .SUM(\hash/CA2/_1115_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2307_  (.A(\hash/CA2/_0664_ ),
    .B(\hash/CA2/_0671_ ),
    .COUT(\hash/CA2/_1116_ ),
    .SUM(\hash/CA2/_1117_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2308_  (.A(\hash/CA2/_0670_ ),
    .B(\hash/CA2/_0677_ ),
    .COUT(\hash/CA2/_1118_ ),
    .SUM(\hash/CA2/_1119_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2309_  (.A(\hash/CA2/_0676_ ),
    .B(\hash/CA2/_1120_ ),
    .COUT(\hash/CA2/_1121_ ),
    .SUM(\hash/CA2/_1122_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2310_  (.A(\hash/CA2/_1123_ ),
    .B(\hash/CA2/_1124_ ),
    .COUT(\hash/CA2/_1125_ ),
    .SUM(\hash/CA2/_1126_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2311_  (.A(\hash/CA2/_1127_ ),
    .B(\hash/CA2/_1128_ ),
    .COUT(\hash/CA2/_1129_ ),
    .SUM(\hash/CA2/_1130_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2312_  (.A(\hash/CA2/_1131_ ),
    .B(\hash/CA2/_1132_ ),
    .COUT(\hash/CA2/_1133_ ),
    .SUM(\hash/CA2/_1134_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2313_  (.A(\hash/CA2/_1135_ ),
    .B(\hash/CA2/_1136_ ),
    .COUT(\hash/CA2/_1137_ ),
    .SUM(\hash/CA2/_1138_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2314_  (.A(\hash/CA2/_1139_ ),
    .B(\hash/CA2/_1140_ ),
    .COUT(\hash/CA2/_1141_ ),
    .SUM(\hash/CA2/_1142_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2315_  (.A(\hash/CA2/_1143_ ),
    .B(\hash/CA2/_1144_ ),
    .COUT(\hash/CA2/_1145_ ),
    .SUM(\hash/CA2/_1146_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2316_  (.A(\hash/CA2/_1147_ ),
    .B(\hash/CA2/_1148_ ),
    .COUT(\hash/CA2/_1149_ ),
    .SUM(\hash/CA2/_1150_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2317_  (.A(\hash/CA2/_1151_ ),
    .B(\hash/CA2/_1152_ ),
    .COUT(\hash/CA2/_1153_ ),
    .SUM(\hash/CA2/_1154_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2318_  (.A(\hash/CA2/_1155_ ),
    .B(\hash/CA2/_1156_ ),
    .COUT(\hash/CA2/_1157_ ),
    .SUM(\hash/CA2/_1158_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2319_  (.A(\hash/CA2/_1159_ ),
    .B(\hash/CA2/_1160_ ),
    .COUT(\hash/CA2/_1161_ ),
    .SUM(\hash/CA2/_1162_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2320_  (.A(\hash/CA2/_1163_ ),
    .B(\hash/CA2/_1164_ ),
    .COUT(\hash/CA2/_1165_ ),
    .SUM(\hash/CA2/_1166_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2321_  (.A(\hash/CA2/_1167_ ),
    .B(\hash/CA2/_1168_ ),
    .COUT(\hash/CA2/_1169_ ),
    .SUM(\hash/CA2/_1170_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2322_  (.A(\hash/CA2/_1171_ ),
    .B(\hash/CA2/_1172_ ),
    .COUT(\hash/CA2/_1173_ ),
    .SUM(\hash/CA2/_1174_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2323_  (.A(\hash/CA2/_1175_ ),
    .B(\hash/CA2/_1176_ ),
    .COUT(\hash/CA2/_1177_ ),
    .SUM(\hash/CA2/_1178_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2324_  (.A(\hash/CA2/_1179_ ),
    .B(\hash/CA2/_1180_ ),
    .COUT(\hash/CA2/_1181_ ),
    .SUM(\hash/CA2/_1182_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2325_  (.A(\hash/CA2/_1183_ ),
    .B(\hash/CA2/_1184_ ),
    .COUT(\hash/CA2/_1185_ ),
    .SUM(\hash/CA2/_1186_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2326_  (.A(\hash/CA2/_1187_ ),
    .B(\hash/CA2/_1188_ ),
    .COUT(\hash/CA2/_1189_ ),
    .SUM(\hash/CA2/_1190_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2327_  (.A(\hash/CA2/_1191_ ),
    .B(\hash/CA2/_1192_ ),
    .COUT(\hash/CA2/_1193_ ),
    .SUM(\hash/CA2/_1194_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2328_  (.A(\hash/CA2/_1195_ ),
    .B(\hash/CA2/_1196_ ),
    .COUT(\hash/CA2/_1197_ ),
    .SUM(\hash/CA2/_1198_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2329_  (.A(\hash/CA2/_1199_ ),
    .B(\hash/CA2/_1200_ ),
    .COUT(\hash/CA2/_1201_ ),
    .SUM(\hash/CA2/_1202_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2330_  (.A(\hash/CA2/_1203_ ),
    .B(\hash/CA2/_1204_ ),
    .COUT(\hash/CA2/_1205_ ),
    .SUM(\hash/CA2/_1206_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2331_  (.A(\hash/CA2/_1207_ ),
    .B(\hash/CA2/_0865_ ),
    .COUT(\hash/CA2/_1208_ ),
    .SUM(\hash/CA2/_1209_ ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2332_  (.A(\hash/CA2/_0933_ ),
    .B(\hash/CA2/_1210_ ),
    .COUT(\hash/CA2/_1211_ ),
    .SUM(\hash/a_new[0] ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2333_  (.A(\hash/CA2/_1211_ ),
    .B(\hash/CA2/_1212_ ),
    .COUT(\hash/CA2/_1213_ ),
    .SUM(\hash/a_new[1] ));
 sky130_fd_sc_hd__ha_1 \hash/CA2/_2334_  (.A(\hash/p5_cap[0] ),
    .B(\hash/CA2/_0933_ ),
    .COUT(\hash/CA2/_0869_ ),
    .SUM(\hash/e_new[0] ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1957_  (.A1(\hash/_1720_ ),
    .A2(\hash/_0826_ ),
    .B1(\hash/_1719_ ),
    .Y(\hash/_0827_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_1958_  (.A(\hash/_1724_ ),
    .B(\hash/_0827_ ),
    .Y(\hash/_0144_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_1960_  (.A1(\hash/_1719_ ),
    .A2(\hash/_0822_ ),
    .B1(\hash/_1724_ ),
    .X(\hash/_0829_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_1961_  (.A(\hash/_1723_ ),
    .B(\hash/_0829_ ),
    .Y(\hash/_0830_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_1962_  (.A(\hash/_1726_ ),
    .B(\hash/_0830_ ),
    .Y(\hash/_0145_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_1963_  (.A(\hash/_1724_ ),
    .B(\hash/_1726_ ),
    .Y(\hash/_0831_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1964_  (.A1(\hash/_1726_ ),
    .A2(\hash/_1723_ ),
    .B1(\hash/_1725_ ),
    .Y(\hash/_0832_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_1965_  (.A1(\hash/_0827_ ),
    .A2(\hash/_0831_ ),
    .B1(\hash/_0832_ ),
    .Y(\hash/_0833_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_1966_  (.A(\hash/_1728_ ),
    .B(\hash/_0833_ ),
    .X(\hash/_0146_ ));
 sky130_fd_sc_hd__inv_1 \hash/_1967_  (.A(\hash/_1726_ ),
    .Y(\hash/_0834_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_1968_  (.A1(\hash/_0834_ ),
    .A2(\hash/_0830_ ),
    .B1_N(\hash/_1725_ ),
    .Y(\hash/_0835_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1969_  (.A1(\hash/_1728_ ),
    .A2(\hash/_0835_ ),
    .B1(\hash/_1727_ ),
    .Y(\hash/_0836_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_1970_  (.A(\hash/_1730_ ),
    .B(\hash/_0836_ ),
    .Y(\hash/_0147_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_1971_  (.A1(\hash/_1728_ ),
    .A2(\hash/_0833_ ),
    .B1(\hash/_1727_ ),
    .X(\hash/_0837_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1972_  (.A1(\hash/_1730_ ),
    .A2(\hash/_0837_ ),
    .B1(\hash/_1729_ ),
    .Y(\hash/_0838_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_1973_  (.A(\hash/_1732_ ),
    .B(\hash/_0838_ ),
    .Y(\hash/_0148_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1974_  (.A1(\hash/_1728_ ),
    .A2(\hash/_1725_ ),
    .B1(\hash/_1727_ ),
    .Y(\hash/_0839_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_1975_  (.A(\hash/_1730_ ),
    .B(\hash/_1732_ ),
    .Y(\hash/_0840_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1976_  (.A1(\hash/_1732_ ),
    .A2(\hash/_1729_ ),
    .B1(\hash/_1731_ ),
    .Y(\hash/_0841_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_1977_  (.A1(\hash/_0839_ ),
    .A2(\hash/_0840_ ),
    .B1(\hash/_0841_ ),
    .Y(\hash/_0842_ ));
 sky130_fd_sc_hd__and3_1 \hash/_1978_  (.A(\hash/_1728_ ),
    .B(\hash/_1730_ ),
    .C(\hash/_1732_ ),
    .X(\hash/_0843_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_1979_  (.A(\hash/_1726_ ),
    .B(\hash/_1723_ ),
    .Y(\hash/_0844_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_1980_  (.A(\hash/_1724_ ),
    .B(\hash/_1726_ ),
    .C(\hash/_1719_ ),
    .Y(\hash/_0845_ ));
 sky130_fd_sc_hd__a21boi_1 \hash/_1981_  (.A1(\hash/_0844_ ),
    .A2(\hash/_0845_ ),
    .B1_N(\hash/_0843_ ),
    .Y(\hash/_0846_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_1982_  (.A1(\hash/_1724_ ),
    .A2(\hash/_1726_ ),
    .A3(\hash/_0822_ ),
    .A4(\hash/_0843_ ),
    .B1(\hash/_0846_ ),
    .Y(\hash/_0847_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_1983_  (.A(\hash/_0842_ ),
    .B_N(\hash/_0847_ ),
    .Y(\hash/_0848_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_1984_  (.A(\hash/_1734_ ),
    .B(\hash/_0848_ ),
    .Y(\hash/_0149_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_1985_  (.A1(\hash/_1730_ ),
    .A2(\hash/_1727_ ),
    .B1(\hash/_1729_ ),
    .X(\hash/_0849_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1986_  (.A1(\hash/_1732_ ),
    .A2(\hash/_0849_ ),
    .B1(\hash/_1731_ ),
    .Y(\hash/_0850_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_1987_  (.A(\hash/_0833_ ),
    .B(\hash/_0843_ ),
    .Y(\hash/_0851_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_1988_  (.A(\hash/_0850_ ),
    .B(\hash/_0851_ ),
    .Y(\hash/_0852_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1989_  (.A1(\hash/_1734_ ),
    .A2(\hash/_0852_ ),
    .B1(\hash/_1733_ ),
    .Y(\hash/_0853_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_1990_  (.A(\hash/_1736_ ),
    .B(\hash/_0853_ ),
    .Y(\hash/_0120_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_1991_  (.A(\hash/_1733_ ),
    .B(\hash/_1735_ ),
    .C(\hash/_0842_ ),
    .Y(\hash/_0854_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_1992_  (.A1(\hash/_1734_ ),
    .A2(\hash/_1733_ ),
    .B1(\hash/_1736_ ),
    .X(\hash/_0855_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \hash/_1993_  (.A1_N(\hash/_0847_ ),
    .A2_N(\hash/_0854_ ),
    .B1(\hash/_0855_ ),
    .B2(\hash/_1735_ ),
    .Y(\hash/_0856_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_1994_  (.A(\hash/_1738_ ),
    .B(\hash/_0856_ ),
    .Y(\hash/_0121_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_1995_  (.A(\hash/_1734_ ),
    .B(\hash/_1736_ ),
    .Y(\hash/_0857_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_1996_  (.A1(\hash/_1736_ ),
    .A2(\hash/_1733_ ),
    .B1(\hash/_1735_ ),
    .Y(\hash/_0858_ ));
 sky130_fd_sc_hd__inv_1 \hash/_1997_  (.A(\hash/_1737_ ),
    .Y(\hash/_0859_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_1998_  (.A1(\hash/_0850_ ),
    .A2(\hash/_0857_ ),
    .B1(\hash/_0858_ ),
    .C1(\hash/_0859_ ),
    .Y(\hash/_0860_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_1999_  (.A1(\hash/_1734_ ),
    .A2(\hash/_1736_ ),
    .A3(\hash/_0833_ ),
    .A4(\hash/_0843_ ),
    .B1(\hash/_0860_ ),
    .Y(\hash/_0861_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2000_  (.A(\hash/_1738_ ),
    .B(\hash/_1737_ ),
    .Y(\hash/_0862_ ));
 sky130_fd_sc_hd__or2_2 \hash/_2001_  (.A(\hash/_0861_ ),
    .B(\hash/_0862_ ),
    .X(\hash/_0863_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2002_  (.A(\hash/_1740_ ),
    .B(\hash/_0863_ ),
    .Y(\hash/_0122_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2003_  (.A(\hash/_1738_ ),
    .Y(\hash/_0864_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2004_  (.A1(\hash/_0864_ ),
    .A2(\hash/_0856_ ),
    .B1(\hash/_0859_ ),
    .Y(\hash/_0865_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2005_  (.A1(\hash/_1740_ ),
    .A2(\hash/_0865_ ),
    .B1(\hash/_1739_ ),
    .Y(\hash/_0866_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2006_  (.A(\hash/_1742_ ),
    .B(\hash/_0866_ ),
    .Y(\hash/_0123_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2007_  (.A(\hash/_1744_ ),
    .Y(\hash/_0867_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2008_  (.A(\hash/_1740_ ),
    .B(\hash/_1742_ ),
    .Y(\hash/_0868_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2009_  (.A1(\hash/_1742_ ),
    .A2(\hash/_1739_ ),
    .B1(\hash/_1741_ ),
    .Y(\hash/_0869_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2010_  (.A1(\hash/_0863_ ),
    .A2(\hash/_0868_ ),
    .B1(\hash/_0869_ ),
    .Y(\hash/_0870_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2011_  (.A(\hash/_0867_ ),
    .B(\hash/_0870_ ),
    .Y(\hash/_0124_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2012_  (.A(\hash/_1738_ ),
    .B(\hash/_1740_ ),
    .C(\hash/_1742_ ),
    .Y(\hash/_0871_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2013_  (.A1(\hash/_1740_ ),
    .A2(\hash/_1737_ ),
    .B1(\hash/_1739_ ),
    .X(\hash/_0872_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2014_  (.A1(\hash/_1742_ ),
    .A2(\hash/_0872_ ),
    .B1(\hash/_1741_ ),
    .Y(\hash/_0873_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2015_  (.A1(\hash/_0856_ ),
    .A2(\hash/_0871_ ),
    .B1(\hash/_0873_ ),
    .Y(\hash/_0874_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2016_  (.A1(\hash/_1744_ ),
    .A2(\hash/_0874_ ),
    .B1(\hash/_1743_ ),
    .X(\hash/_0875_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2017_  (.A(\hash/_1748_ ),
    .B(\hash/_0875_ ),
    .X(\hash/_0125_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2019_  (.A(\hash/_1740_ ),
    .B(\hash/_1742_ ),
    .C(\hash/_1744_ ),
    .D(\hash/_1748_ ),
    .Y(\hash/_0877_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2020_  (.A1(\hash/_0867_ ),
    .A2(\hash/_0869_ ),
    .B1_N(\hash/_1743_ ),
    .Y(\hash/_0878_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2021_  (.A1(\hash/_1748_ ),
    .A2(\hash/_0878_ ),
    .B1(\hash/_1747_ ),
    .Y(\hash/_0879_ ));
 sky130_fd_sc_hd__o31a_1 \hash/_2022_  (.A1(\hash/_0861_ ),
    .A2(\hash/_0862_ ),
    .A3(\hash/_0877_ ),
    .B1(\hash/_0879_ ),
    .X(\hash/_0880_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2023_  (.A(\hash/_1746_ ),
    .B(\hash/_0880_ ),
    .Y(\hash/_0126_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2024_  (.A1(\hash/_0858_ ),
    .A2(\hash/_0871_ ),
    .B1(\hash/_0873_ ),
    .Y(\hash/_0881_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2025_  (.A1(\hash/_1744_ ),
    .A2(\hash/_0881_ ),
    .B1(\hash/_1743_ ),
    .X(\hash/_0882_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2026_  (.A1(\hash/_1748_ ),
    .A2(\hash/_0882_ ),
    .B1(\hash/_1747_ ),
    .X(\hash/_0883_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2027_  (.A(\hash/_1738_ ),
    .B(\hash/_1746_ ),
    .Y(\hash/_0884_ ));
 sky130_fd_sc_hd__nor4_1 \hash/_2028_  (.A(\hash/_0848_ ),
    .B(\hash/_0857_ ),
    .C(\hash/_0877_ ),
    .D(\hash/_0884_ ),
    .Y(\hash/_0885_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_2029_  (.A1(\hash/_1746_ ),
    .A2(\hash/_0883_ ),
    .B1(\hash/_0885_ ),
    .C1(\hash/_1745_ ),
    .Y(\hash/_0886_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2030_  (.A(\hash/_1750_ ),
    .B(\hash/_0886_ ),
    .Y(\hash/_0127_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2031_  (.A(\hash/_1752_ ),
    .Y(\hash/_0887_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2032_  (.A(\hash/_1746_ ),
    .B(\hash/_1750_ ),
    .Y(\hash/_0888_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2033_  (.A1(\hash/_1750_ ),
    .A2(\hash/_1745_ ),
    .B1(\hash/_1749_ ),
    .Y(\hash/_0889_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2034_  (.A1(\hash/_0880_ ),
    .A2(\hash/_0888_ ),
    .B1(\hash/_0889_ ),
    .Y(\hash/_0890_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2035_  (.A(\hash/_0887_ ),
    .B(\hash/_0890_ ),
    .Y(\hash/_0128_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2036_  (.A1(\hash/_1746_ ),
    .A2(\hash/_1747_ ),
    .B1(\hash/_1745_ ),
    .X(\hash/_0891_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2037_  (.A1(\hash/_1750_ ),
    .A2(\hash/_0891_ ),
    .B1(\hash/_1749_ ),
    .X(\hash/_0892_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2038_  (.A1(\hash/_1752_ ),
    .A2(\hash/_0892_ ),
    .B1(\hash/_1751_ ),
    .Y(\hash/_0893_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2039_  (.A(\hash/_1743_ ),
    .B_N(\hash/_0893_ ),
    .Y(\hash/_0894_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2040_  (.A(\hash/_1748_ ),
    .B(\hash/_1746_ ),
    .C(\hash/_1750_ ),
    .X(\hash/_0895_ ));
 sky130_fd_sc_hd__nand3b_1 \hash/_2041_  (.A_N(\hash/_1743_ ),
    .B(\hash/_0873_ ),
    .C(\hash/_0871_ ),
    .Y(\hash/_0896_ ));
 sky130_fd_sc_hd__o2111ai_1 \hash/_2042_  (.A1(\hash/_1744_ ),
    .A2(\hash/_1743_ ),
    .B1(\hash/_0895_ ),
    .C1(\hash/_0896_ ),
    .D1(\hash/_1752_ ),
    .Y(\hash/_0897_ ));
 sky130_fd_sc_hd__a32oi_1 \hash/_2043_  (.A1(\hash/_0856_ ),
    .A2(\hash/_0873_ ),
    .A3(\hash/_0894_ ),
    .B1(\hash/_0897_ ),
    .B2(\hash/_0893_ ),
    .Y(\hash/_0898_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2044_  (.A(\hash/_1754_ ),
    .B(\hash/_0898_ ),
    .X(\hash/_0129_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2046_  (.A(\hash/_1746_ ),
    .B(\hash/_1750_ ),
    .C(\hash/_1752_ ),
    .D(\hash/_1754_ ),
    .Y(\hash/_0900_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2047_  (.A1(\hash/_0887_ ),
    .A2(\hash/_0889_ ),
    .B1_N(\hash/_1751_ ),
    .Y(\hash/_0901_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2048_  (.A1(\hash/_1754_ ),
    .A2(\hash/_0901_ ),
    .B1(\hash/_1753_ ),
    .Y(\hash/_0902_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2049_  (.A1(\hash/_0880_ ),
    .A2(\hash/_0900_ ),
    .B1(\hash/_0902_ ),
    .Y(\hash/_0903_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2050_  (.A(\hash/_1756_ ),
    .B(\hash/_0903_ ),
    .X(\hash/_0130_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2051_  (.A1(\hash/_1754_ ),
    .A2(\hash/_0898_ ),
    .B1(\hash/_1753_ ),
    .X(\hash/_0904_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2052_  (.A1(\hash/_1756_ ),
    .A2(\hash/_0904_ ),
    .B1(\hash/_1755_ ),
    .Y(\hash/_0905_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2053_  (.A(\hash/_1758_ ),
    .B(\hash/_0905_ ),
    .Y(\hash/_0131_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2054_  (.A1(\hash/_1758_ ),
    .A2(\hash/_1755_ ),
    .B1(\hash/_1757_ ),
    .Y(\hash/_0906_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2055_  (.A(\hash/_1756_ ),
    .B(\hash/_1758_ ),
    .C(\hash/_0903_ ),
    .Y(\hash/_0907_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2056_  (.A(\hash/_0906_ ),
    .B(\hash/_0907_ ),
    .Y(\hash/_0908_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2057_  (.A(\hash/_1760_ ),
    .B(\hash/_0908_ ),
    .X(\hash/_0132_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2058_  (.A(\hash/_1758_ ),
    .B(\hash/_1760_ ),
    .Y(\hash/_0909_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2059_  (.A(\hash/_1754_ ),
    .B(\hash/_1756_ ),
    .Y(\hash/_0910_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2060_  (.A(\hash/_0909_ ),
    .B(\hash/_0910_ ),
    .Y(\hash/_0911_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2061_  (.A1(\hash/_1756_ ),
    .A2(\hash/_1753_ ),
    .B1(\hash/_1755_ ),
    .Y(\hash/_0912_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2062_  (.A1(\hash/_1760_ ),
    .A2(\hash/_1757_ ),
    .B1(\hash/_1759_ ),
    .Y(\hash/_0913_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2063_  (.A1(\hash/_0909_ ),
    .A2(\hash/_0912_ ),
    .B1(\hash/_0913_ ),
    .Y(\hash/_0914_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2064_  (.A1(\hash/_0898_ ),
    .A2(\hash/_0911_ ),
    .B1(\hash/_0914_ ),
    .Y(\hash/_0915_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2065_  (.A(\hash/_1762_ ),
    .B(\hash/_0915_ ),
    .Y(\hash/_0133_ ));
 sky130_fd_sc_hd__and2_1 \hash/_2067_  (.A(\hash/_1760_ ),
    .B(\hash/_1762_ ),
    .X(\hash/_0917_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2068_  (.A(\hash/_1756_ ),
    .B(\hash/_1758_ ),
    .C(\hash/_0903_ ),
    .D(\hash/_0917_ ),
    .Y(\hash/_0918_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2069_  (.A1(\hash/_1762_ ),
    .A2(\hash/_1759_ ),
    .B1(\hash/_1761_ ),
    .X(\hash/_0919_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2070_  (.A(\hash/_0906_ ),
    .B_N(\hash/_0917_ ),
    .Y(\hash/_0920_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2071_  (.A(\hash/_0919_ ),
    .B(\hash/_0920_ ),
    .Y(\hash/_0921_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2072_  (.A(\hash/_0918_ ),
    .B(\hash/_0921_ ),
    .Y(\hash/_0922_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2073_  (.A(\hash/_1764_ ),
    .B(\hash/_0922_ ),
    .X(\hash/_0134_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2074_  (.A(\hash/_1766_ ),
    .Y(\hash/_0923_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2075_  (.A(\hash/_1762_ ),
    .B(\hash/_1764_ ),
    .Y(\hash/_0924_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2076_  (.A1(\hash/_1764_ ),
    .A2(\hash/_1761_ ),
    .B1(\hash/_1763_ ),
    .Y(\hash/_0925_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2077_  (.A1(\hash/_0915_ ),
    .A2(\hash/_0924_ ),
    .B1(\hash/_0925_ ),
    .Y(\hash/_0926_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2078_  (.A(\hash/_0923_ ),
    .B(\hash/_0926_ ),
    .Y(\hash/_0135_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2079_  (.A(\hash/_1768_ ),
    .Y(\hash/_0927_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_2080_  (.A1(\hash/_1756_ ),
    .A2(\hash/_1758_ ),
    .A3(\hash/_0903_ ),
    .A4(\hash/_0917_ ),
    .B1(\hash/_0920_ ),
    .Y(\hash/_0928_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2081_  (.A(\hash/_1764_ ),
    .B(\hash/_1766_ ),
    .Y(\hash/_0929_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2082_  (.A1(\hash/_1764_ ),
    .A2(\hash/_0919_ ),
    .B1(\hash/_1763_ ),
    .Y(\hash/_0930_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2083_  (.A(\hash/_0923_ ),
    .B(\hash/_0930_ ),
    .Y(\hash/_0931_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2084_  (.A(\hash/_1765_ ),
    .B(\hash/_0931_ ),
    .Y(\hash/_0932_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2085_  (.A1(\hash/_0928_ ),
    .A2(\hash/_0929_ ),
    .B1(\hash/_0932_ ),
    .Y(\hash/_0933_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2086_  (.A(\hash/_0927_ ),
    .B(\hash/_0933_ ),
    .Y(\hash/_0136_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2087_  (.A(\hash/_1762_ ),
    .B(\hash/_1764_ ),
    .C(\hash/_1766_ ),
    .D(\hash/_1768_ ),
    .Y(\hash/_0934_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2088_  (.A1(\hash/_0923_ ),
    .A2(\hash/_0925_ ),
    .B1_N(\hash/_1765_ ),
    .Y(\hash/_0935_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2089_  (.A1(\hash/_1768_ ),
    .A2(\hash/_0935_ ),
    .B1(\hash/_1767_ ),
    .Y(\hash/_0936_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2090_  (.A1(\hash/_0915_ ),
    .A2(\hash/_0934_ ),
    .B1(\hash/_0936_ ),
    .Y(\hash/_0937_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2091_  (.A(\hash/_1770_ ),
    .B(\hash/_0937_ ),
    .X(\hash/_0137_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2092_  (.A(\hash/_1764_ ),
    .B(\hash/_1766_ ),
    .C(\hash/_1768_ ),
    .D(\hash/_1770_ ),
    .Y(\hash/_0938_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2093_  (.A1(\hash/_1766_ ),
    .A2(\hash/_1763_ ),
    .B1(\hash/_1765_ ),
    .Y(\hash/_0939_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2094_  (.A(\hash/_1767_ ),
    .Y(\hash/_0940_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2095_  (.A1(\hash/_0927_ ),
    .A2(\hash/_0939_ ),
    .B1(\hash/_0940_ ),
    .Y(\hash/_0941_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2096_  (.A(\hash/_0921_ ),
    .B(\hash/_0938_ ),
    .Y(\hash/_0942_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_2097_  (.A1(\hash/_1770_ ),
    .A2(\hash/_0941_ ),
    .B1(\hash/_0942_ ),
    .C1(\hash/_1769_ ),
    .Y(\hash/_0943_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2098_  (.A1(\hash/_0918_ ),
    .A2(\hash/_0938_ ),
    .B1(\hash/_0943_ ),
    .Y(\hash/_0944_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2099_  (.A(\hash/_1772_ ),
    .B(\hash/_0944_ ),
    .X(\hash/_0138_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2100_  (.A(\hash/_1770_ ),
    .B(\hash/_1772_ ),
    .Y(\hash/_0945_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2101_  (.A1(\hash/_0913_ ),
    .A2(\hash/_0924_ ),
    .B1(\hash/_0925_ ),
    .Y(\hash/_0946_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2102_  (.A1(\hash/_1766_ ),
    .A2(\hash/_0946_ ),
    .B1(\hash/_1765_ ),
    .Y(\hash/_0947_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2103_  (.A(\hash/_0927_ ),
    .B(\hash/_0947_ ),
    .Y(\hash/_0948_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2104_  (.A(\hash/_1767_ ),
    .B(\hash/_0948_ ),
    .Y(\hash/_0949_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2105_  (.A1(\hash/_1772_ ),
    .A2(\hash/_1769_ ),
    .B1(\hash/_1771_ ),
    .Y(\hash/_0950_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2106_  (.A1(\hash/_0949_ ),
    .A2(\hash/_0945_ ),
    .B1(\hash/_0950_ ),
    .X(\hash/_0951_ ));
 sky130_fd_sc_hd__o41ai_1 \hash/_2107_  (.A1(\hash/_0905_ ),
    .A2(\hash/_0909_ ),
    .A3(\hash/_0934_ ),
    .A4(\hash/_0945_ ),
    .B1(\hash/_0951_ ),
    .Y(\hash/_0952_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2108_  (.A(\hash/_1774_ ),
    .B(\hash/_0952_ ),
    .X(\hash/_0139_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2109_  (.A(\hash/_1770_ ),
    .B(\hash/_1772_ ),
    .C(\hash/_1774_ ),
    .X(\hash/_0953_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2110_  (.A(\hash/_1764_ ),
    .B(\hash/_1766_ ),
    .C(\hash/_1768_ ),
    .D(\hash/_0953_ ),
    .Y(\hash/_0954_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2111_  (.A1(\hash/_0927_ ),
    .A2(\hash/_0932_ ),
    .B1(\hash/_0950_ ),
    .C1(\hash/_0940_ ),
    .Y(\hash/_0955_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2112_  (.A1(\hash/_1770_ ),
    .A2(\hash/_1769_ ),
    .B1(\hash/_1772_ ),
    .Y(\hash/_0956_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2113_  (.A_N(\hash/_1771_ ),
    .B(\hash/_0956_ ),
    .Y(\hash/_0957_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2114_  (.A1(\hash/_1774_ ),
    .A2(\hash/_0955_ ),
    .A3(\hash/_0957_ ),
    .B1(\hash/_1773_ ),
    .Y(\hash/_0958_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2115_  (.A1(\hash/_0928_ ),
    .A2(\hash/_0954_ ),
    .B1(\hash/_0958_ ),
    .Y(\hash/_0959_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2116_  (.A(\hash/_1776_ ),
    .B(\hash/_0959_ ),
    .X(\hash/_0141_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_2117_  (.A0(\hash/e_new[31] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[31] ));
 sky130_fd_sc_hd__nor2_1 \hash/_2118_  (.A(\hash/_0915_ ),
    .B(\hash/_0934_ ),
    .Y(\hash/_0960_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2119_  (.A1(\hash/_0936_ ),
    .A2(\hash/_0945_ ),
    .B1(\hash/_0950_ ),
    .Y(\hash/_0961_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2120_  (.A1(\hash/_1774_ ),
    .A2(\hash/_0961_ ),
    .B1(\hash/_1773_ ),
    .Y(\hash/_0962_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2121_  (.A(\hash/_0962_ ),
    .B_N(\hash/_1776_ ),
    .Y(\hash/_0963_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/_2122_  (.A1(\hash/_1776_ ),
    .A2(\hash/_0960_ ),
    .A3(\hash/_0953_ ),
    .B1(\hash/_0963_ ),
    .C1(\hash/_1775_ ),
    .Y(\hash/_0964_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2123_  (.A(_09578_),
    .B(\hash/e_new[31] ),
    .Y(\hash/_0965_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2124_  (.A(reset_hash_dash),
    .B(\hash/_0965_ ),
    .Y(\hash/_0966_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2125_  (.A(\hash/_0964_ ),
    .B(\hash/_0966_ ),
    .Y(\hash/_0142_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2126_  (.A(\hash/_1472_ ),
    .B(\hash/_1782_ ),
    .X(\hash/_0170_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2127_  (.A1(\hash/_1471_ ),
    .A2(\hash/_1778_ ),
    .B1(\hash/_1777_ ),
    .X(\hash/_0967_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2128_  (.A1(\hash/_1782_ ),
    .A2(\hash/_0967_ ),
    .B1(\hash/_1781_ ),
    .Y(\hash/_0968_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2129_  (.A(\hash/_1780_ ),
    .B(\hash/_0968_ ),
    .Y(\hash/_0173_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2130_  (.A1(\hash/_1472_ ),
    .A2(\hash/_1782_ ),
    .B1(\hash/_1781_ ),
    .X(\hash/_0969_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2131_  (.A1(\hash/_1780_ ),
    .A2(\hash/_0969_ ),
    .B1(\hash/_1779_ ),
    .Y(\hash/_0970_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2132_  (.A(\hash/_1784_ ),
    .B(\hash/_0970_ ),
    .Y(\hash/_0174_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2133_  (.A(\hash/_1784_ ),
    .Y(\hash/_0971_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2134_  (.A(\hash/_0968_ ),
    .B_N(\hash/_1780_ ),
    .Y(\hash/_0972_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2135_  (.A(\hash/_1779_ ),
    .B(\hash/_0972_ ),
    .Y(\hash/_0973_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2136_  (.A(\hash/_0971_ ),
    .B(\hash/_0973_ ),
    .Y(\hash/_0974_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2137_  (.A(\hash/_1783_ ),
    .B(\hash/_0974_ ),
    .Y(\hash/_0975_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2138_  (.A(\hash/_1786_ ),
    .B(\hash/_0975_ ),
    .Y(\hash/_0175_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2139_  (.A1(\hash/_0971_ ),
    .A2(\hash/_0970_ ),
    .B1_N(\hash/_1783_ ),
    .Y(\hash/_0976_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2140_  (.A1(\hash/_1786_ ),
    .A2(\hash/_0976_ ),
    .B1(\hash/_1785_ ),
    .Y(\hash/_0977_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2141_  (.A(\hash/_1788_ ),
    .B(\hash/_0977_ ),
    .Y(\hash/_0176_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2142_  (.A(\hash/_1786_ ),
    .Y(\hash/_0978_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2143_  (.A1(\hash/_0978_ ),
    .A2(\hash/_0975_ ),
    .B1_N(\hash/_1785_ ),
    .Y(\hash/_0979_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2144_  (.A1(\hash/_1788_ ),
    .A2(\hash/_0979_ ),
    .B1(\hash/_1787_ ),
    .Y(\hash/_0980_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2145_  (.A(\hash/_1790_ ),
    .B(\hash/_0980_ ),
    .Y(\hash/_0177_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2146_  (.A(\hash/_1788_ ),
    .Y(\hash/_0981_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2147_  (.A1(\hash/_0981_ ),
    .A2(\hash/_0977_ ),
    .B1_N(\hash/_1787_ ),
    .Y(\hash/_0982_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2148_  (.A1(\hash/_1790_ ),
    .A2(\hash/_0982_ ),
    .B1(\hash/_1789_ ),
    .Y(\hash/_0983_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2149_  (.A(\hash/_1792_ ),
    .B(\hash/_0983_ ),
    .Y(\hash/_0178_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2150_  (.A(\hash/_1788_ ),
    .B(\hash/_1790_ ),
    .C(\hash/_1792_ ),
    .Y(\hash/_0984_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2151_  (.A(\hash/_0971_ ),
    .B(\hash/_0978_ ),
    .C(\hash/_0984_ ),
    .Y(\hash/_0985_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2152_  (.A(\hash/_1786_ ),
    .B(\hash/_1783_ ),
    .Y(\hash/_0986_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2153_  (.A(\hash/_1784_ ),
    .B(\hash/_1786_ ),
    .C(\hash/_1779_ ),
    .Y(\hash/_0987_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2154_  (.A1(\hash/_0986_ ),
    .A2(\hash/_0987_ ),
    .B1(\hash/_0984_ ),
    .Y(\hash/_0988_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2155_  (.A1(\hash/_0972_ ),
    .A2(\hash/_0985_ ),
    .B1(\hash/_0988_ ),
    .Y(\hash/_0989_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2156_  (.A1(\hash/_1788_ ),
    .A2(\hash/_1785_ ),
    .B1(\hash/_1787_ ),
    .X(\hash/_0990_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2157_  (.A1(\hash/_1790_ ),
    .A2(\hash/_0990_ ),
    .B1(\hash/_1789_ ),
    .X(\hash/_0991_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2158_  (.A1(\hash/_1792_ ),
    .A2(\hash/_0991_ ),
    .B1(\hash/_1791_ ),
    .Y(\hash/_0992_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2159_  (.A(\hash/_0989_ ),
    .B(\hash/_0992_ ),
    .Y(\hash/_0993_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2160_  (.A(\hash/_1794_ ),
    .B(\hash/_0993_ ),
    .X(\hash/_0179_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2161_  (.A(\hash/_1792_ ),
    .Y(\hash/_0994_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2162_  (.A1(\hash/_0994_ ),
    .A2(\hash/_0983_ ),
    .B1_N(\hash/_1791_ ),
    .Y(\hash/_0995_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2163_  (.A1(\hash/_1794_ ),
    .A2(\hash/_0995_ ),
    .B1(\hash/_1793_ ),
    .Y(\hash/_0996_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2164_  (.A(\hash/_1796_ ),
    .B(\hash/_0996_ ),
    .Y(\hash/_0150_ ));
 sky130_fd_sc_hd__nor3b_1 \hash/_2165_  (.A(\hash/_1793_ ),
    .B(\hash/_1795_ ),
    .C_N(\hash/_0992_ ),
    .Y(\hash/_0997_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2166_  (.A1(\hash/_1794_ ),
    .A2(\hash/_1793_ ),
    .B1(\hash/_1796_ ),
    .X(\hash/_0998_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2167_  (.A(\hash/_1795_ ),
    .B(\hash/_0998_ ),
    .Y(\hash/_0999_ ));
 sky130_fd_sc_hd__a21oi_2 \hash/_2168_  (.A1(\hash/_0989_ ),
    .A2(\hash/_0997_ ),
    .B1(\hash/_0999_ ),
    .Y(\hash/_1000_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2169_  (.A(\hash/_1798_ ),
    .B(\hash/_1000_ ),
    .X(\hash/_0151_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2171_  (.A(\hash/_1783_ ),
    .B(\hash/_1785_ ),
    .Y(\hash/_1002_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2172_  (.A1(\hash/_0971_ ),
    .A2(\hash/_0970_ ),
    .B1(\hash/_1002_ ),
    .Y(\hash/_1003_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2173_  (.A(\hash/_1794_ ),
    .B(\hash/_1796_ ),
    .Y(\hash/_1004_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2174_  (.A(\hash/_1786_ ),
    .B(\hash/_1785_ ),
    .Y(\hash/_1005_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2175_  (.A(\hash/_0984_ ),
    .B(\hash/_1004_ ),
    .C(\hash/_1005_ ),
    .Y(\hash/_1006_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2176_  (.A1(\hash/_1790_ ),
    .A2(\hash/_1787_ ),
    .B1(\hash/_1789_ ),
    .X(\hash/_1007_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2177_  (.A1(\hash/_1792_ ),
    .A2(\hash/_1007_ ),
    .B1(\hash/_1791_ ),
    .Y(\hash/_1008_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2178_  (.A(\hash/_1796_ ),
    .B(\hash/_1793_ ),
    .Y(\hash/_1009_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2179_  (.A1(\hash/_1004_ ),
    .A2(\hash/_1008_ ),
    .B1(\hash/_1009_ ),
    .Y(\hash/_1010_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_2180_  (.A1(\hash/_1003_ ),
    .A2(\hash/_1006_ ),
    .B1(\hash/_1010_ ),
    .C1(\hash/_1795_ ),
    .Y(\hash/_1011_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2181_  (.A(\hash/_1011_ ),
    .Y(\hash/_1012_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2182_  (.A1(\hash/_1798_ ),
    .A2(\hash/_1012_ ),
    .B1(\hash/_1797_ ),
    .Y(\hash/_1013_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2183_  (.A(\hash/_1800_ ),
    .B(\hash/_1013_ ),
    .Y(\hash/_0152_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2185_  (.A1(\hash/_1798_ ),
    .A2(\hash/_1000_ ),
    .B1(\hash/_1797_ ),
    .X(\hash/_1015_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2186_  (.A1(\hash/_1800_ ),
    .A2(\hash/_1015_ ),
    .B1(\hash/_1799_ ),
    .Y(\hash/_1016_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2187_  (.A(\hash/_1802_ ),
    .B(\hash/_1016_ ),
    .Y(\hash/_0153_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2188_  (.A(\hash/_1798_ ),
    .B(\hash/_1800_ ),
    .C(\hash/_1802_ ),
    .Y(\hash/_1017_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2189_  (.A1(\hash/_1802_ ),
    .A2(\hash/_1799_ ),
    .B1(\hash/_1801_ ),
    .X(\hash/_1018_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2190_  (.A1(\hash/_1800_ ),
    .A2(\hash/_1802_ ),
    .A3(\hash/_1797_ ),
    .B1(\hash/_1018_ ),
    .Y(\hash/_1019_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2191_  (.A1(\hash/_1011_ ),
    .A2(\hash/_1017_ ),
    .B1(\hash/_1019_ ),
    .Y(\hash/_1020_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2192_  (.A(\hash/_1804_ ),
    .B(\hash/_1020_ ),
    .X(\hash/_0154_ ));
 sky130_fd_sc_hd__a31o_2 \hash/_2193_  (.A1(\hash/_1800_ ),
    .A2(\hash/_1802_ ),
    .A3(\hash/_1797_ ),
    .B1(\hash/_1018_ ),
    .X(\hash/_1021_ ));
 sky130_fd_sc_hd__a41o_1 \hash/_2194_  (.A1(\hash/_1798_ ),
    .A2(\hash/_1800_ ),
    .A3(\hash/_1802_ ),
    .A4(\hash/_1000_ ),
    .B1(\hash/_1021_ ),
    .X(\hash/_1022_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2195_  (.A1(\hash/_1804_ ),
    .A2(\hash/_1022_ ),
    .B1(\hash/_1803_ ),
    .Y(\hash/_1023_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2196_  (.A(\hash/_1808_ ),
    .B(\hash/_1023_ ),
    .Y(\hash/_0155_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2197_  (.A(\hash/_1804_ ),
    .B(\hash/_1808_ ),
    .Y(\hash/_1024_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2198_  (.A(\hash/_1024_ ),
    .Y(\hash/_1025_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2199_  (.A(\hash/_1800_ ),
    .B(\hash/_1802_ ),
    .C(\hash/_1025_ ),
    .Y(\hash/_1026_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2200_  (.A(\hash/_1803_ ),
    .Y(\hash/_1027_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2201_  (.A(\hash/_1804_ ),
    .B(\hash/_1018_ ),
    .Y(\hash/_1028_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2202_  (.A(\hash/_1027_ ),
    .B(\hash/_1028_ ),
    .Y(\hash/_1029_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2203_  (.A1(\hash/_1808_ ),
    .A2(\hash/_1029_ ),
    .B1(\hash/_1807_ ),
    .Y(\hash/_1030_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2204_  (.A1(\hash/_1013_ ),
    .A2(\hash/_1026_ ),
    .B1(\hash/_1030_ ),
    .Y(\hash/_1031_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2205_  (.A(\hash/_1806_ ),
    .B(\hash/_1031_ ),
    .X(\hash/_0156_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2206_  (.A(\hash/_1004_ ),
    .B(\hash/_1017_ ),
    .C(\hash/_1024_ ),
    .Y(\hash/_1032_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2207_  (.A1(\hash/_1796_ ),
    .A2(\hash/_1793_ ),
    .B1(\hash/_1795_ ),
    .Y(\hash/_1033_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2208_  (.A(\hash/_1017_ ),
    .B(\hash/_1033_ ),
    .Y(\hash/_1034_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2209_  (.A1(\hash/_1021_ ),
    .A2(\hash/_1034_ ),
    .B1(\hash/_1804_ ),
    .Y(\hash/_1035_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2210_  (.A(\hash/_1027_ ),
    .B(\hash/_1035_ ),
    .Y(\hash/_1036_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2211_  (.A1(\hash/_1808_ ),
    .A2(\hash/_1036_ ),
    .B1(\hash/_1807_ ),
    .Y(\hash/_1037_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2212_  (.A(\hash/_1037_ ),
    .B_N(\hash/_1806_ ),
    .Y(\hash/_1038_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/_2213_  (.A1(\hash/_1806_ ),
    .A2(\hash/_0993_ ),
    .A3(\hash/_1032_ ),
    .B1(\hash/_1038_ ),
    .C1(\hash/_1805_ ),
    .Y(\hash/_1039_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2214_  (.A(\hash/_1810_ ),
    .B(\hash/_1039_ ),
    .Y(\hash/_0157_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2215_  (.A1(\hash/_1808_ ),
    .A2(\hash/_1803_ ),
    .B1(\hash/_1807_ ),
    .X(\hash/_1040_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2216_  (.A1(\hash/_1806_ ),
    .A2(\hash/_1040_ ),
    .B1(\hash/_1805_ ),
    .X(\hash/_1041_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2217_  (.A1(\hash/_1810_ ),
    .A2(\hash/_1041_ ),
    .B1(\hash/_1809_ ),
    .Y(\hash/_1042_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2218_  (.A(\hash/_1806_ ),
    .B(\hash/_1810_ ),
    .C(\hash/_1020_ ),
    .D(\hash/_1025_ ),
    .Y(\hash/_1043_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2219_  (.A(\hash/_1042_ ),
    .B(\hash/_1043_ ),
    .Y(\hash/_1044_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2220_  (.A(\hash/_1812_ ),
    .B(\hash/_1044_ ),
    .X(\hash/_0158_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2221_  (.A1(\hash/_1806_ ),
    .A2(\hash/_1807_ ),
    .B1(\hash/_1805_ ),
    .X(\hash/_1045_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2222_  (.A1(\hash/_1810_ ),
    .A2(\hash/_1045_ ),
    .B1(\hash/_1809_ ),
    .X(\hash/_1046_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2223_  (.A1(\hash/_1812_ ),
    .A2(\hash/_1046_ ),
    .B1(\hash/_1811_ ),
    .X(\hash/_1047_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2224_  (.A(\hash/_1806_ ),
    .B(\hash/_1810_ ),
    .C(\hash/_1812_ ),
    .X(\hash/_1048_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2225_  (.A1(\hash/_1804_ ),
    .A2(\hash/_1803_ ),
    .B1(\hash/_1048_ ),
    .C1(\hash/_1808_ ),
    .Y(\hash/_1049_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2226_  (.A1(\hash/_1027_ ),
    .A2(\hash/_1019_ ),
    .A3(\hash/_1017_ ),
    .B1(\hash/_1049_ ),
    .Y(\hash/_1050_ ));
 sky130_fd_sc_hd__or2_2 \hash/_2227_  (.A(\hash/_1047_ ),
    .B(\hash/_1050_ ),
    .X(\hash/_1051_ ));
 sky130_fd_sc_hd__o41ai_1 \hash/_2228_  (.A1(\hash/_1803_ ),
    .A2(\hash/_1000_ ),
    .A3(\hash/_1021_ ),
    .A4(\hash/_1047_ ),
    .B1(\hash/_1051_ ),
    .Y(\hash/_1052_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2229_  (.A(\hash/_1814_ ),
    .B(\hash/_1052_ ),
    .Y(\hash/_0159_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2230_  (.A(\hash/_1814_ ),
    .B(\hash/_1025_ ),
    .C(\hash/_1048_ ),
    .X(\hash/_1053_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2231_  (.A(\hash/_1812_ ),
    .B(\hash/_1814_ ),
    .Y(\hash/_1054_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2232_  (.A1(\hash/_1814_ ),
    .A2(\hash/_1811_ ),
    .B1(\hash/_1813_ ),
    .Y(\hash/_1055_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2233_  (.A1(\hash/_1042_ ),
    .A2(\hash/_1054_ ),
    .B1(\hash/_1055_ ),
    .Y(\hash/_1056_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2234_  (.A1(\hash/_1020_ ),
    .A2(\hash/_1053_ ),
    .B1(\hash/_1056_ ),
    .Y(\hash/_1057_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2235_  (.A(\hash/_1816_ ),
    .B(\hash/_1057_ ),
    .Y(\hash/_0160_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2236_  (.A(\hash/_1814_ ),
    .B(\hash/_1816_ ),
    .Y(\hash/_1058_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2237_  (.A(\hash/_1058_ ),
    .B_N(\hash/_1051_ ),
    .Y(\hash/_1059_ ));
 sky130_fd_sc_hd__o41ai_1 \hash/_2238_  (.A1(\hash/_1803_ ),
    .A2(\hash/_1000_ ),
    .A3(\hash/_1021_ ),
    .A4(\hash/_1047_ ),
    .B1(\hash/_1059_ ),
    .Y(\hash/_1060_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2239_  (.A1(\hash/_1816_ ),
    .A2(\hash/_1813_ ),
    .B1(\hash/_1815_ ),
    .Y(\hash/_1061_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2240_  (.A(\hash/_1060_ ),
    .B(\hash/_1061_ ),
    .Y(\hash/_1062_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2241_  (.A(\hash/_1818_ ),
    .B(\hash/_1062_ ),
    .X(\hash/_0161_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2242_  (.A(\hash/_1816_ ),
    .B(\hash/_1818_ ),
    .Y(\hash/_1063_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2243_  (.A1(\hash/_1818_ ),
    .A2(\hash/_1815_ ),
    .B1(\hash/_1817_ ),
    .Y(\hash/_1064_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2244_  (.A1(\hash/_1057_ ),
    .A2(\hash/_1063_ ),
    .B1(\hash/_1064_ ),
    .Y(\hash/_1065_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2245_  (.A(\hash/_1820_ ),
    .B(\hash/_1065_ ),
    .X(\hash/_0162_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2246_  (.A(\hash/_1818_ ),
    .B(\hash/_1820_ ),
    .Y(\hash/_1066_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2247_  (.A1(\hash/_1820_ ),
    .A2(\hash/_1817_ ),
    .B1(\hash/_1819_ ),
    .Y(\hash/_1067_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2248_  (.A1(\hash/_1061_ ),
    .A2(\hash/_1066_ ),
    .B1(\hash/_1067_ ),
    .X(\hash/_1068_ ));
 sky130_fd_sc_hd__o31a_1 \hash/_2249_  (.A1(\hash/_1052_ ),
    .A2(\hash/_1058_ ),
    .A3(\hash/_1066_ ),
    .B1(\hash/_1068_ ),
    .X(\hash/_1069_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2250_  (.A(\hash/_1822_ ),
    .B(\hash/_1069_ ),
    .Y(\hash/_0163_ ));
 sky130_fd_sc_hd__and2_1 \hash/_2252_  (.A(\hash/_1820_ ),
    .B(\hash/_1822_ ),
    .X(\hash/_1071_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2253_  (.A1(\hash/_1822_ ),
    .A2(\hash/_1819_ ),
    .B1(\hash/_1821_ ),
    .Y(\hash/_1072_ ));
 sky130_fd_sc_hd__a21boi_1 \hash/_2254_  (.A1(\hash/_1065_ ),
    .A2(\hash/_1071_ ),
    .B1_N(\hash/_1072_ ),
    .Y(\hash/_1073_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2255_  (.A(\hash/_1824_ ),
    .B(\hash/_1073_ ),
    .Y(\hash/_0164_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2256_  (.A(\hash/_1826_ ),
    .Y(\hash/_1074_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2257_  (.A(\hash/_1822_ ),
    .B(\hash/_1824_ ),
    .Y(\hash/_1075_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2258_  (.A1(\hash/_1824_ ),
    .A2(\hash/_1821_ ),
    .B1(\hash/_1823_ ),
    .Y(\hash/_1076_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2259_  (.A1(\hash/_1069_ ),
    .A2(\hash/_1075_ ),
    .B1(\hash/_1076_ ),
    .Y(\hash/_1077_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2260_  (.A(\hash/_1074_ ),
    .B(\hash/_1077_ ),
    .Y(\hash/_0165_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2261_  (.A(\hash/_1072_ ),
    .B_N(\hash/_1824_ ),
    .Y(\hash/_1078_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2262_  (.A1(\hash/_1823_ ),
    .A2(\hash/_1078_ ),
    .B1(\hash/_1826_ ),
    .Y(\hash/_1079_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2263_  (.A_N(\hash/_1825_ ),
    .B(\hash/_1079_ ),
    .Y(\hash/_1080_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_2264_  (.A1(\hash/_1824_ ),
    .A2(\hash/_1826_ ),
    .A3(\hash/_1065_ ),
    .A4(\hash/_1071_ ),
    .B1(\hash/_1080_ ),
    .Y(\hash/_1081_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2265_  (.A(\hash/_1828_ ),
    .B(\hash/_1081_ ),
    .Y(\hash/_0166_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2266_  (.A(\hash/_1822_ ),
    .B(\hash/_1824_ ),
    .C(\hash/_1826_ ),
    .D(\hash/_1828_ ),
    .Y(\hash/_1082_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2267_  (.A1(\hash/_1074_ ),
    .A2(\hash/_1076_ ),
    .B1_N(\hash/_1825_ ),
    .Y(\hash/_1083_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2268_  (.A1(\hash/_1828_ ),
    .A2(\hash/_1083_ ),
    .B1(\hash/_1827_ ),
    .Y(\hash/_1084_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2269_  (.A1(\hash/_1069_ ),
    .A2(\hash/_1082_ ),
    .B1(\hash/_1084_ ),
    .Y(\hash/_1085_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2270_  (.A(\hash/_1830_ ),
    .B(\hash/_1085_ ),
    .X(\hash/_0167_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2271_  (.A_N(\hash/_1829_ ),
    .B(\hash/_1832_ ),
    .Y(\hash/_1086_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2272_  (.A(\hash/_1828_ ),
    .Y(\hash/_1087_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2273_  (.A1(\hash/_1826_ ),
    .A2(\hash/_1823_ ),
    .B1(\hash/_1825_ ),
    .Y(\hash/_1088_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2274_  (.A(\hash/_1827_ ),
    .Y(\hash/_1089_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2275_  (.A1(\hash/_1087_ ),
    .A2(\hash/_1088_ ),
    .B1(\hash/_1089_ ),
    .Y(\hash/_1090_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2276_  (.A1(\hash/_1830_ ),
    .A2(\hash/_1090_ ),
    .B1(\hash/_1829_ ),
    .Y(\hash/_1091_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2277_  (.A(\hash/_1090_ ),
    .B(\hash/_1086_ ),
    .Y(\hash/_1092_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2278_  (.A(\hash/_1832_ ),
    .B_N(\hash/_1830_ ),
    .Y(\hash/_1093_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2279_  (.A(\hash/_1820_ ),
    .B(\hash/_1822_ ),
    .Y(\hash/_1094_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2280_  (.A(\hash/_1824_ ),
    .B(\hash/_1826_ ),
    .C(\hash/_1828_ ),
    .Y(\hash/_1095_ ));
 sky130_fd_sc_hd__or3_1 \hash/_2281_  (.A(\hash/_1063_ ),
    .B(\hash/_1094_ ),
    .C(\hash/_1095_ ),
    .X(\hash/_1096_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2282_  (.A(\hash/_1064_ ),
    .B(\hash/_1095_ ),
    .Y(\hash/_1097_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2283_  (.A(\hash/_1072_ ),
    .B(\hash/_1095_ ),
    .Y(\hash/_1098_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2284_  (.A1(\hash/_1071_ ),
    .A2(\hash/_1097_ ),
    .B1(\hash/_1098_ ),
    .Y(\hash/_1099_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2285_  (.A1(\hash/_1057_ ),
    .A2(\hash/_1096_ ),
    .B1(\hash/_1099_ ),
    .Y(\hash/_1100_ ));
 sky130_fd_sc_hd__mux2i_1 \hash/_2286_  (.A0(\hash/_1092_ ),
    .A1(\hash/_1093_ ),
    .S(\hash/_1100_ ),
    .Y(\hash/_1101_ ));
 sky130_fd_sc_hd__o221ai_1 \hash/_2287_  (.A1(\hash/_1830_ ),
    .A2(\hash/_1086_ ),
    .B1(\hash/_1091_ ),
    .B2(\hash/_1832_ ),
    .C1(\hash/_1101_ ),
    .Y(\hash/_0168_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2288_  (.A1(\hash/_1060_ ),
    .A2(\hash/_1061_ ),
    .B1(\hash/_1066_ ),
    .Y(\hash/_1102_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2289_  (.A(\hash/_1830_ ),
    .B(\hash/_1832_ ),
    .Y(\hash/_1103_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2290_  (.A(\hash/_1082_ ),
    .B(\hash/_1103_ ),
    .Y(\hash/_1104_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2291_  (.A1(\hash/_1067_ ),
    .A2(\hash/_1075_ ),
    .B1(\hash/_1076_ ),
    .Y(\hash/_1105_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2292_  (.A1(\hash/_1826_ ),
    .A2(\hash/_1105_ ),
    .B1(\hash/_1825_ ),
    .Y(\hash/_1106_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2293_  (.A(\hash/_1087_ ),
    .B(\hash/_1106_ ),
    .Y(\hash/_1107_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2294_  (.A(\hash/_1827_ ),
    .B(\hash/_1107_ ),
    .Y(\hash/_1108_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2295_  (.A1(\hash/_1832_ ),
    .A2(\hash/_1829_ ),
    .B1(\hash/_1831_ ),
    .Y(\hash/_1109_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2296_  (.A1(\hash/_1108_ ),
    .A2(\hash/_1103_ ),
    .B1(\hash/_1109_ ),
    .Y(\hash/_1110_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2297_  (.A1(\hash/_1102_ ),
    .A2(\hash/_1104_ ),
    .B1(\hash/_1110_ ),
    .Y(\hash/_1111_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2298_  (.A(\hash/_1834_ ),
    .B(\hash/_1111_ ),
    .Y(\hash/_0169_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2299_  (.A(\hash/_1824_ ),
    .B(\hash/_1071_ ),
    .Y(\hash/_1112_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2300_  (.A(\hash/_1830_ ),
    .B(\hash/_1832_ ),
    .C(\hash/_1834_ ),
    .Y(\hash/_1113_ ));
 sky130_fd_sc_hd__nor4_1 \hash/_2301_  (.A(\hash/_1074_ ),
    .B(\hash/_1087_ ),
    .C(\hash/_1112_ ),
    .D(\hash/_1113_ ),
    .Y(\hash/_1114_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2302_  (.A(\hash/_1828_ ),
    .B(\hash/_1080_ ),
    .Y(\hash/_1115_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2303_  (.A1(\hash/_1830_ ),
    .A2(\hash/_1829_ ),
    .B1(\hash/_1832_ ),
    .Y(\hash/_1116_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2304_  (.A_N(\hash/_1831_ ),
    .B(\hash/_1116_ ),
    .Y(\hash/_1117_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2305_  (.A(\hash/_1834_ ),
    .B(\hash/_1117_ ),
    .Y(\hash/_1118_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2306_  (.A1(\hash/_1089_ ),
    .A2(\hash/_1109_ ),
    .A3(\hash/_1115_ ),
    .B1(\hash/_1118_ ),
    .Y(\hash/_1119_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_2307_  (.A1(\hash/_1065_ ),
    .A2(\hash/_1114_ ),
    .B1(\hash/_1119_ ),
    .C1(\hash/_1833_ ),
    .Y(\hash/_1120_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2308_  (.A(\hash/_1836_ ),
    .B(\hash/_1120_ ),
    .Y(\hash/_0171_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_2309_  (.A0(\hash/p2_cap[31] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2310_  (.A(_09577_),
    .B(\hash/p2_cap[31] ),
    .Y(\hash/_1121_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2311_  (.A(reset_hash_dash),
    .B(\hash/_1121_ ),
    .Y(\hash/_1122_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2312_  (.A(\hash/_1836_ ),
    .Y(\hash/_1123_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2313_  (.A1(\hash/_1084_ ),
    .A2(\hash/_1103_ ),
    .B1(\hash/_1109_ ),
    .Y(\hash/_1124_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2314_  (.A1(\hash/_1834_ ),
    .A2(\hash/_1124_ ),
    .B1(\hash/_1833_ ),
    .X(\hash/_1125_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2315_  (.A1(\hash/_1836_ ),
    .A2(\hash/_1125_ ),
    .B1(\hash/_1835_ ),
    .Y(\hash/_1126_ ));
 sky130_fd_sc_hd__o41ai_1 \hash/_2316_  (.A1(\hash/_1123_ ),
    .A2(\hash/_1069_ ),
    .A3(\hash/_1082_ ),
    .A4(\hash/_1113_ ),
    .B1(\hash/_1126_ ),
    .Y(\hash/_1127_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2317_  (.A(\hash/_1122_ ),
    .B(\hash/_1127_ ),
    .X(\hash/_0172_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2318_  (.A(\hash/_1474_ ),
    .B(\hash/_1842_ ),
    .X(\hash/_0200_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2319_  (.A1(\hash/_1473_ ),
    .A2(\hash/_1838_ ),
    .B1(\hash/_1837_ ),
    .X(\hash/_1128_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2320_  (.A1(\hash/_1842_ ),
    .A2(\hash/_1128_ ),
    .B1(\hash/_1841_ ),
    .X(\hash/_1129_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2321_  (.A(\hash/_1840_ ),
    .B(\hash/_1129_ ),
    .X(\hash/_0203_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2322_  (.A1(\hash/_1474_ ),
    .A2(\hash/_1842_ ),
    .B1(\hash/_1841_ ),
    .X(\hash/_1130_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2323_  (.A1(\hash/_1840_ ),
    .A2(\hash/_1130_ ),
    .B1(\hash/_1839_ ),
    .Y(\hash/_1131_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2324_  (.A(\hash/_1844_ ),
    .B(\hash/_1131_ ),
    .Y(\hash/_0204_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2325_  (.A1(\hash/_1840_ ),
    .A2(\hash/_1129_ ),
    .B1(\hash/_1839_ ),
    .Y(\hash/_1132_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2326_  (.A(\hash/_1132_ ),
    .B_N(\hash/_1844_ ),
    .Y(\hash/_1133_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2327_  (.A(\hash/_1843_ ),
    .B(\hash/_1133_ ),
    .Y(\hash/_1134_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2328_  (.A(\hash/_1846_ ),
    .B(\hash/_1134_ ),
    .Y(\hash/_0205_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_2329_  (.A1(\hash/_1474_ ),
    .A2(\hash/_1842_ ),
    .B1(\hash/_1839_ ),
    .C1(\hash/_1841_ ),
    .Y(\hash/_1135_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2330_  (.A1(\hash/_1840_ ),
    .A2(\hash/_1839_ ),
    .B1(\hash/_1844_ ),
    .Y(\hash/_1136_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2331_  (.A1(\hash/_1135_ ),
    .A2(\hash/_1136_ ),
    .B1_N(\hash/_1843_ ),
    .Y(\hash/_1137_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2332_  (.A1(\hash/_1846_ ),
    .A2(\hash/_1137_ ),
    .B1(\hash/_1845_ ),
    .Y(\hash/_1138_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2333_  (.A(\hash/_1848_ ),
    .B(\hash/_1138_ ),
    .Y(\hash/_0206_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2334_  (.A1(\hash/_1843_ ),
    .A2(\hash/_1133_ ),
    .B1(\hash/_1846_ ),
    .Y(\hash/_1139_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2335_  (.A_N(\hash/_1845_ ),
    .B(\hash/_1139_ ),
    .Y(\hash/_1140_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2336_  (.A1(\hash/_1848_ ),
    .A2(\hash/_1140_ ),
    .B1(\hash/_1847_ ),
    .Y(\hash/_1141_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2337_  (.A(\hash/_1850_ ),
    .B(\hash/_1141_ ),
    .Y(\hash/_0207_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2338_  (.A(\hash/_1848_ ),
    .Y(\hash/_1142_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2339_  (.A1(\hash/_1142_ ),
    .A2(\hash/_1138_ ),
    .B1_N(\hash/_1847_ ),
    .Y(\hash/_1143_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2340_  (.A1(\hash/_1850_ ),
    .A2(\hash/_1143_ ),
    .B1(\hash/_1849_ ),
    .Y(\hash/_1144_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2341_  (.A(\hash/_1852_ ),
    .B(\hash/_1144_ ),
    .Y(\hash/_0208_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2342_  (.A(\hash/_1848_ ),
    .B(\hash/_1850_ ),
    .C(\hash/_1852_ ),
    .Y(\hash/_1145_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2343_  (.A(\hash/_1844_ ),
    .B(\hash/_1846_ ),
    .Y(\hash/_1146_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2344_  (.A(\hash/_1145_ ),
    .B(\hash/_1146_ ),
    .Y(\hash/_1147_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2345_  (.A(\hash/_1846_ ),
    .B(\hash/_1843_ ),
    .Y(\hash/_1148_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2346_  (.A(\hash/_1844_ ),
    .B(\hash/_1846_ ),
    .C(\hash/_1839_ ),
    .Y(\hash/_1149_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2347_  (.A1(\hash/_1148_ ),
    .A2(\hash/_1149_ ),
    .B1(\hash/_1145_ ),
    .Y(\hash/_1150_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2348_  (.A1(\hash/_1840_ ),
    .A2(\hash/_1129_ ),
    .A3(\hash/_1147_ ),
    .B1(\hash/_1150_ ),
    .Y(\hash/_1151_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2349_  (.A1(\hash/_1848_ ),
    .A2(\hash/_1845_ ),
    .B1(\hash/_1847_ ),
    .X(\hash/_1152_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2350_  (.A1(\hash/_1850_ ),
    .A2(\hash/_1152_ ),
    .B1(\hash/_1849_ ),
    .X(\hash/_1153_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2351_  (.A1(\hash/_1852_ ),
    .A2(\hash/_1153_ ),
    .B1(\hash/_1851_ ),
    .Y(\hash/_1154_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2352_  (.A(\hash/_1151_ ),
    .B(\hash/_1154_ ),
    .Y(\hash/_1155_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2353_  (.A(\hash/_1854_ ),
    .B(\hash/_1155_ ),
    .X(\hash/_0209_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2354_  (.A(\hash/_1852_ ),
    .Y(\hash/_1156_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2355_  (.A1(\hash/_1156_ ),
    .A2(\hash/_1144_ ),
    .B1_N(\hash/_1851_ ),
    .Y(\hash/_1157_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2356_  (.A1(\hash/_1854_ ),
    .A2(\hash/_1157_ ),
    .B1(\hash/_1853_ ),
    .Y(\hash/_1158_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2357_  (.A(\hash/_1856_ ),
    .B(\hash/_1158_ ),
    .Y(\hash/_0180_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2358_  (.A1(\hash/_1856_ ),
    .A2(\hash/_1853_ ),
    .B1(\hash/_1855_ ),
    .Y(\hash/_1159_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2359_  (.A(\hash/_1854_ ),
    .B(\hash/_1856_ ),
    .C(\hash/_1155_ ),
    .Y(\hash/_1160_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2360_  (.A(\hash/_1159_ ),
    .B(\hash/_1160_ ),
    .Y(\hash/_1161_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2361_  (.A(\hash/_1858_ ),
    .B(\hash/_1161_ ),
    .X(\hash/_0181_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2362_  (.A(\hash/_1854_ ),
    .B(\hash/_1856_ ),
    .Y(\hash/_1162_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2363_  (.A1(\hash/_1850_ ),
    .A2(\hash/_1847_ ),
    .B1(\hash/_1849_ ),
    .X(\hash/_1163_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2364_  (.A1(\hash/_1852_ ),
    .A2(\hash/_1163_ ),
    .B1(\hash/_1851_ ),
    .Y(\hash/_1164_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2365_  (.A1(\hash/_1162_ ),
    .A2(\hash/_1164_ ),
    .B1(\hash/_1159_ ),
    .X(\hash/_1165_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_2366_  (.A1(\hash/_1138_ ),
    .A2(\hash/_1145_ ),
    .A3(\hash/_1162_ ),
    .B1(\hash/_1165_ ),
    .Y(\hash/_1166_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2367_  (.A1(\hash/_1858_ ),
    .A2(\hash/_1166_ ),
    .B1(\hash/_1857_ ),
    .Y(\hash/_1167_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2368_  (.A(\hash/_1860_ ),
    .B(\hash/_1167_ ),
    .Y(\hash/_0182_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2369_  (.A(\hash/_1858_ ),
    .B(\hash/_1860_ ),
    .Y(\hash/_1168_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2370_  (.A1(\hash/_1159_ ),
    .A2(\hash/_1162_ ),
    .B1(\hash/_1168_ ),
    .Y(\hash/_1169_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2371_  (.A1(\hash/_1860_ ),
    .A2(\hash/_1857_ ),
    .B1(\hash/_1859_ ),
    .Y(\hash/_1170_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2372_  (.A(\hash/_1169_ ),
    .B_N(\hash/_1170_ ),
    .Y(\hash/_1171_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2373_  (.A(\hash/_1159_ ),
    .B(\hash/_1170_ ),
    .Y(\hash/_1172_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_2374_  (.A1(\hash/_1852_ ),
    .A2(\hash/_1153_ ),
    .B1(\hash/_1172_ ),
    .C1(\hash/_1851_ ),
    .Y(\hash/_1173_ ));
 sky130_fd_sc_hd__and2_1 \hash/_2375_  (.A(\hash/_1151_ ),
    .B(\hash/_1173_ ),
    .X(\hash/_1174_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2376_  (.A(\hash/_1171_ ),
    .B(\hash/_1174_ ),
    .Y(\hash/_1175_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2377_  (.A(\hash/_1862_ ),
    .B(\hash/_1175_ ),
    .X(\hash/_0183_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2378_  (.A(\hash/_1860_ ),
    .B(\hash/_1862_ ),
    .Y(\hash/_1176_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2379_  (.A1(\hash/_1862_ ),
    .A2(\hash/_1859_ ),
    .B1(\hash/_1861_ ),
    .Y(\hash/_1177_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2380_  (.A1(\hash/_1167_ ),
    .A2(\hash/_1176_ ),
    .B1(\hash/_1177_ ),
    .Y(\hash/_1178_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2381_  (.A(\hash/_1864_ ),
    .B(\hash/_1178_ ),
    .X(\hash/_0184_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2382_  (.A(\hash/_1862_ ),
    .B(\hash/_1864_ ),
    .Y(\hash/_1179_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2383_  (.A1(\hash/_1864_ ),
    .A2(\hash/_1861_ ),
    .B1(\hash/_1863_ ),
    .Y(\hash/_1180_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_2384_  (.A1(\hash/_1171_ ),
    .A2(\hash/_1174_ ),
    .A3(\hash/_1179_ ),
    .B1(\hash/_1180_ ),
    .Y(\hash/_1181_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2385_  (.A(\hash/_1868_ ),
    .B(\hash/_1181_ ),
    .X(\hash/_0185_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2386_  (.A1(\hash/_1868_ ),
    .A2(\hash/_1863_ ),
    .B1(\hash/_1867_ ),
    .X(\hash/_1182_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2387_  (.A1(\hash/_1864_ ),
    .A2(\hash/_1868_ ),
    .A3(\hash/_1178_ ),
    .B1(\hash/_1182_ ),
    .Y(\hash/_1183_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2388_  (.A(\hash/_1866_ ),
    .B(\hash/_1183_ ),
    .Y(\hash/_0186_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2389_  (.A1(\hash/_1868_ ),
    .A2(\hash/_1181_ ),
    .B1(\hash/_1867_ ),
    .X(\hash/_1184_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2390_  (.A1(\hash/_1866_ ),
    .A2(\hash/_1184_ ),
    .B1(\hash/_1865_ ),
    .Y(\hash/_1185_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2391_  (.A(\hash/_1870_ ),
    .B(\hash/_1185_ ),
    .Y(\hash/_0187_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2392_  (.A(\hash/_1168_ ),
    .B(\hash/_1179_ ),
    .Y(\hash/_1186_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2393_  (.A(\hash/_1864_ ),
    .B(\hash/_1861_ ),
    .Y(\hash/_1187_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2394_  (.A1(\hash/_1170_ ),
    .A2(\hash/_1179_ ),
    .B1(\hash/_1187_ ),
    .Y(\hash/_1188_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2395_  (.A1(\hash/_1166_ ),
    .A2(\hash/_1186_ ),
    .B1(\hash/_1188_ ),
    .Y(\hash/_1189_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2396_  (.A(\hash/_1868_ ),
    .B(\hash/_1866_ ),
    .C(\hash/_1870_ ),
    .Y(\hash/_1190_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2397_  (.A1(\hash/_1866_ ),
    .A2(\hash/_1182_ ),
    .B1(\hash/_1865_ ),
    .X(\hash/_1191_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2398_  (.A1(\hash/_1870_ ),
    .A2(\hash/_1191_ ),
    .B1(\hash/_1869_ ),
    .Y(\hash/_1192_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2399_  (.A1(\hash/_1189_ ),
    .A2(\hash/_1190_ ),
    .B1(\hash/_1192_ ),
    .Y(\hash/_1193_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2400_  (.A(\hash/_1872_ ),
    .B(\hash/_1193_ ),
    .X(\hash/_0188_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2401_  (.A1(\hash/_1866_ ),
    .A2(\hash/_1867_ ),
    .B1(\hash/_1865_ ),
    .X(\hash/_1194_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2402_  (.A1(\hash/_1870_ ),
    .A2(\hash/_1194_ ),
    .B1(\hash/_1869_ ),
    .X(\hash/_1195_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2403_  (.A(\hash/_1868_ ),
    .B(\hash/_1866_ ),
    .C(\hash/_1870_ ),
    .D(\hash/_1872_ ),
    .Y(\hash/_1196_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2404_  (.A(\hash/_1180_ ),
    .B(\hash/_1196_ ),
    .Y(\hash/_1197_ ));
 sky130_fd_sc_hd__a211o_1 \hash/_2405_  (.A1(\hash/_1872_ ),
    .A2(\hash/_1195_ ),
    .B1(\hash/_1197_ ),
    .C1(\hash/_1871_ ),
    .X(\hash/_1198_ ));
 sky130_fd_sc_hd__a2111oi_1 \hash/_2406_  (.A1(\hash/_1151_ ),
    .A2(\hash/_1173_ ),
    .B1(\hash/_1179_ ),
    .C1(\hash/_1196_ ),
    .D1(\hash/_1171_ ),
    .Y(\hash/_1199_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2407_  (.A(\hash/_1198_ ),
    .B(\hash/_1199_ ),
    .Y(\hash/_1200_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2408_  (.A(\hash/_1874_ ),
    .B(\hash/_1200_ ),
    .Y(\hash/_0189_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2409_  (.A1(\hash/_1872_ ),
    .A2(\hash/_1193_ ),
    .B1(\hash/_1871_ ),
    .X(\hash/_1201_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2410_  (.A1(\hash/_1874_ ),
    .A2(\hash/_1201_ ),
    .B1(\hash/_1873_ ),
    .Y(\hash/_1202_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2411_  (.A(\hash/_1876_ ),
    .B(\hash/_1202_ ),
    .Y(\hash/_0190_ ));
 sky130_fd_sc_hd__or3_1 \hash/_2412_  (.A(\hash/_1873_ ),
    .B(\hash/_1875_ ),
    .C(\hash/_1198_ ),
    .X(\hash/_1203_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2413_  (.A(\hash/_1874_ ),
    .B(\hash/_1873_ ),
    .C(\hash/_1875_ ),
    .Y(\hash/_1204_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2414_  (.A(\hash/_1876_ ),
    .B(\hash/_1875_ ),
    .Y(\hash/_1205_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2415_  (.A(\hash/_1204_ ),
    .B(\hash/_1205_ ),
    .Y(\hash/_1206_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2416_  (.A1(\hash/_1199_ ),
    .A2(\hash/_1203_ ),
    .B1(\hash/_1206_ ),
    .Y(\hash/_1207_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2417_  (.A(\hash/_1878_ ),
    .B(\hash/_1207_ ),
    .Y(\hash/_0191_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2418_  (.A(\hash/_1880_ ),
    .Y(\hash/_1208_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2419_  (.A(\hash/_1872_ ),
    .B(\hash/_1874_ ),
    .C(\hash/_1876_ ),
    .Y(\hash/_1209_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2420_  (.A(\hash/_1874_ ),
    .B(\hash/_1876_ ),
    .C(\hash/_1871_ ),
    .X(\hash/_1210_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2421_  (.A1(\hash/_1876_ ),
    .A2(\hash/_1873_ ),
    .B1(\hash/_1210_ ),
    .Y(\hash/_1211_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2422_  (.A(\hash/_1875_ ),
    .B(\hash/_1877_ ),
    .Y(\hash/_1212_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2423_  (.A1(\hash/_1192_ ),
    .A2(\hash/_1209_ ),
    .B1(\hash/_1211_ ),
    .C1(\hash/_1212_ ),
    .Y(\hash/_1213_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_2424_  (.A1(\hash/_1166_ ),
    .A2(\hash/_1186_ ),
    .B1(\hash/_1188_ ),
    .C1(\hash/_1213_ ),
    .Y(\hash/_1214_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2425_  (.A1(\hash/_1192_ ),
    .A2(\hash/_1209_ ),
    .B1(\hash/_1211_ ),
    .Y(\hash/_1215_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2426_  (.A(\hash/_1874_ ),
    .B(\hash/_1876_ ),
    .Y(\hash/_1216_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2427_  (.A1(\hash/_1196_ ),
    .A2(\hash/_1216_ ),
    .B1(\hash/_1212_ ),
    .Y(\hash/_1217_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/_2428_  (.A1(\hash/_1878_ ),
    .A2(\hash/_1877_ ),
    .B1(\hash/_1215_ ),
    .B2(\hash/_1217_ ),
    .Y(\hash/_1218_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2429_  (.A(\hash/_1214_ ),
    .B(\hash/_1218_ ),
    .Y(\hash/_1219_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2430_  (.A(\hash/_1208_ ),
    .B(\hash/_1219_ ),
    .Y(\hash/_0192_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2431_  (.A1(\hash/_1199_ ),
    .A2(\hash/_1203_ ),
    .B1(\hash/_1206_ ),
    .C1(\hash/_1878_ ),
    .Y(\hash/_1220_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2432_  (.A(\hash/_1877_ ),
    .B_N(\hash/_1220_ ),
    .Y(\hash/_1221_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2433_  (.A1(\hash/_1208_ ),
    .A2(\hash/_1221_ ),
    .B1_N(\hash/_1879_ ),
    .Y(\hash/_1222_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2434_  (.A(\hash/_1882_ ),
    .B(\hash/_1222_ ),
    .X(\hash/_0193_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2435_  (.A1(\hash/_1882_ ),
    .A2(\hash/_1879_ ),
    .B1(\hash/_1881_ ),
    .Y(\hash/_1223_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2436_  (.A(\hash/_1880_ ),
    .B(\hash/_1882_ ),
    .Y(\hash/_1224_ ));
 sky130_fd_sc_hd__or3_1 \hash/_2437_  (.A(\hash/_1214_ ),
    .B(\hash/_1218_ ),
    .C(\hash/_1224_ ),
    .X(\hash/_1225_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2438_  (.A(\hash/_1223_ ),
    .B(\hash/_1225_ ),
    .Y(\hash/_1226_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2439_  (.A(\hash/_1884_ ),
    .B(\hash/_1226_ ),
    .X(\hash/_0194_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2440_  (.A1(\hash/_1884_ ),
    .A2(\hash/_1881_ ),
    .B1(\hash/_1883_ ),
    .X(\hash/_1227_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2441_  (.A1(\hash/_1882_ ),
    .A2(\hash/_1884_ ),
    .A3(\hash/_1222_ ),
    .B1(\hash/_1227_ ),
    .Y(\hash/_1228_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2442_  (.A(\hash/_1886_ ),
    .B(\hash/_1228_ ),
    .Y(\hash/_0195_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2443_  (.A(\hash/_1883_ ),
    .B(\hash/_1885_ ),
    .Y(\hash/_1229_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2444_  (.A(\hash/_1884_ ),
    .B(\hash/_1883_ ),
    .C(\hash/_1885_ ),
    .Y(\hash/_1230_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2445_  (.A(\hash/_1886_ ),
    .B(\hash/_1885_ ),
    .Y(\hash/_1231_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/_2446_  (.A1(\hash/_1223_ ),
    .A2(\hash/_1225_ ),
    .A3(\hash/_1229_ ),
    .B1(\hash/_1230_ ),
    .C1(\hash/_1231_ ),
    .Y(\hash/_1232_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2447_  (.A(\hash/_1888_ ),
    .B(\hash/_1232_ ),
    .X(\hash/_0196_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2448_  (.A(\hash/_1882_ ),
    .B(\hash/_1884_ ),
    .Y(\hash/_1233_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2449_  (.A(\hash/_1886_ ),
    .B(\hash/_1888_ ),
    .Y(\hash/_1234_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2450_  (.A(\hash/_1233_ ),
    .B(\hash/_1234_ ),
    .Y(\hash/_1235_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2451_  (.A1(\hash/_1886_ ),
    .A2(\hash/_1227_ ),
    .B1(\hash/_1885_ ),
    .X(\hash/_1236_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2452_  (.A1(\hash/_1888_ ),
    .A2(\hash/_1236_ ),
    .B1(\hash/_1887_ ),
    .X(\hash/_1237_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2453_  (.A1(\hash/_1222_ ),
    .A2(\hash/_1235_ ),
    .B1(\hash/_1237_ ),
    .Y(\hash/_1238_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2454_  (.A(\hash/_1890_ ),
    .B(\hash/_1238_ ),
    .Y(\hash/_0197_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2455_  (.A1(\hash/_1886_ ),
    .A2(\hash/_1883_ ),
    .B1(\hash/_1885_ ),
    .X(\hash/_1239_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2456_  (.A1(\hash/_1888_ ),
    .A2(\hash/_1239_ ),
    .B1(\hash/_1887_ ),
    .X(\hash/_1240_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2457_  (.A(\hash/_1884_ ),
    .B(\hash/_1890_ ),
    .Y(\hash/_1241_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2458_  (.A(\hash/_1234_ ),
    .B(\hash/_1241_ ),
    .Y(\hash/_1242_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/_2459_  (.A1(\hash/_1890_ ),
    .A2(\hash/_1240_ ),
    .B1(\hash/_1242_ ),
    .B2(\hash/_1226_ ),
    .C1(\hash/_1889_ ),
    .Y(\hash/_1243_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2460_  (.A(\hash/_1892_ ),
    .B(\hash/_1243_ ),
    .Y(\hash/_0198_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2461_  (.A(\hash/_1890_ ),
    .B(\hash/_1892_ ),
    .C(\hash/_1235_ ),
    .X(\hash/_1244_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2462_  (.A(\hash/_1880_ ),
    .B(\hash/_1244_ ),
    .Y(\hash/_1245_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2463_  (.A1(\hash/_1880_ ),
    .A2(\hash/_1877_ ),
    .B1(\hash/_1879_ ),
    .Y(\hash/_1246_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2464_  (.A1(\hash/_1233_ ),
    .A2(\hash/_1246_ ),
    .B1_N(\hash/_1227_ ),
    .Y(\hash/_1247_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2465_  (.A1(\hash/_1886_ ),
    .A2(\hash/_1247_ ),
    .B1(\hash/_1885_ ),
    .Y(\hash/_1248_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2466_  (.A(\hash/_1248_ ),
    .B_N(\hash/_1888_ ),
    .Y(\hash/_1249_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2467_  (.A1(\hash/_1887_ ),
    .A2(\hash/_1249_ ),
    .B1(\hash/_1890_ ),
    .Y(\hash/_1250_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2468_  (.A_N(\hash/_1889_ ),
    .B(\hash/_1250_ ),
    .Y(\hash/_1251_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2469_  (.A1(\hash/_1892_ ),
    .A2(\hash/_1251_ ),
    .B1(\hash/_1891_ ),
    .Y(\hash/_1252_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2470_  (.A1(\hash/_1220_ ),
    .A2(\hash/_1245_ ),
    .B1(\hash/_1252_ ),
    .Y(\hash/_1253_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2471_  (.A(\hash/_1894_ ),
    .B(\hash/_1253_ ),
    .X(\hash/_0199_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2472_  (.A1(\hash/_1890_ ),
    .A2(\hash/_1237_ ),
    .B1(\hash/_1889_ ),
    .X(\hash/_1254_ ));
 sky130_fd_sc_hd__a221o_1 \hash/_2473_  (.A1(\hash/_1879_ ),
    .A2(\hash/_1244_ ),
    .B1(\hash/_1254_ ),
    .B2(\hash/_1892_ ),
    .C1(\hash/_1891_ ),
    .X(\hash/_1255_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2474_  (.A(\hash/_1214_ ),
    .B(\hash/_1218_ ),
    .C(\hash/_1245_ ),
    .Y(\hash/_1256_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2475_  (.A1(\hash/_1255_ ),
    .A2(\hash/_1256_ ),
    .B1(\hash/_1894_ ),
    .X(\hash/_1257_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2476_  (.A(\hash/_1893_ ),
    .B(\hash/_1257_ ),
    .Y(\hash/_1258_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2477_  (.A(\hash/_1896_ ),
    .B(\hash/_1258_ ),
    .Y(\hash/_0201_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_2478_  (.A0(\hash/e_cap[31] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[31] ));
 sky130_fd_sc_hd__nand2_1 \hash/_2479_  (.A(\hash/_1894_ ),
    .B(\hash/_1896_ ),
    .Y(\hash/_1259_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2480_  (.A(\hash/_1894_ ),
    .B(\hash/_1896_ ),
    .C(\hash/_1255_ ),
    .Y(\hash/_1260_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2481_  (.A1(\hash/_1896_ ),
    .A2(\hash/_1893_ ),
    .B1(\hash/_1895_ ),
    .Y(\hash/_1261_ ));
 sky130_fd_sc_hd__o311ai_1 \hash/_2482_  (.A1(\hash/_1221_ ),
    .A2(\hash/_1245_ ),
    .A3(\hash/_1259_ ),
    .B1(\hash/_1260_ ),
    .C1(\hash/_1261_ ),
    .Y(\hash/_1262_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2483_  (.A(_09578_),
    .B(\hash/e_cap[31] ),
    .Y(\hash/_1263_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2484_  (.A(reset_hash_dash),
    .B(\hash/_1263_ ),
    .Y(\hash/_1264_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2485_  (.A(\hash/_1262_ ),
    .B(\hash/_1264_ ),
    .X(\hash/_0202_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2486_  (.A(\hash/_1476_ ),
    .B(\hash/_1902_ ),
    .X(\hash/_0230_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2487_  (.A1(\hash/_1475_ ),
    .A2(\hash/_1898_ ),
    .B1(\hash/_1897_ ),
    .X(\hash/_1265_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2488_  (.A1(\hash/_1902_ ),
    .A2(\hash/_1265_ ),
    .B1(\hash/_1901_ ),
    .Y(\hash/_1266_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2489_  (.A(\hash/_1900_ ),
    .B(\hash/_1266_ ),
    .Y(\hash/_0233_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2490_  (.A1(\hash/_1476_ ),
    .A2(\hash/_1902_ ),
    .B1(\hash/_1901_ ),
    .X(\hash/_1267_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2491_  (.A1(\hash/_1900_ ),
    .A2(\hash/_1267_ ),
    .B1(\hash/_1899_ ),
    .Y(\hash/_1268_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2492_  (.A(\hash/_1904_ ),
    .B(\hash/_1268_ ),
    .Y(\hash/_0234_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2493_  (.A(\hash/_1904_ ),
    .Y(\hash/_1269_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2494_  (.A(\hash/_1266_ ),
    .B_N(\hash/_1900_ ),
    .Y(\hash/_1270_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2495_  (.A(\hash/_1899_ ),
    .B(\hash/_1270_ ),
    .Y(\hash/_1271_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2496_  (.A(\hash/_1269_ ),
    .B(\hash/_1271_ ),
    .Y(\hash/_1272_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2497_  (.A(\hash/_1903_ ),
    .B(\hash/_1272_ ),
    .Y(\hash/_1273_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2498_  (.A(\hash/_1906_ ),
    .B(\hash/_1273_ ),
    .Y(\hash/_0235_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2499_  (.A1(\hash/_1269_ ),
    .A2(\hash/_1268_ ),
    .B1_N(\hash/_1903_ ),
    .Y(\hash/_1274_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2500_  (.A1(\hash/_1906_ ),
    .A2(\hash/_1274_ ),
    .B1(\hash/_1905_ ),
    .Y(\hash/_1275_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2501_  (.A(\hash/_1908_ ),
    .B(\hash/_1275_ ),
    .Y(\hash/_0236_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2502_  (.A(\hash/_1906_ ),
    .Y(\hash/_1276_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2503_  (.A1(\hash/_1276_ ),
    .A2(\hash/_1273_ ),
    .B1_N(\hash/_1905_ ),
    .Y(\hash/_1277_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2504_  (.A1(\hash/_1908_ ),
    .A2(\hash/_1277_ ),
    .B1(\hash/_1907_ ),
    .Y(\hash/_1278_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2505_  (.A(\hash/_1910_ ),
    .B(\hash/_1278_ ),
    .Y(\hash/_0237_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2506_  (.A(\hash/_1908_ ),
    .Y(\hash/_1279_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2507_  (.A1(\hash/_1279_ ),
    .A2(\hash/_1275_ ),
    .B1_N(\hash/_1907_ ),
    .Y(\hash/_1280_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2508_  (.A1(\hash/_1910_ ),
    .A2(\hash/_1280_ ),
    .B1(\hash/_1909_ ),
    .Y(\hash/_1281_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2509_  (.A(\hash/_1912_ ),
    .B(\hash/_1281_ ),
    .Y(\hash/_0238_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2510_  (.A(\hash/_1908_ ),
    .B(\hash/_1910_ ),
    .C(\hash/_1912_ ),
    .Y(\hash/_1282_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2511_  (.A(\hash/_1269_ ),
    .B(\hash/_1276_ ),
    .C(\hash/_1282_ ),
    .Y(\hash/_1283_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2512_  (.A(\hash/_1906_ ),
    .B(\hash/_1903_ ),
    .Y(\hash/_1284_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2513_  (.A(\hash/_1904_ ),
    .B(\hash/_1906_ ),
    .C(\hash/_1899_ ),
    .Y(\hash/_1285_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2514_  (.A1(\hash/_1284_ ),
    .A2(\hash/_1285_ ),
    .B1(\hash/_1282_ ),
    .Y(\hash/_1286_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2515_  (.A1(\hash/_1270_ ),
    .A2(\hash/_1283_ ),
    .B1(\hash/_1286_ ),
    .X(\hash/_1287_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2516_  (.A1(\hash/_1908_ ),
    .A2(\hash/_1905_ ),
    .B1(\hash/_1907_ ),
    .X(\hash/_1288_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2517_  (.A1(\hash/_1910_ ),
    .A2(\hash/_1288_ ),
    .B1(\hash/_1909_ ),
    .X(\hash/_1289_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2518_  (.A1(\hash/_1912_ ),
    .A2(\hash/_1289_ ),
    .B1(\hash/_1911_ ),
    .Y(\hash/_1290_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2519_  (.A(\hash/_1287_ ),
    .B_N(\hash/_1290_ ),
    .Y(\hash/_1291_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2520_  (.A(\hash/_1914_ ),
    .B(\hash/_1291_ ),
    .Y(\hash/_0239_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2521_  (.A(\hash/_1912_ ),
    .Y(\hash/_1292_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2522_  (.A1(\hash/_1292_ ),
    .A2(\hash/_1281_ ),
    .B1_N(\hash/_1911_ ),
    .Y(\hash/_1293_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2523_  (.A1(\hash/_1914_ ),
    .A2(\hash/_1293_ ),
    .B1(\hash/_1913_ ),
    .Y(\hash/_1294_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2524_  (.A(\hash/_1916_ ),
    .B(\hash/_1294_ ),
    .Y(\hash/_0210_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2525_  (.A(\hash/_1913_ ),
    .B(\hash/_1915_ ),
    .Y(\hash/_1295_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2526_  (.A(\hash/_1290_ ),
    .B(\hash/_1295_ ),
    .Y(\hash/_1296_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2527_  (.A1(\hash/_1914_ ),
    .A2(\hash/_1913_ ),
    .B1(\hash/_1916_ ),
    .X(\hash/_1297_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2528_  (.A(\hash/_1915_ ),
    .B(\hash/_1297_ ),
    .Y(\hash/_1298_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2529_  (.A(\hash/_1298_ ),
    .Y(\hash/_1299_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2530_  (.A1(\hash/_1287_ ),
    .A2(\hash/_1296_ ),
    .B1(\hash/_1299_ ),
    .Y(\hash/_1300_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2531_  (.A(\hash/_1918_ ),
    .B(\hash/_1300_ ),
    .Y(\hash/_0211_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2532_  (.A(\hash/_1903_ ),
    .B(\hash/_1905_ ),
    .Y(\hash/_1301_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2533_  (.A1(\hash/_1269_ ),
    .A2(\hash/_1268_ ),
    .B1(\hash/_1301_ ),
    .X(\hash/_1302_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2534_  (.A(\hash/_1914_ ),
    .B(\hash/_1916_ ),
    .Y(\hash/_1303_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2535_  (.A(\hash/_1282_ ),
    .B(\hash/_1303_ ),
    .Y(\hash/_1304_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2536_  (.A1(\hash/_1906_ ),
    .A2(\hash/_1905_ ),
    .B1(\hash/_1304_ ),
    .Y(\hash/_1305_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2537_  (.A(\hash/_1303_ ),
    .Y(\hash/_1306_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2538_  (.A1(\hash/_1910_ ),
    .A2(\hash/_1907_ ),
    .B1(\hash/_1909_ ),
    .Y(\hash/_1307_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2539_  (.A1(\hash/_1292_ ),
    .A2(\hash/_1307_ ),
    .B1_N(\hash/_1911_ ),
    .Y(\hash/_1308_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/_2540_  (.A1(\hash/_1916_ ),
    .A2(\hash/_1913_ ),
    .B1(\hash/_1306_ ),
    .B2(\hash/_1308_ ),
    .C1(\hash/_1915_ ),
    .Y(\hash/_1309_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2541_  (.A1(\hash/_1302_ ),
    .A2(\hash/_1305_ ),
    .B1(\hash/_1309_ ),
    .Y(\hash/_1310_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2542_  (.A1(\hash/_1918_ ),
    .A2(\hash/_1310_ ),
    .B1(\hash/_1917_ ),
    .Y(\hash/_1311_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2543_  (.A(\hash/_1920_ ),
    .B(\hash/_1311_ ),
    .Y(\hash/_0212_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2544_  (.A1(\hash/_1287_ ),
    .A2(\hash/_1296_ ),
    .B1(\hash/_1299_ ),
    .C1(\hash/_1918_ ),
    .Y(\hash/_1312_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2545_  (.A_N(\hash/_1917_ ),
    .B(\hash/_1312_ ),
    .Y(\hash/_1313_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2546_  (.A1(\hash/_1920_ ),
    .A2(\hash/_1313_ ),
    .B1(\hash/_1919_ ),
    .Y(\hash/_1314_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2547_  (.A(\hash/_1922_ ),
    .B(\hash/_1314_ ),
    .Y(\hash/_0213_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2548_  (.A(\hash/_1920_ ),
    .B(\hash/_1922_ ),
    .Y(\hash/_1315_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2549_  (.A(\hash/_1918_ ),
    .B(\hash/_1917_ ),
    .Y(\hash/_1316_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2550_  (.A(\hash/_1922_ ),
    .B(\hash/_1919_ ),
    .Y(\hash/_1317_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2551_  (.A1(\hash/_1315_ ),
    .A2(\hash/_1316_ ),
    .B1(\hash/_1317_ ),
    .Y(\hash/_1318_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2552_  (.A(\hash/_1917_ ),
    .B(\hash/_1919_ ),
    .Y(\hash/_1319_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2553_  (.A1(\hash/_1302_ ),
    .A2(\hash/_1305_ ),
    .B1(\hash/_1309_ ),
    .C1(\hash/_1319_ ),
    .Y(\hash/_1320_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2554_  (.A1(\hash/_1318_ ),
    .A2(\hash/_1320_ ),
    .B1(\hash/_1921_ ),
    .Y(\hash/_1321_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2555_  (.A(\hash/_1924_ ),
    .B(\hash/_1321_ ),
    .Y(\hash/_0214_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2556_  (.A(\hash/_1920_ ),
    .B(\hash/_1922_ ),
    .C(\hash/_1917_ ),
    .Y(\hash/_1322_ ));
 sky130_fd_sc_hd__and2_1 \hash/_2557_  (.A(\hash/_1317_ ),
    .B(\hash/_1322_ ),
    .X(\hash/_1323_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_2558_  (.A1(\hash/_1312_ ),
    .A2(\hash/_1315_ ),
    .B1(\hash/_1323_ ),
    .X(\hash/_1324_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2559_  (.A_N(\hash/_1921_ ),
    .B(\hash/_1324_ ),
    .Y(\hash/_1325_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2560_  (.A1(\hash/_1924_ ),
    .A2(\hash/_1325_ ),
    .B1(\hash/_1923_ ),
    .Y(\hash/_1326_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2561_  (.A(\hash/_1928_ ),
    .B(\hash/_1326_ ),
    .Y(\hash/_0215_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2562_  (.A(\hash/_1318_ ),
    .B(\hash/_1320_ ),
    .Y(\hash/_1327_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2563_  (.A(\hash/_1921_ ),
    .B(\hash/_1923_ ),
    .Y(\hash/_1328_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2564_  (.A1(\hash/_1924_ ),
    .A2(\hash/_1923_ ),
    .B1(\hash/_1928_ ),
    .Y(\hash/_1329_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2565_  (.A1(\hash/_1327_ ),
    .A2(\hash/_1328_ ),
    .B1(\hash/_1329_ ),
    .Y(\hash/_1330_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2566_  (.A(\hash/_1927_ ),
    .B(\hash/_1330_ ),
    .Y(\hash/_1331_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2567_  (.A(\hash/_1926_ ),
    .B(\hash/_1331_ ),
    .Y(\hash/_0216_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2568_  (.A1(\hash/_1928_ ),
    .A2(\hash/_1923_ ),
    .B1(\hash/_1927_ ),
    .X(\hash/_1332_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2569_  (.A1(\hash/_1926_ ),
    .A2(\hash/_1332_ ),
    .B1(\hash/_1925_ ),
    .X(\hash/_1333_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_2570_  (.A1(\hash/_1924_ ),
    .A2(\hash/_1928_ ),
    .A3(\hash/_1926_ ),
    .A4(\hash/_1325_ ),
    .B1(\hash/_1333_ ),
    .Y(\hash/_1334_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2571_  (.A(\hash/_1930_ ),
    .B(\hash/_1334_ ),
    .Y(\hash/_0217_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2572_  (.A(\hash/_1932_ ),
    .Y(\hash/_1335_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2573_  (.A(\hash/_1924_ ),
    .B(\hash/_1928_ ),
    .C(\hash/_1926_ ),
    .D(\hash/_1930_ ),
    .Y(\hash/_1336_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2574_  (.A1(\hash/_1930_ ),
    .A2(\hash/_1333_ ),
    .B1(\hash/_1929_ ),
    .Y(\hash/_1337_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2575_  (.A1(\hash/_1321_ ),
    .A2(\hash/_1336_ ),
    .B1(\hash/_1337_ ),
    .Y(\hash/_1338_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2576_  (.A(\hash/_1335_ ),
    .B(\hash/_1338_ ),
    .Y(\hash/_0218_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2577_  (.A1(\hash/_1926_ ),
    .A2(\hash/_1927_ ),
    .B1(\hash/_1925_ ),
    .X(\hash/_1339_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2578_  (.A1(\hash/_1930_ ),
    .A2(\hash/_1339_ ),
    .B1(\hash/_1929_ ),
    .Y(\hash/_1340_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2579_  (.A(\hash/_1335_ ),
    .B(\hash/_1340_ ),
    .Y(\hash/_1341_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2580_  (.A(\hash/_1931_ ),
    .B(\hash/_1341_ ),
    .Y(\hash/_1342_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2581_  (.A(\hash/_1926_ ),
    .B(\hash/_1930_ ),
    .C(\hash/_1932_ ),
    .Y(\hash/_1343_ ));
 sky130_fd_sc_hd__or2_2 \hash/_2582_  (.A(\hash/_1329_ ),
    .B(\hash/_1343_ ),
    .X(\hash/_1344_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2583_  (.A(\hash/_1342_ ),
    .B(\hash/_1344_ ),
    .Y(\hash/_1345_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2584_  (.A(\hash/_1323_ ),
    .B(\hash/_1328_ ),
    .C(\hash/_1342_ ),
    .X(\hash/_1346_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2585_  (.A1(\hash/_1312_ ),
    .A2(\hash/_1315_ ),
    .B1(\hash/_1346_ ),
    .Y(\hash/_1347_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2586_  (.A(\hash/_1345_ ),
    .B(\hash/_1347_ ),
    .Y(\hash/_1348_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2587_  (.A(\hash/_1934_ ),
    .B(\hash/_1348_ ),
    .Y(\hash/_0219_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2588_  (.A1(\hash/_1932_ ),
    .A2(\hash/_1338_ ),
    .B1(\hash/_1931_ ),
    .X(\hash/_1349_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2589_  (.A1(\hash/_1934_ ),
    .A2(\hash/_1349_ ),
    .B1(\hash/_1933_ ),
    .Y(\hash/_1350_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2590_  (.A(\hash/_1936_ ),
    .B(\hash/_1350_ ),
    .Y(\hash/_0220_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2591_  (.A1(\hash/_1936_ ),
    .A2(\hash/_1933_ ),
    .B1(\hash/_1935_ ),
    .Y(\hash/_1351_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2592_  (.A(\hash/_1934_ ),
    .B(\hash/_1936_ ),
    .Y(\hash/_1352_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2593_  (.A(\hash/_1351_ ),
    .B(\hash/_1352_ ),
    .Y(\hash/_1353_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2594_  (.A(\hash/_1342_ ),
    .B(\hash/_1344_ ),
    .C(\hash/_1351_ ),
    .Y(\hash/_1354_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2595_  (.A(\hash/_1353_ ),
    .B(\hash/_1354_ ),
    .Y(\hash/_1355_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_2596_  (.A1(\hash/_1324_ ),
    .A2(\hash/_1328_ ),
    .A3(\hash/_1342_ ),
    .A4(\hash/_1351_ ),
    .B1(\hash/_1355_ ),
    .Y(\hash/_1356_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2597_  (.A(\hash/_1938_ ),
    .B(\hash/_1356_ ),
    .X(\hash/_0221_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2598_  (.A(\hash/_1343_ ),
    .B(\hash/_1352_ ),
    .Y(\hash/_1357_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2599_  (.A(\hash/_1924_ ),
    .B(\hash/_1928_ ),
    .C(\hash/_1938_ ),
    .D(\hash/_1357_ ),
    .Y(\hash/_1358_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2600_  (.A(\hash/_1931_ ),
    .B(\hash/_1933_ ),
    .C(\hash/_1935_ ),
    .Y(\hash/_1359_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2601_  (.A1(\hash/_1335_ ),
    .A2(\hash/_1337_ ),
    .B1(\hash/_1359_ ),
    .Y(\hash/_1360_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2602_  (.A1(\hash/_1938_ ),
    .A2(\hash/_1353_ ),
    .A3(\hash/_1360_ ),
    .B1(\hash/_1937_ ),
    .Y(\hash/_1361_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2603_  (.A1(\hash/_1321_ ),
    .A2(\hash/_1358_ ),
    .B1(\hash/_1361_ ),
    .Y(\hash/_1362_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2604_  (.A(\hash/_1940_ ),
    .B(\hash/_1362_ ),
    .X(\hash/_0222_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2605_  (.A(\hash/_1938_ ),
    .B(\hash/_1940_ ),
    .Y(\hash/_1363_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2606_  (.A(\hash/_1352_ ),
    .B(\hash/_1363_ ),
    .Y(\hash/_1364_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2607_  (.A(\hash/_1351_ ),
    .B_N(\hash/_1938_ ),
    .Y(\hash/_1365_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2608_  (.A1(\hash/_1937_ ),
    .A2(\hash/_1365_ ),
    .B1(\hash/_1940_ ),
    .Y(\hash/_1366_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2609_  (.A_N(\hash/_1939_ ),
    .B(\hash/_1366_ ),
    .Y(\hash/_1367_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2610_  (.A1(\hash/_1345_ ),
    .A2(\hash/_1347_ ),
    .A3(\hash/_1364_ ),
    .B1(\hash/_1367_ ),
    .Y(\hash/_1368_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2611_  (.A(\hash/_1942_ ),
    .B(\hash/_1368_ ),
    .Y(\hash/_0223_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2612_  (.A(\hash/_1944_ ),
    .Y(\hash/_1369_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2613_  (.A1(\hash/_1942_ ),
    .A2(\hash/_1939_ ),
    .B1(\hash/_1941_ ),
    .Y(\hash/_1370_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2614_  (.A(\hash/_1940_ ),
    .B(\hash/_1942_ ),
    .C(\hash/_1362_ ),
    .Y(\hash/_1371_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2615_  (.A(\hash/_1370_ ),
    .B(\hash/_1371_ ),
    .Y(\hash/_1372_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2616_  (.A(\hash/_1369_ ),
    .B(\hash/_1372_ ),
    .Y(\hash/_0224_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2617_  (.A(\hash/_1946_ ),
    .Y(\hash/_1373_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2618_  (.A(\hash/_1942_ ),
    .B(\hash/_1944_ ),
    .Y(\hash/_1374_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2619_  (.A1(\hash/_1944_ ),
    .A2(\hash/_1941_ ),
    .B1(\hash/_1943_ ),
    .Y(\hash/_1375_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2620_  (.A1(\hash/_1368_ ),
    .A2(\hash/_1374_ ),
    .B1(\hash/_1375_ ),
    .Y(\hash/_1376_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2621_  (.A(\hash/_1373_ ),
    .B(\hash/_1376_ ),
    .Y(\hash/_0225_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2622_  (.A(\hash/_1948_ ),
    .Y(\hash/_1377_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2623_  (.A(\hash/_1944_ ),
    .B(\hash/_1946_ ),
    .Y(\hash/_1378_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2624_  (.A1(\hash/_1369_ ),
    .A2(\hash/_1370_ ),
    .B1_N(\hash/_1943_ ),
    .Y(\hash/_1379_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2625_  (.A1(\hash/_1946_ ),
    .A2(\hash/_1379_ ),
    .B1(\hash/_1945_ ),
    .Y(\hash/_1380_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2626_  (.A1(\hash/_1371_ ),
    .A2(\hash/_1378_ ),
    .B1(\hash/_1380_ ),
    .Y(\hash/_1381_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2627_  (.A(\hash/_1377_ ),
    .B(\hash/_1381_ ),
    .Y(\hash/_0226_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2628_  (.A(\hash/_1942_ ),
    .B(\hash/_1944_ ),
    .C(\hash/_1946_ ),
    .D(\hash/_1948_ ),
    .Y(\hash/_1382_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2629_  (.A1(\hash/_1373_ ),
    .A2(\hash/_1375_ ),
    .B1_N(\hash/_1945_ ),
    .Y(\hash/_1383_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2630_  (.A1(\hash/_1948_ ),
    .A2(\hash/_1383_ ),
    .B1(\hash/_1947_ ),
    .Y(\hash/_1384_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2631_  (.A1(\hash/_1368_ ),
    .A2(\hash/_1382_ ),
    .B1(\hash/_1384_ ),
    .Y(\hash/_1385_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2632_  (.A(\hash/_1950_ ),
    .B(\hash/_1385_ ),
    .X(\hash/_0227_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2633_  (.A(\hash/_1944_ ),
    .B(\hash/_1946_ ),
    .C(\hash/_1948_ ),
    .Y(\hash/_1386_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2634_  (.A1(\hash/_1950_ ),
    .A2(\hash/_1949_ ),
    .B1(\hash/_1940_ ),
    .C1(\hash/_1942_ ),
    .Y(\hash/_1387_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2635_  (.A(\hash/_1386_ ),
    .B(\hash/_1387_ ),
    .Y(\hash/_1388_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2636_  (.A1(\hash/_1946_ ),
    .A2(\hash/_1943_ ),
    .B1(\hash/_1945_ ),
    .Y(\hash/_1389_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2637_  (.A(\hash/_1947_ ),
    .B(\hash/_1949_ ),
    .Y(\hash/_1390_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2638_  (.A1(\hash/_1377_ ),
    .A2(\hash/_1389_ ),
    .B1(\hash/_1390_ ),
    .Y(\hash/_1391_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2639_  (.A(\hash/_1370_ ),
    .B(\hash/_1386_ ),
    .Y(\hash/_1392_ ));
 sky130_fd_sc_hd__o22a_1 \hash/_2640_  (.A1(\hash/_1950_ ),
    .A2(\hash/_1949_ ),
    .B1(\hash/_1391_ ),
    .B2(\hash/_1392_ ),
    .X(\hash/_1393_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2641_  (.A1(\hash/_1362_ ),
    .A2(\hash/_1388_ ),
    .B1(\hash/_1393_ ),
    .Y(\hash/_1394_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2642_  (.A(\hash/_1952_ ),
    .B(\hash/_1394_ ),
    .Y(\hash/_0228_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2643_  (.A(\hash/_1950_ ),
    .B(\hash/_1952_ ),
    .Y(\hash/_1395_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_2644_  (.A(\hash/_1363_ ),
    .B(\hash/_1382_ ),
    .C(\hash/_1395_ ),
    .Y(\hash/_1396_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2645_  (.A1(\hash/_1940_ ),
    .A2(\hash/_1937_ ),
    .B1(\hash/_1939_ ),
    .Y(\hash/_1397_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2646_  (.A1(\hash/_1374_ ),
    .A2(\hash/_1397_ ),
    .B1(\hash/_1375_ ),
    .Y(\hash/_1398_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2647_  (.A1(\hash/_1946_ ),
    .A2(\hash/_1398_ ),
    .B1(\hash/_1945_ ),
    .Y(\hash/_1399_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2648_  (.A(\hash/_1377_ ),
    .B(\hash/_1399_ ),
    .Y(\hash/_1400_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2649_  (.A(\hash/_1947_ ),
    .B(\hash/_1400_ ),
    .Y(\hash/_1401_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2650_  (.A1(\hash/_1952_ ),
    .A2(\hash/_1949_ ),
    .B1(\hash/_1951_ ),
    .Y(\hash/_1402_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2651_  (.A1(\hash/_1401_ ),
    .A2(\hash/_1395_ ),
    .B1(\hash/_1402_ ),
    .Y(\hash/_1403_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2652_  (.A1(\hash/_1356_ ),
    .A2(\hash/_1396_ ),
    .B1(\hash/_1403_ ),
    .Y(\hash/_1404_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2653_  (.A(\hash/_1954_ ),
    .B(\hash/_1404_ ),
    .Y(\hash/_0229_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2654_  (.A(\hash/_1956_ ),
    .Y(\hash/_1405_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_2655_  (.A(\hash/_1950_ ),
    .B(\hash/_1952_ ),
    .C(\hash/_1954_ ),
    .Y(\hash/_1406_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2656_  (.A(\hash/_1947_ ),
    .Y(\hash/_1407_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2657_  (.A1(\hash/_1377_ ),
    .A2(\hash/_1380_ ),
    .B1(\hash/_1402_ ),
    .C1(\hash/_1407_ ),
    .Y(\hash/_1408_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2658_  (.A1(\hash/_1950_ ),
    .A2(\hash/_1949_ ),
    .B1(\hash/_1952_ ),
    .Y(\hash/_1409_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2659_  (.A_N(\hash/_1951_ ),
    .B(\hash/_1409_ ),
    .Y(\hash/_1410_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2660_  (.A1(\hash/_1954_ ),
    .A2(\hash/_1408_ ),
    .A3(\hash/_1410_ ),
    .B1(\hash/_1953_ ),
    .Y(\hash/_1411_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_2661_  (.A1(\hash/_1371_ ),
    .A2(\hash/_1386_ ),
    .A3(\hash/_1406_ ),
    .B1(\hash/_1411_ ),
    .Y(\hash/_1412_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2662_  (.A(\hash/_1405_ ),
    .B(\hash/_1412_ ),
    .Y(\hash/_0231_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_2663_  (.A0(\hash/f_cap[31] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2664_  (.A(_09578_),
    .B(\hash/f_cap[31] ),
    .Y(\hash/_1413_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2665_  (.A(reset_hash_dash),
    .B(\hash/_1413_ ),
    .Y(\hash/_1414_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2666_  (.A1(\hash/_1384_ ),
    .A2(\hash/_1395_ ),
    .B1(\hash/_1402_ ),
    .Y(\hash/_1415_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2667_  (.A1(\hash/_1954_ ),
    .A2(\hash/_1415_ ),
    .B1(\hash/_1953_ ),
    .X(\hash/_1416_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2668_  (.A1(\hash/_1956_ ),
    .A2(\hash/_1416_ ),
    .B1(\hash/_1955_ ),
    .Y(\hash/_1417_ ));
 sky130_fd_sc_hd__o41ai_1 \hash/_2669_  (.A1(\hash/_1405_ ),
    .A2(\hash/_1368_ ),
    .A3(\hash/_1382_ ),
    .A4(\hash/_1406_ ),
    .B1(\hash/_1417_ ),
    .Y(\hash/_1418_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2670_  (.A(\hash/_1414_ ),
    .B(\hash/_1418_ ),
    .X(\hash/_0232_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_2671_  (.A0(\hash/a_new[0] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2672_  (.A0(\hash/a_new[10] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2673_  (.A0(\hash/a_new[11] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2674_  (.A0(\hash/a_new[12] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2676_  (.A0(\hash/a_new[13] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2677_  (.A0(\hash/a_new[14] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2678_  (.A0(\hash/a_new[15] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2679_  (.A0(\hash/a_new[16] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2680_  (.A0(\hash/a_new[17] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2681_  (.A0(\hash/a_new[18] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2682_  (.A0(\hash/a_new[19] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2683_  (.A0(\hash/a_new[1] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2684_  (.A0(\hash/a_new[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2685_  (.A0(\hash/a_new[21] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2687_  (.A0(\hash/a_new[22] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2688_  (.A0(\hash/a_new[23] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2689_  (.A0(\hash/a_new[24] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2690_  (.A0(\hash/a_new[25] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2691_  (.A0(\hash/a_new[26] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2692_  (.A0(\hash/a_new[27] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2693_  (.A0(\hash/a_new[28] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2694_  (.A0(\hash/a_new[29] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2695_  (.A0(\hash/a_new[2] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2696_  (.A0(\hash/a_new[30] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2698_  (.A0(\hash/a_new[3] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2699_  (.A0(\hash/a_new[4] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2700_  (.A0(\hash/a_new[5] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2701_  (.A0(\hash/a_new[6] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2702_  (.A0(\hash/a_new[7] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2703_  (.A0(\hash/a_new[8] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2704_  (.A0(\hash/a_new[9] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/a[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2705_  (.A0(\hash/b_new[0] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2706_  (.A0(\hash/b_new[10] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2707_  (.A0(\hash/b_new[11] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2709_  (.A0(\hash/b_new[12] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2710_  (.A0(\hash/b_new[13] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2711_  (.A0(\hash/b_new[14] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2712_  (.A0(\hash/b_new[15] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2713_  (.A0(\hash/b_new[16] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2714_  (.A0(\hash/b_new[17] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2715_  (.A0(\hash/b_new[18] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2716_  (.A0(\hash/b_new[19] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2717_  (.A0(\hash/b_new[1] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2718_  (.A0(\hash/b_new[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2721_  (.A0(\hash/b_new[21] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2722_  (.A0(\hash/b_new[22] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2723_  (.A0(\hash/b_new[23] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2724_  (.A0(\hash/b_new[24] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2725_  (.A0(\hash/b_new[25] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2726_  (.A0(\hash/b_new[26] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2727_  (.A0(\hash/b_new[27] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2728_  (.A0(\hash/b_new[28] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2729_  (.A0(\hash/b_new[29] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2730_  (.A0(\hash/b_new[2] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2732_  (.A0(\hash/b_new[30] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2733_  (.A0(\hash/b_new[3] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2734_  (.A0(\hash/b_new[4] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2735_  (.A0(\hash/b_new[5] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2736_  (.A0(\hash/b_new[6] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2737_  (.A0(\hash/b_new[7] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2738_  (.A0(\hash/b_new[8] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/b[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2739_  (.A0(\hash/b_new[9] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2740_  (.A0(\hash/a_cap[0] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2741_  (.A0(\hash/a_cap[10] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2743_  (.A0(\hash/a_cap[11] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2744_  (.A0(\hash/a_cap[12] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2745_  (.A0(\hash/a_cap[13] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2746_  (.A0(\hash/a_cap[14] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2747_  (.A0(\hash/a_cap[15] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2748_  (.A0(\hash/a_cap[16] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2749_  (.A0(\hash/a_cap[17] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2750_  (.A0(\hash/a_cap[18] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2751_  (.A0(\hash/a_cap[19] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2752_  (.A0(\hash/a_cap[1] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2754_  (.A0(\hash/a_cap[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2755_  (.A0(\hash/a_cap[21] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2756_  (.A0(\hash/a_cap[22] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2757_  (.A0(\hash/a_cap[23] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2758_  (.A0(\hash/a_cap[24] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2759_  (.A0(\hash/a_cap[25] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2760_  (.A0(\hash/a_cap[26] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2761_  (.A0(\hash/a_cap[27] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2762_  (.A0(\hash/a_cap[28] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2763_  (.A0(\hash/a_cap[29] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2765_  (.A0(\hash/a_cap[2] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2766_  (.A0(\hash/a_cap[30] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2767_  (.A0(\hash/a_cap[3] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2768_  (.A0(\hash/a_cap[4] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2769_  (.A0(\hash/a_cap[5] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2770_  (.A0(\hash/a_cap[6] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2771_  (.A0(\hash/a_cap[7] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2772_  (.A0(\hash/a_cap[8] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2773_  (.A0(\hash/a_cap[9] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/c[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2774_  (.A0(\hash/b_cap[0] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2776_  (.A0(\hash/b_cap[10] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2777_  (.A0(\hash/b_cap[11] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2778_  (.A0(\hash/b_cap[12] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2779_  (.A0(\hash/b_cap[13] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2780_  (.A0(\hash/b_cap[14] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2781_  (.A0(\hash/b_cap[15] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2782_  (.A0(\hash/b_cap[16] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2783_  (.A0(\hash/b_cap[17] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2784_  (.A0(\hash/b_cap[18] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2785_  (.A0(\hash/b_cap[19] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2787_  (.A0(\hash/b_cap[1] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2788_  (.A0(\hash/b_cap[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2789_  (.A0(\hash/b_cap[21] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2790_  (.A0(\hash/b_cap[22] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2791_  (.A0(\hash/b_cap[23] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2792_  (.A0(\hash/b_cap[24] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2793_  (.A0(\hash/b_cap[25] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2794_  (.A0(\hash/b_cap[26] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2795_  (.A0(\hash/b_cap[27] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2796_  (.A0(\hash/b_cap[28] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2798_  (.A0(\hash/b_cap[29] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2799_  (.A0(\hash/b_cap[2] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2800_  (.A0(\hash/b_cap[30] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2801_  (.A0(\hash/b_cap[3] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2802_  (.A0(\hash/b_cap[4] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2803_  (.A0(\hash/b_cap[5] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2804_  (.A0(\hash/b_cap[6] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2805_  (.A0(\hash/b_cap[7] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2806_  (.A0(\hash/b_cap[8] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2807_  (.A0(\hash/b_cap[9] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/d[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2809_  (.A0(\hash/e_new[0] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2810_  (.A0(\hash/e_new[10] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2811_  (.A0(\hash/e_new[11] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2812_  (.A0(\hash/e_new[12] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2813_  (.A0(\hash/e_new[13] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2814_  (.A0(\hash/e_new[14] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2815_  (.A0(\hash/e_new[15] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2816_  (.A0(\hash/e_new[16] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2817_  (.A0(\hash/e_new[17] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2818_  (.A0(\hash/e_new[18] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2820_  (.A0(\hash/e_new[19] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2821_  (.A0(\hash/e_new[1] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2822_  (.A0(\hash/e_new[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2823_  (.A0(\hash/e_new[21] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2824_  (.A0(\hash/e_new[22] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2825_  (.A0(\hash/e_new[23] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2826_  (.A0(\hash/e_new[24] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2827_  (.A0(\hash/e_new[25] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2828_  (.A0(\hash/e_new[26] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2829_  (.A0(\hash/e_new[27] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2832_  (.A0(\hash/e_new[28] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2833_  (.A0(\hash/e_new[29] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2834_  (.A0(\hash/e_new[2] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2835_  (.A0(\hash/e_new[30] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2836_  (.A0(\hash/e_new[3] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2837_  (.A0(\hash/e_new[4] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2838_  (.A0(\hash/e_new[5] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2839_  (.A0(\hash/e_new[6] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2840_  (.A0(\hash/e_new[7] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2841_  (.A0(\hash/e_new[8] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/e[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2843_  (.A0(\hash/e_new[9] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/e[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2844_  (.A0(\hash/p2_cap[0] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2845_  (.A0(\hash/p2_cap[10] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2846_  (.A0(\hash/p2_cap[11] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2847_  (.A0(\hash/p2_cap[12] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2848_  (.A0(\hash/p2_cap[13] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2849_  (.A0(\hash/p2_cap[14] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2850_  (.A0(\hash/p2_cap[15] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2851_  (.A0(\hash/p2_cap[16] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2852_  (.A0(\hash/p2_cap[17] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2854_  (.A0(\hash/p2_cap[18] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2855_  (.A0(\hash/p2_cap[19] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2856_  (.A0(\hash/p2_cap[1] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2857_  (.A0(\hash/p2_cap[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2858_  (.A0(\hash/p2_cap[21] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2859_  (.A0(\hash/p2_cap[22] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2860_  (.A0(\hash/p2_cap[23] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2861_  (.A0(\hash/p2_cap[24] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2862_  (.A0(\hash/p2_cap[25] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2863_  (.A0(\hash/p2_cap[26] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2865_  (.A0(\hash/p2_cap[27] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2866_  (.A0(\hash/p2_cap[28] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2867_  (.A0(\hash/p2_cap[29] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2868_  (.A0(\hash/p2_cap[2] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2869_  (.A0(\hash/p2_cap[30] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2870_  (.A0(\hash/p2_cap[3] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2871_  (.A0(\hash/p2_cap[4] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2872_  (.A0(\hash/p2_cap[5] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2873_  (.A0(\hash/p2_cap[6] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2874_  (.A0(\hash/p2_cap[7] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/f[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2876_  (.A0(\hash/p2_cap[8] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2877_  (.A0(\hash/p2_cap[9] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/f[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2878_  (.A0(\hash/e_cap[0] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2879_  (.A0(\hash/e_cap[10] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2880_  (.A0(\hash/e_cap[11] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2881_  (.A0(\hash/e_cap[12] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2882_  (.A0(\hash/e_cap[13] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2883_  (.A0(\hash/e_cap[14] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2884_  (.A0(\hash/e_cap[15] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2885_  (.A0(\hash/e_cap[16] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2887_  (.A0(\hash/e_cap[17] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2888_  (.A0(\hash/e_cap[18] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2889_  (.A0(\hash/e_cap[19] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2890_  (.A0(\hash/e_cap[1] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2891_  (.A0(\hash/e_cap[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2892_  (.A0(\hash/e_cap[21] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2893_  (.A0(\hash/e_cap[22] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2894_  (.A0(\hash/e_cap[23] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2895_  (.A0(\hash/e_cap[24] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2896_  (.A0(\hash/e_cap[25] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2898_  (.A0(\hash/e_cap[26] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2899_  (.A0(\hash/e_cap[27] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2900_  (.A0(\hash/e_cap[28] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2901_  (.A0(\hash/e_cap[29] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2902_  (.A0(\hash/e_cap[2] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2903_  (.A0(\hash/e_cap[30] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2904_  (.A0(\hash/e_cap[3] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2905_  (.A0(\hash/e_cap[4] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2906_  (.A0(\hash/e_cap[5] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2907_  (.A0(\hash/e_cap[6] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2909_  (.A0(\hash/e_cap[7] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2910_  (.A0(\hash/e_cap[8] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/g[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2911_  (.A0(\hash/e_cap[9] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/g[9] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2912_  (.A0(\hash/f_cap[0] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[0] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2913_  (.A0(\hash/f_cap[10] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[10] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2914_  (.A0(\hash/f_cap[11] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[11] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2915_  (.A0(\hash/f_cap[12] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[12] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2916_  (.A0(\hash/f_cap[13] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[13] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2917_  (.A0(\hash/f_cap[14] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[14] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2918_  (.A0(\hash/f_cap[15] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[15] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2920_  (.A0(\hash/f_cap[16] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[16] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2921_  (.A0(\hash/f_cap[17] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[17] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2922_  (.A0(\hash/f_cap[18] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[18] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2923_  (.A0(\hash/f_cap[19] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[19] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2924_  (.A0(\hash/f_cap[1] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[1] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2925_  (.A0(\hash/f_cap[20] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[20] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2926_  (.A0(\hash/f_cap[21] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[21] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2927_  (.A0(\hash/f_cap[22] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[22] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2928_  (.A0(\hash/f_cap[23] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[23] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2929_  (.A0(\hash/f_cap[24] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[24] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2931_  (.A0(\hash/f_cap[25] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[25] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2932_  (.A0(\hash/f_cap[26] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[26] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2933_  (.A0(\hash/f_cap[27] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[27] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2934_  (.A0(\hash/f_cap[28] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[28] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2935_  (.A0(\hash/f_cap[29] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[29] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2936_  (.A0(\hash/f_cap[2] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[2] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2937_  (.A0(\hash/f_cap[30] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[30] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2938_  (.A0(\hash/f_cap[3] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[3] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2939_  (.A0(\hash/f_cap[4] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[4] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2940_  (.A0(\hash/f_cap[5] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[5] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2941_  (.A0(\hash/f_cap[6] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[6] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2942_  (.A0(\hash/f_cap[7] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[7] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2943_  (.A0(\hash/f_cap[8] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/h[8] ));
 sky130_fd_sc_hd__mux2_2 \hash/_2944_  (.A0(\hash/f_cap[9] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/h[9] ));
 sky130_fd_sc_hd__xor2_1 \hash/_2945_  (.A(\hash/_1462_ ),
    .B(\hash/_1482_ ),
    .X(\hash/_0020_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2946_  (.A1(\hash/_1461_ ),
    .A2(\hash/_1478_ ),
    .B1(\hash/_1477_ ),
    .X(\hash/_0240_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2947_  (.A1(\hash/_1482_ ),
    .A2(\hash/_0240_ ),
    .B1(\hash/_1481_ ),
    .Y(\hash/_0241_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2948_  (.A(\hash/_1480_ ),
    .B(\hash/_0241_ ),
    .Y(\hash/_0023_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2949_  (.A1(\hash/_1462_ ),
    .A2(\hash/_1482_ ),
    .B1(\hash/_1481_ ),
    .Y(\hash/_0242_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2950_  (.A(\hash/_0242_ ),
    .Y(\hash/_0243_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2951_  (.A1(\hash/_1480_ ),
    .A2(\hash/_0243_ ),
    .B1(\hash/_1479_ ),
    .Y(\hash/_0244_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2952_  (.A(\hash/_1484_ ),
    .B(\hash/_0244_ ),
    .Y(\hash/_0024_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2953_  (.A(\hash/_1480_ ),
    .B(\hash/_1484_ ),
    .Y(\hash/_0245_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2954_  (.A1(\hash/_1484_ ),
    .A2(\hash/_1479_ ),
    .B1(\hash/_1483_ ),
    .Y(\hash/_0246_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2955_  (.A1(\hash/_0241_ ),
    .A2(\hash/_0245_ ),
    .B1(\hash/_0246_ ),
    .Y(\hash/_0247_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_2956_  (.A(\hash/_1486_ ),
    .B(\hash/_0247_ ),
    .X(\hash/_0025_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2957_  (.A1(\hash/_0242_ ),
    .A2(\hash/_0245_ ),
    .B1(\hash/_0246_ ),
    .Y(\hash/_0248_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2958_  (.A1(\hash/_1486_ ),
    .A2(\hash/_0248_ ),
    .B1(\hash/_1485_ ),
    .Y(\hash/_0249_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2959_  (.A(\hash/_1488_ ),
    .B(\hash/_0249_ ),
    .Y(\hash/_0026_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2960_  (.A1(\hash/_1486_ ),
    .A2(\hash/_0247_ ),
    .B1(\hash/_1485_ ),
    .X(\hash/_0250_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2961_  (.A1(\hash/_1488_ ),
    .A2(\hash/_0250_ ),
    .B1(\hash/_1487_ ),
    .Y(\hash/_0251_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2962_  (.A(\hash/_1490_ ),
    .B(\hash/_0251_ ),
    .Y(\hash/_0027_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2963_  (.A(\hash/_1485_ ),
    .B(\hash/_1487_ ),
    .Y(\hash/_0252_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_2964_  (.A1(\hash/_0242_ ),
    .A2(\hash/_0245_ ),
    .B1(\hash/_0252_ ),
    .C1(\hash/_0246_ ),
    .Y(\hash/_0253_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2965_  (.A(\hash/_1487_ ),
    .Y(\hash/_0254_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_2966_  (.A1(\hash/_1486_ ),
    .A2(\hash/_1485_ ),
    .B1(\hash/_1488_ ),
    .Y(\hash/_0255_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2967_  (.A(\hash/_0254_ ),
    .B(\hash/_0255_ ),
    .Y(\hash/_0256_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_2968_  (.A1(\hash/_1490_ ),
    .A2(\hash/_0253_ ),
    .A3(\hash/_0256_ ),
    .B1(\hash/_1489_ ),
    .Y(\hash/_0257_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2969_  (.A(\hash/_1492_ ),
    .B(\hash/_0257_ ),
    .Y(\hash/_0028_ ));
 sky130_fd_sc_hd__and3_1 \hash/_2970_  (.A(\hash/_1488_ ),
    .B(\hash/_1490_ ),
    .C(\hash/_1492_ ),
    .X(\hash/_0258_ ));
 sky130_fd_sc_hd__inv_1 \hash/_2971_  (.A(\hash/_1492_ ),
    .Y(\hash/_0259_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2972_  (.A1(\hash/_1488_ ),
    .A2(\hash/_1485_ ),
    .B1(\hash/_1487_ ),
    .X(\hash/_0260_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2973_  (.A1(\hash/_1490_ ),
    .A2(\hash/_0260_ ),
    .B1(\hash/_1489_ ),
    .Y(\hash/_0261_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2974_  (.A(\hash/_0259_ ),
    .B(\hash/_0261_ ),
    .Y(\hash/_0262_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/_2975_  (.A1(\hash/_1486_ ),
    .A2(\hash/_0247_ ),
    .A3(\hash/_0258_ ),
    .B1(\hash/_0262_ ),
    .C1(\hash/_1491_ ),
    .Y(\hash/_0263_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2976_  (.A(\hash/_1494_ ),
    .B(\hash/_0263_ ),
    .Y(\hash/_0029_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_2977_  (.A1(\hash/_0259_ ),
    .A2(\hash/_0257_ ),
    .B1_N(\hash/_1491_ ),
    .Y(\hash/_0264_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2978_  (.A1(\hash/_1494_ ),
    .A2(\hash/_0264_ ),
    .B1(\hash/_1493_ ),
    .Y(\hash/_0265_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2979_  (.A(\hash/_1496_ ),
    .B(\hash/_0265_ ),
    .Y(\hash/_0000_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_2980_  (.A1(\hash/_1494_ ),
    .A2(\hash/_1493_ ),
    .B1(\hash/_1496_ ),
    .Y(\hash/_0266_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_2981_  (.A_N(\hash/_1495_ ),
    .B(\hash/_0266_ ),
    .Y(\hash/_0267_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_2982_  (.A(\hash/_1493_ ),
    .B(\hash/_1495_ ),
    .Y(\hash/_0268_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2983_  (.A(\hash/_0263_ ),
    .B(\hash/_0268_ ),
    .Y(\hash/_0269_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_2984_  (.A(\hash/_0267_ ),
    .B(\hash/_0269_ ),
    .Y(\hash/_0270_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2985_  (.A(\hash/_1498_ ),
    .B(\hash/_0270_ ),
    .Y(\hash/_0001_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_2986_  (.A(\hash/_1494_ ),
    .B(\hash/_1496_ ),
    .C(\hash/_1490_ ),
    .D(\hash/_1492_ ),
    .Y(\hash/_0271_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2987_  (.A1(\hash/_0254_ ),
    .A2(\hash/_0255_ ),
    .B1(\hash/_0271_ ),
    .Y(\hash/_0272_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2988_  (.A1(\hash/_1492_ ),
    .A2(\hash/_1489_ ),
    .B1(\hash/_1491_ ),
    .X(\hash/_0273_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2989_  (.A1(\hash/_1494_ ),
    .A2(\hash/_0273_ ),
    .B1(\hash/_1493_ ),
    .X(\hash/_0274_ ));
 sky130_fd_sc_hd__a221o_1 \hash/_2990_  (.A1(\hash/_0253_ ),
    .A2(\hash/_0272_ ),
    .B1(\hash/_0274_ ),
    .B2(\hash/_1496_ ),
    .C1(\hash/_1495_ ),
    .X(\hash/_0275_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_2991_  (.A1(\hash/_1498_ ),
    .A2(\hash/_0275_ ),
    .B1(\hash/_1497_ ),
    .Y(\hash/_0276_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2992_  (.A(\hash/_1500_ ),
    .B(\hash/_0276_ ),
    .Y(\hash/_0002_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2994_  (.A1(\hash/_1500_ ),
    .A2(\hash/_1497_ ),
    .B1(\hash/_1499_ ),
    .X(\hash/_0278_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_2995_  (.A1(\hash/_1498_ ),
    .A2(\hash/_1500_ ),
    .A3(\hash/_0267_ ),
    .A4(\hash/_0269_ ),
    .B1(\hash/_0278_ ),
    .Y(\hash/_0279_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_2996_  (.A(\hash/_1502_ ),
    .B(\hash/_0279_ ),
    .Y(\hash/_0003_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_2998_  (.A(\hash/_0276_ ),
    .B_N(\hash/_1500_ ),
    .Y(\hash/_0281_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_2999_  (.A1(\hash/_1502_ ),
    .A2(\hash/_1499_ ),
    .B1(\hash/_1501_ ),
    .X(\hash/_0282_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3000_  (.A1(\hash/_1502_ ),
    .A2(\hash/_0281_ ),
    .B1(\hash/_0282_ ),
    .Y(\hash/_0283_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3001_  (.A(\hash/_1504_ ),
    .B(\hash/_0283_ ),
    .Y(\hash/_0004_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3003_  (.A(\hash/_1498_ ),
    .B(\hash/_1500_ ),
    .C(\hash/_1502_ ),
    .D(\hash/_1504_ ),
    .Y(\hash/_0285_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3004_  (.A(\hash/_1500_ ),
    .B(\hash/_1502_ ),
    .C(\hash/_1504_ ),
    .D(\hash/_1497_ ),
    .Y(\hash/_0286_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3005_  (.A1(\hash/_1504_ ),
    .A2(\hash/_0282_ ),
    .B1(\hash/_1503_ ),
    .Y(\hash/_0287_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_3006_  (.A1(\hash/_0270_ ),
    .A2(\hash/_0285_ ),
    .B1(\hash/_0286_ ),
    .C1(\hash/_0287_ ),
    .Y(\hash/_0288_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3007_  (.A(\hash/_1508_ ),
    .B(\hash/_0288_ ),
    .X(\hash/_0005_ ));
 sky130_fd_sc_hd__and4_1 \hash/_3009_  (.A(\hash/_1498_ ),
    .B(\hash/_1500_ ),
    .C(\hash/_1502_ ),
    .D(\hash/_1504_ ),
    .X(\hash/_0290_ ));
 sky130_fd_sc_hd__a21boi_1 \hash/_3010_  (.A1(\hash/_0275_ ),
    .A2(\hash/_0290_ ),
    .B1_N(\hash/_0286_ ),
    .Y(\hash/_0291_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3011_  (.A(\hash/_0287_ ),
    .B(\hash/_0291_ ),
    .Y(\hash/_0292_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3012_  (.A1(\hash/_1508_ ),
    .A2(\hash/_0292_ ),
    .B1(\hash/_1507_ ),
    .Y(\hash/_0293_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3013_  (.A(\hash/_1506_ ),
    .B(\hash/_0293_ ),
    .Y(\hash/_0006_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3014_  (.A(\hash/_1502_ ),
    .B(\hash/_1504_ ),
    .C(\hash/_1508_ ),
    .D(\hash/_1506_ ),
    .Y(\hash/_0294_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3015_  (.A1(\hash/_1504_ ),
    .A2(\hash/_1501_ ),
    .B1(\hash/_1503_ ),
    .X(\hash/_0295_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3016_  (.A1(\hash/_1508_ ),
    .A2(\hash/_0295_ ),
    .B1(\hash/_1507_ ),
    .X(\hash/_0296_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3017_  (.A1(\hash/_1506_ ),
    .A2(\hash/_0296_ ),
    .B1(\hash/_1505_ ),
    .Y(\hash/_0297_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3018_  (.A1(\hash/_0279_ ),
    .A2(\hash/_0294_ ),
    .B1(\hash/_0297_ ),
    .Y(\hash/_0298_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3019_  (.A(\hash/_1510_ ),
    .B(\hash/_0298_ ),
    .X(\hash/_0007_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3020_  (.A(\hash/_1504_ ),
    .B(\hash/_1508_ ),
    .C(\hash/_1506_ ),
    .Y(\hash/_0299_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3021_  (.A1(\hash/_1508_ ),
    .A2(\hash/_1503_ ),
    .B1(\hash/_1507_ ),
    .X(\hash/_0300_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3022_  (.A1(\hash/_1506_ ),
    .A2(\hash/_0300_ ),
    .B1(\hash/_1505_ ),
    .Y(\hash/_0301_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3023_  (.A1(\hash/_0283_ ),
    .A2(\hash/_0299_ ),
    .B1(\hash/_0301_ ),
    .Y(\hash/_0302_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3024_  (.A1(\hash/_1510_ ),
    .A2(\hash/_0302_ ),
    .B1(\hash/_1509_ ),
    .Y(\hash/_0303_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3025_  (.A(\hash/_1512_ ),
    .B(\hash/_0303_ ),
    .Y(\hash/_0008_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3026_  (.A(\hash/_1508_ ),
    .B(\hash/_1506_ ),
    .Y(\hash/_0304_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3027_  (.A(\hash/_1510_ ),
    .B(\hash/_1512_ ),
    .Y(\hash/_0305_ ));
 sky130_fd_sc_hd__nor4b_1 \hash/_3028_  (.A(\hash/_0285_ ),
    .B(\hash/_0304_ ),
    .C(\hash/_0305_ ),
    .D_N(\hash/_0267_ ),
    .Y(\hash/_0306_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3029_  (.A1(\hash/_1502_ ),
    .A2(\hash/_0278_ ),
    .B1(\hash/_1501_ ),
    .X(\hash/_0307_ ));
 sky130_fd_sc_hd__a2111oi_0 \hash/_3030_  (.A1(\hash/_1504_ ),
    .A2(\hash/_0307_ ),
    .B1(\hash/_1507_ ),
    .C1(\hash/_1505_ ),
    .D1(\hash/_1503_ ),
    .Y(\hash/_0308_ ));
 sky130_fd_sc_hd__or3_1 \hash/_3031_  (.A(\hash/_1508_ ),
    .B(\hash/_1505_ ),
    .C(\hash/_1507_ ),
    .X(\hash/_0309_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3032_  (.A1(\hash/_1506_ ),
    .A2(\hash/_1505_ ),
    .B1(\hash/_0309_ ),
    .Y(\hash/_0310_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3033_  (.A1(\hash/_1512_ ),
    .A2(\hash/_1509_ ),
    .B1(\hash/_1511_ ),
    .Y(\hash/_0311_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_3034_  (.A1(\hash/_0305_ ),
    .A2(\hash/_0308_ ),
    .A3(\hash/_0310_ ),
    .B1(\hash/_0311_ ),
    .Y(\hash/_0312_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3035_  (.A1(\hash/_0269_ ),
    .A2(\hash/_0306_ ),
    .B1(\hash/_0312_ ),
    .Y(\hash/_0313_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3036_  (.A(\hash/_1514_ ),
    .B(\hash/_0313_ ),
    .Y(\hash/_0009_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3037_  (.A1(\hash/_1510_ ),
    .A2(\hash/_1505_ ),
    .B1(\hash/_1509_ ),
    .X(\hash/_0314_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3038_  (.A1(\hash/_1512_ ),
    .A2(\hash/_0314_ ),
    .B1(\hash/_1511_ ),
    .Y(\hash/_0315_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3039_  (.A(\hash/_0287_ ),
    .B(\hash/_0315_ ),
    .Y(\hash/_0316_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3040_  (.A(\hash/_1507_ ),
    .B(\hash/_0316_ ),
    .Y(\hash/_0317_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3041_  (.A(\hash/_1506_ ),
    .B(\hash/_1510_ ),
    .C(\hash/_1512_ ),
    .Y(\hash/_0318_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3042_  (.A(\hash/_1508_ ),
    .B(\hash/_1507_ ),
    .Y(\hash/_0319_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3043_  (.A1(\hash/_0318_ ),
    .A2(\hash/_0319_ ),
    .B1(\hash/_0315_ ),
    .X(\hash/_0320_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3044_  (.A1(\hash/_0291_ ),
    .A2(\hash/_0317_ ),
    .B1(\hash/_0320_ ),
    .Y(\hash/_0321_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3045_  (.A1(\hash/_1514_ ),
    .A2(\hash/_0321_ ),
    .B1(\hash/_1513_ ),
    .Y(\hash/_0322_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3046_  (.A(\hash/_1516_ ),
    .B(\hash/_0322_ ),
    .Y(\hash/_0010_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3047_  (.A(\hash/_1491_ ),
    .B(\hash/_1493_ ),
    .C(\hash/_1495_ ),
    .Y(\hash/_0323_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3048_  (.A1(\hash/_0259_ ),
    .A2(\hash/_0261_ ),
    .B1(\hash/_0323_ ),
    .Y(\hash/_0324_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3049_  (.A1(\hash/_1486_ ),
    .A2(\hash/_0247_ ),
    .A3(\hash/_0258_ ),
    .B1(\hash/_0324_ ),
    .Y(\hash/_0325_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3050_  (.A(\hash/_1514_ ),
    .B(\hash/_1516_ ),
    .C(\hash/_0306_ ),
    .Y(\hash/_0326_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3051_  (.A(\hash/_1510_ ),
    .B(\hash/_1512_ ),
    .C(\hash/_1514_ ),
    .D(\hash/_1516_ ),
    .Y(\hash/_0327_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3052_  (.A(\hash/_1514_ ),
    .B(\hash/_1516_ ),
    .Y(\hash/_0328_ ));
 sky130_fd_sc_hd__o32a_1 \hash/_3053_  (.A1(\hash/_0308_ ),
    .A2(\hash/_0310_ ),
    .A3(\hash/_0327_ ),
    .B1(\hash/_0328_ ),
    .B2(\hash/_0311_ ),
    .X(\hash/_0329_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3054_  (.A1(\hash/_1516_ ),
    .A2(\hash/_1513_ ),
    .B1(\hash/_1515_ ),
    .Y(\hash/_0330_ ));
 sky130_fd_sc_hd__o211a_2 \hash/_3055_  (.A1(\hash/_0325_ ),
    .A2(\hash/_0326_ ),
    .B1(\hash/_0329_ ),
    .C1(\hash/_0330_ ),
    .X(\hash/_0331_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3056_  (.A(\hash/_1518_ ),
    .B(\hash/_0331_ ),
    .Y(\hash/_0011_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3057_  (.A(\hash/_0330_ ),
    .Y(\hash/_0332_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3058_  (.A(\hash/_1514_ ),
    .B(\hash/_1516_ ),
    .C(\hash/_1518_ ),
    .X(\hash/_0333_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/_3059_  (.A1(\hash/_1518_ ),
    .A2(\hash/_0332_ ),
    .B1(\hash/_0333_ ),
    .B2(\hash/_0321_ ),
    .C1(\hash/_1517_ ),
    .Y(\hash/_0334_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3060_  (.A(\hash/_1520_ ),
    .B(\hash/_0334_ ),
    .Y(\hash/_0012_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3061_  (.A(\hash/_1522_ ),
    .Y(\hash/_0335_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3062_  (.A(\hash/_1518_ ),
    .B(\hash/_1520_ ),
    .Y(\hash/_0336_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3063_  (.A1(\hash/_1520_ ),
    .A2(\hash/_1517_ ),
    .B1(\hash/_1519_ ),
    .Y(\hash/_0337_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3064_  (.A1(\hash/_0331_ ),
    .A2(\hash/_0336_ ),
    .B1(\hash/_0337_ ),
    .Y(\hash/_0338_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3065_  (.A(\hash/_0335_ ),
    .B(\hash/_0338_ ),
    .Y(\hash/_0013_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3066_  (.A(\hash/_1516_ ),
    .B(\hash/_1518_ ),
    .C(\hash/_1520_ ),
    .X(\hash/_0339_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3067_  (.A1(\hash/_1518_ ),
    .A2(\hash/_1515_ ),
    .B1(\hash/_1517_ ),
    .X(\hash/_0340_ ));
 sky130_fd_sc_hd__a221o_1 \hash/_3068_  (.A1(\hash/_1520_ ),
    .A2(\hash/_0340_ ),
    .B1(\hash/_0339_ ),
    .B2(\hash/_1513_ ),
    .C1(\hash/_1519_ ),
    .X(\hash/_0341_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3069_  (.A1(\hash/_1514_ ),
    .A2(\hash/_0321_ ),
    .A3(\hash/_0339_ ),
    .B1(\hash/_0341_ ),
    .Y(\hash/_0342_ ));
 sky130_fd_sc_hd__o21ba_1 \hash/_3070_  (.A1(\hash/_0335_ ),
    .A2(\hash/_0342_ ),
    .B1_N(\hash/_1521_ ),
    .X(\hash/_0343_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3071_  (.A(\hash/_1524_ ),
    .B(\hash/_0343_ ),
    .Y(\hash/_0014_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3072_  (.A1(\hash/_1524_ ),
    .A2(\hash/_1521_ ),
    .B1(\hash/_1523_ ),
    .X(\hash/_0344_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3073_  (.A1(\hash/_1522_ ),
    .A2(\hash/_1524_ ),
    .A3(\hash/_0338_ ),
    .B1(\hash/_0344_ ),
    .Y(\hash/_0345_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3074_  (.A(\hash/_1526_ ),
    .B(\hash/_0345_ ),
    .Y(\hash/_0015_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3076_  (.A1(\hash/_1522_ ),
    .A2(\hash/_1519_ ),
    .B1(\hash/_1521_ ),
    .Y(\hash/_0347_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3077_  (.A(\hash/_0347_ ),
    .B_N(\hash/_1524_ ),
    .Y(\hash/_0348_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3078_  (.A1(\hash/_1523_ ),
    .A2(\hash/_0348_ ),
    .B1(\hash/_1526_ ),
    .Y(\hash/_0349_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3079_  (.A_N(\hash/_1525_ ),
    .B(\hash/_0349_ ),
    .Y(\hash/_0350_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3080_  (.A(\hash/_1520_ ),
    .B(\hash/_1522_ ),
    .C(\hash/_1524_ ),
    .D(\hash/_1526_ ),
    .Y(\hash/_0351_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3081_  (.A(\hash/_0334_ ),
    .B(\hash/_0351_ ),
    .Y(\hash/_0352_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3082_  (.A(\hash/_0350_ ),
    .B(\hash/_0352_ ),
    .Y(\hash/_0353_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3083_  (.A(\hash/_1528_ ),
    .B(\hash/_0353_ ),
    .Y(\hash/_0016_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3084_  (.A(\hash/_1522_ ),
    .B(\hash/_1524_ ),
    .C(\hash/_1526_ ),
    .D(\hash/_1528_ ),
    .Y(\hash/_0354_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3085_  (.A1(\hash/_1526_ ),
    .A2(\hash/_0344_ ),
    .B1(\hash/_1525_ ),
    .X(\hash/_0355_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3086_  (.A1(\hash/_1528_ ),
    .A2(\hash/_0355_ ),
    .B1(\hash/_1527_ ),
    .Y(\hash/_0356_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3087_  (.A1(\hash/_0337_ ),
    .A2(\hash/_0354_ ),
    .B1(\hash/_0356_ ),
    .X(\hash/_0357_ ));
 sky130_fd_sc_hd__o31a_1 \hash/_3088_  (.A1(\hash/_0331_ ),
    .A2(\hash/_0336_ ),
    .A3(\hash/_0354_ ),
    .B1(\hash/_0357_ ),
    .X(\hash/_0358_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3089_  (.A(\hash/_1530_ ),
    .B(\hash/_0358_ ),
    .Y(\hash/_0017_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3091_  (.A1(\hash/_0342_ ),
    .A2(\hash/_0354_ ),
    .B1(\hash/_0356_ ),
    .Y(\hash/_0360_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3092_  (.A1(\hash/_1530_ ),
    .A2(\hash/_0360_ ),
    .B1(\hash/_1529_ ),
    .Y(\hash/_0361_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3093_  (.A(\hash/_1532_ ),
    .B(\hash/_0361_ ),
    .Y(\hash/_0018_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3094_  (.A(\hash/_1526_ ),
    .B(\hash/_1528_ ),
    .C(\hash/_1530_ ),
    .D(\hash/_1532_ ),
    .Y(\hash/_0362_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3095_  (.A1(\hash/_1528_ ),
    .A2(\hash/_1525_ ),
    .B1(\hash/_1527_ ),
    .X(\hash/_0363_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3096_  (.A1(\hash/_1530_ ),
    .A2(\hash/_0363_ ),
    .B1(\hash/_1529_ ),
    .X(\hash/_0364_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3097_  (.A1(\hash/_1532_ ),
    .A2(\hash/_0364_ ),
    .B1(\hash/_1531_ ),
    .Y(\hash/_0365_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3098_  (.A1(\hash/_0345_ ),
    .A2(\hash/_0362_ ),
    .B1(\hash/_0365_ ),
    .Y(\hash/_0366_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3099_  (.A(\hash/_1534_ ),
    .B(\hash/_0366_ ),
    .X(\hash/_0019_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3100_  (.A(\hash/_1530_ ),
    .B(\hash/_1532_ ),
    .C(\hash/_1534_ ),
    .X(\hash/_0367_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3101_  (.A1(\hash/_1528_ ),
    .A2(\hash/_0350_ ),
    .B1(\hash/_1527_ ),
    .X(\hash/_0368_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3102_  (.A1(\hash/_1530_ ),
    .A2(\hash/_0368_ ),
    .B1(\hash/_1529_ ),
    .Y(\hash/_0369_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3103_  (.A(\hash/_1532_ ),
    .B(\hash/_1534_ ),
    .Y(\hash/_0370_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3104_  (.A1(\hash/_1534_ ),
    .A2(\hash/_1531_ ),
    .B1(\hash/_1533_ ),
    .Y(\hash/_0371_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3105_  (.A1(\hash/_0369_ ),
    .A2(\hash/_0370_ ),
    .B1(\hash/_0371_ ),
    .Y(\hash/_0372_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3106_  (.A1(\hash/_1528_ ),
    .A2(\hash/_0352_ ),
    .A3(\hash/_0367_ ),
    .B1(\hash/_0372_ ),
    .Y(\hash/_0373_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3107_  (.A(\hash/_1536_ ),
    .B(\hash/_0373_ ),
    .Y(\hash/_0021_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_3110_  (.A0(\hash/a_new[31] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/a[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3111_  (.A(_09578_),
    .B(\hash/a_new[31] ),
    .Y(\hash/_0376_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3112_  (.A(reset_hash_dash),
    .B(\hash/_0376_ ),
    .Y(\hash/_0377_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3113_  (.A(\hash/_1530_ ),
    .B(\hash/_1532_ ),
    .C(\hash/_1534_ ),
    .Y(\hash/_0378_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3114_  (.A1(\hash/_1532_ ),
    .A2(\hash/_1529_ ),
    .B1(\hash/_1531_ ),
    .X(\hash/_0379_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3115_  (.A1(\hash/_1534_ ),
    .A2(\hash/_0379_ ),
    .B1(\hash/_1533_ ),
    .Y(\hash/_0380_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3116_  (.A1(\hash/_0358_ ),
    .A2(\hash/_0378_ ),
    .B1(\hash/_0380_ ),
    .Y(\hash/_0381_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3117_  (.A1(\hash/_1536_ ),
    .A2(\hash/_0381_ ),
    .B1(\hash/_1535_ ),
    .Y(\hash/_0382_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3118_  (.A(\hash/_0377_ ),
    .B(\hash/_0382_ ),
    .Y(\hash/_0022_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3119_  (.A(\hash/_1464_ ),
    .B(\hash/_1542_ ),
    .X(\hash/_0050_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3120_  (.A1(\hash/_1463_ ),
    .A2(\hash/_1538_ ),
    .B1(\hash/_1537_ ),
    .C1(\hash/_1541_ ),
    .Y(\hash/_0383_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3121_  (.A1(\hash/_1542_ ),
    .A2(\hash/_1541_ ),
    .B1(\hash/_1540_ ),
    .Y(\hash/_0384_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3122_  (.A(\hash/_0383_ ),
    .B(\hash/_0384_ ),
    .Y(\hash/_0385_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3123_  (.A1(\hash/_1463_ ),
    .A2(\hash/_1538_ ),
    .B1(\hash/_1537_ ),
    .X(\hash/_0386_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3124_  (.A1(\hash/_1542_ ),
    .A2(\hash/_0386_ ),
    .B1(\hash/_1541_ ),
    .C1(\hash/_1540_ ),
    .Y(\hash/_0387_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3125_  (.A(\hash/_0385_ ),
    .B(\hash/_0387_ ),
    .Y(\hash/_0053_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3126_  (.A1(\hash/_1464_ ),
    .A2(\hash/_1542_ ),
    .B1(\hash/_1541_ ),
    .X(\hash/_0388_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3127_  (.A1(\hash/_1540_ ),
    .A2(\hash/_0388_ ),
    .B1(\hash/_1539_ ),
    .Y(\hash/_0389_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3128_  (.A(\hash/_1544_ ),
    .B(\hash/_0389_ ),
    .Y(\hash/_0054_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3129_  (.A(\hash/_1544_ ),
    .Y(\hash/_0390_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3130_  (.A(\hash/_1539_ ),
    .B(\hash/_0385_ ),
    .Y(\hash/_0391_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3131_  (.A(\hash/_0390_ ),
    .B(\hash/_0391_ ),
    .Y(\hash/_0392_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3132_  (.A(\hash/_1543_ ),
    .B(\hash/_0392_ ),
    .Y(\hash/_0393_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3133_  (.A(\hash/_1546_ ),
    .B(\hash/_0393_ ),
    .Y(\hash/_0055_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3134_  (.A1(\hash/_0390_ ),
    .A2(\hash/_0389_ ),
    .B1_N(\hash/_1543_ ),
    .Y(\hash/_0394_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3135_  (.A1(\hash/_1546_ ),
    .A2(\hash/_0394_ ),
    .B1(\hash/_1545_ ),
    .Y(\hash/_0395_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3136_  (.A(\hash/_1548_ ),
    .B(\hash/_0395_ ),
    .Y(\hash/_0056_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3137_  (.A1(\hash/_1548_ ),
    .A2(\hash/_1545_ ),
    .B1(\hash/_1547_ ),
    .Y(\hash/_0396_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3138_  (.A(\hash/_1539_ ),
    .B(\hash/_1543_ ),
    .Y(\hash/_0397_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3139_  (.A(\hash/_0396_ ),
    .B(\hash/_0397_ ),
    .Y(\hash/_0398_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3140_  (.A(\hash/_1544_ ),
    .B(\hash/_1543_ ),
    .Y(\hash/_0399_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3141_  (.A(\hash/_1546_ ),
    .B(\hash/_1548_ ),
    .Y(\hash/_0400_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3142_  (.A1(\hash/_0399_ ),
    .A2(\hash/_0400_ ),
    .B1(\hash/_0396_ ),
    .Y(\hash/_0401_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3143_  (.A1(\hash/_0385_ ),
    .A2(\hash/_0398_ ),
    .B1(\hash/_0401_ ),
    .Y(\hash/_0402_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3144_  (.A(\hash/_1550_ ),
    .B(\hash/_0402_ ),
    .Y(\hash/_0057_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3145_  (.A(\hash/_1548_ ),
    .Y(\hash/_0403_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3146_  (.A1(\hash/_0403_ ),
    .A2(\hash/_0395_ ),
    .B1_N(\hash/_1547_ ),
    .Y(\hash/_0404_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3147_  (.A1(\hash/_1550_ ),
    .A2(\hash/_0404_ ),
    .B1(\hash/_1549_ ),
    .Y(\hash/_0405_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3148_  (.A(\hash/_1552_ ),
    .B(\hash/_0405_ ),
    .Y(\hash/_0058_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3149_  (.A(\hash/_1550_ ),
    .Y(\hash/_0406_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3150_  (.A(\hash/_1549_ ),
    .Y(\hash/_0407_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3151_  (.A1(\hash/_0406_ ),
    .A2(\hash/_0402_ ),
    .B1(\hash/_0407_ ),
    .Y(\hash/_0408_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3152_  (.A1(\hash/_1552_ ),
    .A2(\hash/_0408_ ),
    .B1(\hash/_1551_ ),
    .Y(\hash/_0409_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3153_  (.A(\hash/_1554_ ),
    .B(\hash/_0409_ ),
    .Y(\hash/_0059_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3154_  (.A(\hash/_1552_ ),
    .Y(\hash/_0410_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3155_  (.A1(\hash/_0410_ ),
    .A2(\hash/_0405_ ),
    .B1_N(\hash/_1551_ ),
    .Y(\hash/_0411_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3156_  (.A1(\hash/_1554_ ),
    .A2(\hash/_0411_ ),
    .B1(\hash/_1553_ ),
    .Y(\hash/_0412_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3157_  (.A(\hash/_1556_ ),
    .B(\hash/_0412_ ),
    .Y(\hash/_0030_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3158_  (.A1(\hash/_1554_ ),
    .A2(\hash/_1551_ ),
    .B1(\hash/_1553_ ),
    .X(\hash/_0413_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3159_  (.A1(\hash/_1556_ ),
    .A2(\hash/_0413_ ),
    .B1(\hash/_1555_ ),
    .Y(\hash/_0414_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3160_  (.A(\hash/_1554_ ),
    .B(\hash/_1556_ ),
    .C(\hash/_1552_ ),
    .Y(\hash/_0415_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3161_  (.A(\hash/_1550_ ),
    .B(\hash/_1549_ ),
    .Y(\hash/_0416_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3162_  (.A1(\hash/_0415_ ),
    .A2(\hash/_0416_ ),
    .B1(\hash/_0414_ ),
    .X(\hash/_0417_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3163_  (.A1(\hash/_0407_ ),
    .A2(\hash/_0402_ ),
    .A3(\hash/_0414_ ),
    .B1(\hash/_0417_ ),
    .Y(\hash/_0418_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3164_  (.A(\hash/_1558_ ),
    .B(\hash/_0418_ ),
    .X(\hash/_0031_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3165_  (.A1(\hash/_1550_ ),
    .A2(\hash/_1547_ ),
    .B1(\hash/_1549_ ),
    .Y(\hash/_0419_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3166_  (.A1(\hash/_0415_ ),
    .A2(\hash/_0419_ ),
    .B1(\hash/_0414_ ),
    .Y(\hash/_0420_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3167_  (.A(\hash/_0390_ ),
    .B(\hash/_0389_ ),
    .Y(\hash/_0421_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3168_  (.A(\hash/_1554_ ),
    .B(\hash/_1556_ ),
    .C(\hash/_1550_ ),
    .D(\hash/_1552_ ),
    .Y(\hash/_0422_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3169_  (.A(\hash/_0400_ ),
    .B(\hash/_0422_ ),
    .Y(\hash/_0423_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3170_  (.A(\hash/_1548_ ),
    .B(\hash/_1545_ ),
    .Y(\hash/_0424_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3171_  (.A(\hash/_1546_ ),
    .B(\hash/_1548_ ),
    .C(\hash/_1543_ ),
    .Y(\hash/_0425_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3172_  (.A1(\hash/_0424_ ),
    .A2(\hash/_0425_ ),
    .B1(\hash/_0422_ ),
    .Y(\hash/_0426_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3173_  (.A1(\hash/_0421_ ),
    .A2(\hash/_0423_ ),
    .B1(\hash/_0426_ ),
    .Y(\hash/_0427_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3174_  (.A_N(\hash/_0420_ ),
    .B(\hash/_0427_ ),
    .Y(\hash/_0428_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3175_  (.A1(\hash/_1558_ ),
    .A2(\hash/_0428_ ),
    .B1(\hash/_1557_ ),
    .Y(\hash/_0429_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3176_  (.A(\hash/_1560_ ),
    .B(\hash/_0429_ ),
    .Y(\hash/_0032_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3177_  (.A1(\hash/_1560_ ),
    .A2(\hash/_1557_ ),
    .B1(\hash/_1559_ ),
    .X(\hash/_0430_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3178_  (.A(\hash/_1558_ ),
    .B(\hash/_1560_ ),
    .Y(\hash/_0431_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/_3179_  (.A1(\hash/_0407_ ),
    .A2(\hash/_0402_ ),
    .A3(\hash/_0414_ ),
    .B1(\hash/_0417_ ),
    .C1(\hash/_0431_ ),
    .Y(\hash/_0432_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3180_  (.A1(\hash/_0430_ ),
    .A2(\hash/_0432_ ),
    .B1(\hash/_1562_ ),
    .X(\hash/_0433_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3181_  (.A(\hash/_1562_ ),
    .B(\hash/_0430_ ),
    .C(\hash/_0432_ ),
    .Y(\hash/_0434_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3182_  (.A(\hash/_0433_ ),
    .B(\hash/_0434_ ),
    .Y(\hash/_0033_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3184_  (.A(\hash/_1562_ ),
    .Y(\hash/_0436_ ));
 sky130_fd_sc_hd__or2_2 \hash/_3185_  (.A(\hash/_1557_ ),
    .B(\hash/_1559_ ),
    .X(\hash/_0437_ ));
 sky130_fd_sc_hd__a2111oi_2 \hash/_3186_  (.A1(\hash/_0421_ ),
    .A2(\hash/_0423_ ),
    .B1(\hash/_0426_ ),
    .C1(\hash/_0437_ ),
    .D1(\hash/_0420_ ),
    .Y(\hash/_0438_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3187_  (.A(\hash/_1558_ ),
    .B(\hash/_1557_ ),
    .C(\hash/_1559_ ),
    .Y(\hash/_0439_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3188_  (.A(\hash/_1560_ ),
    .B(\hash/_1559_ ),
    .Y(\hash/_0440_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3189_  (.A(\hash/_1561_ ),
    .Y(\hash/_0441_ ));
 sky130_fd_sc_hd__o41ai_2 \hash/_3190_  (.A1(\hash/_0436_ ),
    .A2(\hash/_0438_ ),
    .A3(\hash/_0439_ ),
    .A4(\hash/_0440_ ),
    .B1(\hash/_0441_ ),
    .Y(\hash/_0442_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3191_  (.A(\hash/_1564_ ),
    .B(\hash/_0442_ ),
    .X(\hash/_0034_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3192_  (.A1(\hash/_1561_ ),
    .A2(\hash/_0433_ ),
    .B1(\hash/_1564_ ),
    .X(\hash/_0443_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3193_  (.A(\hash/_1563_ ),
    .B(\hash/_0443_ ),
    .Y(\hash/_0444_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3194_  (.A(\hash/_1568_ ),
    .B(\hash/_0444_ ),
    .Y(\hash/_0035_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3195_  (.A1(\hash/_1564_ ),
    .A2(\hash/_0442_ ),
    .B1(\hash/_1563_ ),
    .X(\hash/_0445_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3196_  (.A1(\hash/_1568_ ),
    .A2(\hash/_0445_ ),
    .B1(\hash/_1567_ ),
    .Y(\hash/_0446_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3197_  (.A(\hash/_1566_ ),
    .B(\hash/_0446_ ),
    .Y(\hash/_0036_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3198_  (.A1(\hash/_1568_ ),
    .A2(\hash/_1563_ ),
    .B1(\hash/_1567_ ),
    .X(\hash/_0447_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_3199_  (.A1(\hash/_1561_ ),
    .A2(\hash/_0433_ ),
    .B1(\hash/_1564_ ),
    .C1(\hash/_1568_ ),
    .Y(\hash/_0448_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3200_  (.A_N(\hash/_0447_ ),
    .B(\hash/_0448_ ),
    .Y(\hash/_0449_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3201_  (.A1(\hash/_1566_ ),
    .A2(\hash/_0449_ ),
    .B1(\hash/_1565_ ),
    .Y(\hash/_0450_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3202_  (.A(\hash/_1570_ ),
    .B(\hash/_0450_ ),
    .Y(\hash/_0037_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3203_  (.A(\hash/_1568_ ),
    .B(\hash/_1566_ ),
    .C(\hash/_1570_ ),
    .X(\hash/_0451_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3204_  (.A(\hash/_1570_ ),
    .Y(\hash/_0452_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3205_  (.A1(\hash/_1566_ ),
    .A2(\hash/_0447_ ),
    .B1(\hash/_1565_ ),
    .Y(\hash/_0453_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3206_  (.A(\hash/_0452_ ),
    .B(\hash/_0453_ ),
    .Y(\hash/_0454_ ));
 sky130_fd_sc_hd__a311o_1 \hash/_3207_  (.A1(\hash/_1564_ ),
    .A2(\hash/_0442_ ),
    .A3(\hash/_0451_ ),
    .B1(\hash/_0454_ ),
    .C1(\hash/_1569_ ),
    .X(\hash/_0455_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3208_  (.A(\hash/_1572_ ),
    .B(\hash/_0455_ ),
    .X(\hash/_0038_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3209_  (.A1(\hash/_1564_ ),
    .A2(\hash/_1561_ ),
    .B1(\hash/_1563_ ),
    .X(\hash/_0456_ ));
 sky130_fd_sc_hd__a31o_1 \hash/_3210_  (.A1(\hash/_1562_ ),
    .A2(\hash/_1564_ ),
    .A3(\hash/_0430_ ),
    .B1(\hash/_0456_ ),
    .X(\hash/_0457_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3211_  (.A(\hash/_1566_ ),
    .B(\hash/_1570_ ),
    .C(\hash/_1567_ ),
    .Y(\hash/_0458_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3212_  (.A1(\hash/_1570_ ),
    .A2(\hash/_1565_ ),
    .B1(\hash/_1569_ ),
    .Y(\hash/_0459_ ));
 sky130_fd_sc_hd__a21boi_0 \hash/_3213_  (.A1(\hash/_0458_ ),
    .A2(\hash/_0459_ ),
    .B1_N(\hash/_1572_ ),
    .Y(\hash/_0460_ ));
 sky130_fd_sc_hd__a311o_1 \hash/_3214_  (.A1(\hash/_1572_ ),
    .A2(\hash/_0451_ ),
    .A3(\hash/_0457_ ),
    .B1(\hash/_0460_ ),
    .C1(\hash/_1571_ ),
    .X(\hash/_0461_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3215_  (.A(\hash/_1564_ ),
    .B(\hash/_1572_ ),
    .C(\hash/_0451_ ),
    .X(\hash/_0462_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3216_  (.A(\hash/_1558_ ),
    .B(\hash/_1560_ ),
    .C(\hash/_1562_ ),
    .D(\hash/_0462_ ),
    .Y(\hash/_0463_ ));
 sky130_fd_sc_hd__a311o_1 \hash/_3217_  (.A1(\hash/_0407_ ),
    .A2(\hash/_0402_ ),
    .A3(\hash/_0414_ ),
    .B1(\hash/_0417_ ),
    .C1(\hash/_0463_ ),
    .X(\hash/_0464_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3218_  (.A(\hash/_0461_ ),
    .B_N(\hash/_0464_ ),
    .Y(\hash/_0465_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3219_  (.A(\hash/_1574_ ),
    .B(\hash/_0465_ ),
    .Y(\hash/_0039_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3220_  (.A1(\hash/_1572_ ),
    .A2(\hash/_0455_ ),
    .B1(\hash/_1571_ ),
    .X(\hash/_0466_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3221_  (.A1(\hash/_1574_ ),
    .A2(\hash/_0466_ ),
    .B1(\hash/_1573_ ),
    .Y(\hash/_0467_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3222_  (.A(\hash/_1576_ ),
    .B(\hash/_0467_ ),
    .Y(\hash/_0040_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3223_  (.A(\hash/_1573_ ),
    .B(\hash/_1575_ ),
    .C(\hash/_0461_ ),
    .Y(\hash/_0468_ ));
 sky130_fd_sc_hd__or2_2 \hash/_3224_  (.A(\hash/_1574_ ),
    .B(\hash/_1573_ ),
    .X(\hash/_0469_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3225_  (.A1(\hash/_1576_ ),
    .A2(\hash/_0469_ ),
    .B1(\hash/_1575_ ),
    .Y(\hash/_0470_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3226_  (.A1(\hash/_0464_ ),
    .A2(\hash/_0468_ ),
    .B1(\hash/_0470_ ),
    .Y(\hash/_0471_ ));
 sky130_fd_sc_hd__and2_1 \hash/_3227_  (.A(\hash/_1578_ ),
    .B(\hash/_0471_ ),
    .X(\hash/_0472_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3228_  (.A(\hash/_1578_ ),
    .B(\hash/_0471_ ),
    .Y(\hash/_0473_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3229_  (.A(\hash/_0472_ ),
    .B(\hash/_0473_ ),
    .Y(\hash/_0041_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3230_  (.A(\hash/_1574_ ),
    .B(\hash/_1576_ ),
    .C(\hash/_1578_ ),
    .X(\hash/_0474_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3231_  (.A(\hash/_1569_ ),
    .B(\hash/_1571_ ),
    .C(\hash/_1573_ ),
    .Y(\hash/_0475_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3232_  (.A1(\hash/_0452_ ),
    .A2(\hash/_0453_ ),
    .B1(\hash/_0475_ ),
    .Y(\hash/_0476_ ));
 sky130_fd_sc_hd__or3_1 \hash/_3233_  (.A(\hash/_1572_ ),
    .B(\hash/_1571_ ),
    .C(\hash/_1573_ ),
    .X(\hash/_0477_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_3234_  (.A1(\hash/_1576_ ),
    .A2(\hash/_0469_ ),
    .A3(\hash/_0476_ ),
    .A4(\hash/_0477_ ),
    .B1(\hash/_1575_ ),
    .Y(\hash/_0478_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3235_  (.A(\hash/_0478_ ),
    .B_N(\hash/_1578_ ),
    .Y(\hash/_0479_ ));
 sky130_fd_sc_hd__a311oi_2 \hash/_3236_  (.A1(\hash/_0442_ ),
    .A2(\hash/_0462_ ),
    .A3(\hash/_0474_ ),
    .B1(\hash/_0479_ ),
    .C1(\hash/_1577_ ),
    .Y(\hash/_0480_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3237_  (.A(\hash/_1580_ ),
    .B(\hash/_0480_ ),
    .Y(\hash/_0042_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3238_  (.A1(\hash/_1577_ ),
    .A2(\hash/_0472_ ),
    .B1(\hash/_1580_ ),
    .X(\hash/_0481_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3239_  (.A(\hash/_1579_ ),
    .B(\hash/_0481_ ),
    .Y(\hash/_0482_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3240_  (.A(\hash/_1582_ ),
    .B(\hash/_0482_ ),
    .Y(\hash/_0043_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3241_  (.A(\hash/_1584_ ),
    .Y(\hash/_0483_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3242_  (.A(\hash/_1580_ ),
    .B(\hash/_1582_ ),
    .Y(\hash/_0484_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3243_  (.A1(\hash/_1582_ ),
    .A2(\hash/_1579_ ),
    .B1(\hash/_1581_ ),
    .Y(\hash/_0485_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3244_  (.A1(\hash/_0480_ ),
    .A2(\hash/_0484_ ),
    .B1(\hash/_0485_ ),
    .Y(\hash/_0486_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3245_  (.A(\hash/_0483_ ),
    .B(\hash/_0486_ ),
    .Y(\hash/_0044_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3246_  (.A1(\hash/_1584_ ),
    .A2(\hash/_1581_ ),
    .B1(\hash/_1583_ ),
    .X(\hash/_0487_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3247_  (.A(\hash/_1582_ ),
    .B(\hash/_1579_ ),
    .Y(\hash/_0488_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3248_  (.A(\hash/_1580_ ),
    .B(\hash/_1582_ ),
    .C(\hash/_1577_ ),
    .Y(\hash/_0489_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3249_  (.A(\hash/_0488_ ),
    .B(\hash/_0489_ ),
    .Y(\hash/_0490_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_3250_  (.A1(\hash/_1578_ ),
    .A2(\hash/_1580_ ),
    .A3(\hash/_1582_ ),
    .A4(\hash/_0471_ ),
    .B1(\hash/_0490_ ),
    .Y(\hash/_0491_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3251_  (.A(\hash/_0483_ ),
    .B(\hash/_0491_ ),
    .Y(\hash/_0492_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3252_  (.A(\hash/_0487_ ),
    .B(\hash/_0492_ ),
    .Y(\hash/_0493_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3253_  (.A(\hash/_1586_ ),
    .B(\hash/_0493_ ),
    .Y(\hash/_0045_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3254_  (.A(\hash/_0480_ ),
    .B(\hash/_0484_ ),
    .Y(\hash/_0494_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3255_  (.A(\hash/_0483_ ),
    .B(\hash/_0485_ ),
    .Y(\hash/_0495_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3256_  (.A1(\hash/_1583_ ),
    .A2(\hash/_0495_ ),
    .B1(\hash/_1586_ ),
    .Y(\hash/_0496_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3257_  (.A_N(\hash/_1585_ ),
    .B(\hash/_0496_ ),
    .Y(\hash/_0497_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3258_  (.A1(\hash/_1584_ ),
    .A2(\hash/_1586_ ),
    .A3(\hash/_0494_ ),
    .B1(\hash/_0497_ ),
    .Y(\hash/_0498_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3259_  (.A(\hash/_1588_ ),
    .B(\hash/_0498_ ),
    .Y(\hash/_0046_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3260_  (.A(\hash/_1584_ ),
    .B(\hash/_1586_ ),
    .C(\hash/_1588_ ),
    .Y(\hash/_0499_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3261_  (.A1(\hash/_1586_ ),
    .A2(\hash/_0487_ ),
    .B1(\hash/_1585_ ),
    .X(\hash/_0500_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3262_  (.A1(\hash/_1588_ ),
    .A2(\hash/_0500_ ),
    .B1(\hash/_1587_ ),
    .X(\hash/_0501_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3263_  (.A1(\hash/_0491_ ),
    .A2(\hash/_0499_ ),
    .B1_N(\hash/_0501_ ),
    .Y(\hash/_0502_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3264_  (.A(\hash/_1590_ ),
    .B(\hash/_0502_ ),
    .X(\hash/_0047_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3265_  (.A1(\hash/_1586_ ),
    .A2(\hash/_1583_ ),
    .B1(\hash/_1585_ ),
    .X(\hash/_0503_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3266_  (.A1(\hash/_1588_ ),
    .A2(\hash/_0503_ ),
    .B1(\hash/_1589_ ),
    .C1(\hash/_1587_ ),
    .Y(\hash/_0504_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3267_  (.A(\hash/_0485_ ),
    .B(\hash/_0504_ ),
    .Y(\hash/_0505_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3268_  (.A(\hash/_1590_ ),
    .B(\hash/_1589_ ),
    .Y(\hash/_0506_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3269_  (.A1(\hash/_0499_ ),
    .A2(\hash/_0504_ ),
    .B1(\hash/_0506_ ),
    .Y(\hash/_0507_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3270_  (.A1(\hash/_0494_ ),
    .A2(\hash/_0505_ ),
    .B1(\hash/_0507_ ),
    .Y(\hash/_0508_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3271_  (.A(\hash/_1592_ ),
    .B(\hash/_0508_ ),
    .Y(\hash/_0048_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3272_  (.A(\hash/_1584_ ),
    .B(\hash/_1586_ ),
    .C(\hash/_1588_ ),
    .X(\hash/_0509_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3273_  (.A(\hash/_1590_ ),
    .B(\hash/_1592_ ),
    .C(\hash/_0509_ ),
    .Y(\hash/_0510_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3274_  (.A1(\hash/_1590_ ),
    .A2(\hash/_0501_ ),
    .B1(\hash/_1589_ ),
    .X(\hash/_0511_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3275_  (.A1(\hash/_1592_ ),
    .A2(\hash/_0511_ ),
    .B1(\hash/_1591_ ),
    .Y(\hash/_0512_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3276_  (.A1(\hash/_0491_ ),
    .A2(\hash/_0510_ ),
    .B1(\hash/_0512_ ),
    .Y(\hash/_0513_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3277_  (.A(\hash/_1594_ ),
    .B(\hash/_0513_ ),
    .X(\hash/_0049_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3278_  (.A(\hash/_1590_ ),
    .B(\hash/_1592_ ),
    .C(\hash/_0509_ ),
    .X(\hash/_0514_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3279_  (.A1(\hash/_1592_ ),
    .A2(\hash/_1589_ ),
    .B1(\hash/_1591_ ),
    .C1(\hash/_1587_ ),
    .Y(\hash/_0515_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3280_  (.A(\hash/_1588_ ),
    .B(\hash/_0497_ ),
    .Y(\hash/_0516_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3281_  (.A(\hash/_0506_ ),
    .B_N(\hash/_1592_ ),
    .Y(\hash/_0517_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3282_  (.A1(\hash/_1591_ ),
    .A2(\hash/_0517_ ),
    .B1(\hash/_1594_ ),
    .Y(\hash/_0518_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3283_  (.A1(\hash/_0515_ ),
    .A2(\hash/_0516_ ),
    .B1(\hash/_0518_ ),
    .Y(\hash/_0519_ ));
 sky130_fd_sc_hd__a311oi_1 \hash/_3284_  (.A1(\hash/_1594_ ),
    .A2(\hash/_0494_ ),
    .A3(\hash/_0514_ ),
    .B1(\hash/_0519_ ),
    .C1(\hash/_1593_ ),
    .Y(\hash/_0520_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3285_  (.A(\hash/_1596_ ),
    .B(\hash/_0520_ ),
    .Y(\hash/_0051_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_3286_  (.A0(\hash/b_new[31] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/b[31] ));
 sky130_fd_sc_hd__nand2_1 \hash/_3287_  (.A(\hash/_1594_ ),
    .B(\hash/_1596_ ),
    .Y(\hash/_0521_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3288_  (.A(\hash/_0512_ ),
    .B(\hash/_0521_ ),
    .Y(\hash/_0522_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3289_  (.A1(\hash/_1596_ ),
    .A2(\hash/_1593_ ),
    .B1(\hash/_1595_ ),
    .C1(\hash/_0522_ ),
    .Y(\hash/_0523_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_3290_  (.A1(\hash/_0491_ ),
    .A2(\hash/_0510_ ),
    .A3(\hash/_0521_ ),
    .B1(\hash/_0523_ ),
    .Y(\hash/_0524_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3291_  (.A(_09577_),
    .B(\hash/b_new[31] ),
    .Y(\hash/_0525_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3292_  (.A(reset_hash_dash),
    .B(\hash/_0525_ ),
    .Y(\hash/_0526_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3293_  (.A(\hash/_0524_ ),
    .B(\hash/_0526_ ),
    .X(\hash/_0052_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3294_  (.A(\hash/_1466_ ),
    .B(\hash/_1602_ ),
    .X(\hash/_0080_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3295_  (.A1(\hash/_1465_ ),
    .A2(\hash/_1598_ ),
    .B1(\hash/_1597_ ),
    .X(\hash/_0527_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3296_  (.A1(\hash/_1602_ ),
    .A2(\hash/_0527_ ),
    .B1(\hash/_1601_ ),
    .Y(\hash/_0528_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3297_  (.A(\hash/_1600_ ),
    .B(\hash/_0528_ ),
    .Y(\hash/_0083_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3298_  (.A1(\hash/_1466_ ),
    .A2(\hash/_1602_ ),
    .B1(\hash/_1601_ ),
    .X(\hash/_0529_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3299_  (.A1(\hash/_1600_ ),
    .A2(\hash/_0529_ ),
    .B1(\hash/_1599_ ),
    .Y(\hash/_0530_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3300_  (.A(\hash/_1604_ ),
    .B(\hash/_0530_ ),
    .Y(\hash/_0084_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3301_  (.A(\hash/_1600_ ),
    .Y(\hash/_0531_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3302_  (.A1(\hash/_0531_ ),
    .A2(\hash/_0528_ ),
    .B1_N(\hash/_1599_ ),
    .Y(\hash/_0532_ ));
 sky130_fd_sc_hd__and2_1 \hash/_3303_  (.A(\hash/_1604_ ),
    .B(\hash/_0532_ ),
    .X(\hash/_0533_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3304_  (.A(\hash/_1603_ ),
    .B(\hash/_0533_ ),
    .Y(\hash/_0534_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3305_  (.A(\hash/_1606_ ),
    .B(\hash/_0534_ ),
    .Y(\hash/_0085_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3306_  (.A(\hash/_1604_ ),
    .Y(\hash/_0535_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3307_  (.A1(\hash/_0535_ ),
    .A2(\hash/_0530_ ),
    .B1_N(\hash/_1603_ ),
    .Y(\hash/_0536_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3308_  (.A1(\hash/_1606_ ),
    .A2(\hash/_0536_ ),
    .B1(\hash/_1605_ ),
    .Y(\hash/_0537_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3309_  (.A(\hash/_1608_ ),
    .B(\hash/_0537_ ),
    .Y(\hash/_0086_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3310_  (.A1(\hash/_1603_ ),
    .A2(\hash/_0533_ ),
    .B1(\hash/_1606_ ),
    .Y(\hash/_0538_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3311_  (.A_N(\hash/_1605_ ),
    .B(\hash/_0538_ ),
    .Y(\hash/_0539_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3312_  (.A1(\hash/_1608_ ),
    .A2(\hash/_0539_ ),
    .B1(\hash/_1607_ ),
    .Y(\hash/_0540_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3313_  (.A(\hash/_1610_ ),
    .B(\hash/_0540_ ),
    .Y(\hash/_0087_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3314_  (.A(\hash/_1608_ ),
    .Y(\hash/_0541_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3315_  (.A1(\hash/_0541_ ),
    .A2(\hash/_0537_ ),
    .B1_N(\hash/_1607_ ),
    .Y(\hash/_0542_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3316_  (.A1(\hash/_1610_ ),
    .A2(\hash/_0542_ ),
    .B1(\hash/_1609_ ),
    .Y(\hash/_0543_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3317_  (.A(\hash/_1612_ ),
    .B(\hash/_0543_ ),
    .Y(\hash/_0088_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3318_  (.A(\hash/_1608_ ),
    .B(\hash/_1610_ ),
    .C(\hash/_1612_ ),
    .X(\hash/_0544_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3319_  (.A(\hash/_1612_ ),
    .Y(\hash/_0545_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3320_  (.A1(\hash/_1608_ ),
    .A2(\hash/_1605_ ),
    .B1(\hash/_1607_ ),
    .X(\hash/_0546_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3321_  (.A1(\hash/_1610_ ),
    .A2(\hash/_0546_ ),
    .B1(\hash/_1609_ ),
    .Y(\hash/_0547_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3322_  (.A1(\hash/_1606_ ),
    .A2(\hash/_1603_ ),
    .A3(\hash/_0544_ ),
    .B1(\hash/_1611_ ),
    .Y(\hash/_0548_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3323_  (.A1(\hash/_0545_ ),
    .A2(\hash/_0547_ ),
    .B1(\hash/_0548_ ),
    .Y(\hash/_0549_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_3324_  (.A1(\hash/_1604_ ),
    .A2(\hash/_1606_ ),
    .A3(\hash/_0532_ ),
    .A4(\hash/_0544_ ),
    .B1(\hash/_0549_ ),
    .Y(\hash/_0550_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3325_  (.A(\hash/_1614_ ),
    .B(\hash/_0550_ ),
    .Y(\hash/_0089_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3326_  (.A1(\hash/_0545_ ),
    .A2(\hash/_0543_ ),
    .B1_N(\hash/_1611_ ),
    .Y(\hash/_0551_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3327_  (.A1(\hash/_1614_ ),
    .A2(\hash/_0551_ ),
    .B1(\hash/_1613_ ),
    .Y(\hash/_0552_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3328_  (.A(\hash/_1616_ ),
    .B(\hash/_0552_ ),
    .Y(\hash/_0060_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3329_  (.A(\hash/_1614_ ),
    .B(\hash/_1616_ ),
    .Y(\hash/_0553_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3330_  (.A1(\hash/_1616_ ),
    .A2(\hash/_1613_ ),
    .B1(\hash/_1615_ ),
    .Y(\hash/_0554_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3331_  (.A1(\hash/_0550_ ),
    .A2(\hash/_0553_ ),
    .B1(\hash/_0554_ ),
    .Y(\hash/_0555_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3332_  (.A(\hash/_1618_ ),
    .B(\hash/_0555_ ),
    .X(\hash/_0061_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3333_  (.A(\hash/_1603_ ),
    .B(\hash/_1605_ ),
    .Y(\hash/_0556_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3334_  (.A1(\hash/_0535_ ),
    .A2(\hash/_0530_ ),
    .B1(\hash/_0556_ ),
    .Y(\hash/_0557_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3335_  (.A(\hash/_1606_ ),
    .B(\hash/_1605_ ),
    .Y(\hash/_0558_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3336_  (.A(\hash/_0553_ ),
    .B(\hash/_0558_ ),
    .Y(\hash/_0559_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3337_  (.A1(\hash/_1610_ ),
    .A2(\hash/_1607_ ),
    .B1(\hash/_1609_ ),
    .X(\hash/_0560_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3338_  (.A1(\hash/_1612_ ),
    .A2(\hash/_0560_ ),
    .B1(\hash/_1611_ ),
    .Y(\hash/_0561_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3339_  (.A1(\hash/_0553_ ),
    .A2(\hash/_0561_ ),
    .B1(\hash/_0554_ ),
    .Y(\hash/_0562_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3340_  (.A1(\hash/_0544_ ),
    .A2(\hash/_0557_ ),
    .A3(\hash/_0559_ ),
    .B1(\hash/_0562_ ),
    .Y(\hash/_0563_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3341_  (.A(\hash/_0563_ ),
    .B_N(\hash/_1618_ ),
    .Y(\hash/_0564_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3342_  (.A(\hash/_1617_ ),
    .B(\hash/_0564_ ),
    .Y(\hash/_0565_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3343_  (.A(\hash/_1620_ ),
    .B(\hash/_0565_ ),
    .Y(\hash/_0062_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3345_  (.A1(\hash/_1620_ ),
    .A2(\hash/_1617_ ),
    .B1(\hash/_1619_ ),
    .Y(\hash/_0567_ ));
 sky130_fd_sc_hd__and2_1 \hash/_3346_  (.A(\hash/_0554_ ),
    .B(\hash/_0567_ ),
    .X(\hash/_0568_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3347_  (.A(\hash/_1618_ ),
    .B(\hash/_1620_ ),
    .Y(\hash/_0569_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3348_  (.A1(\hash/_0554_ ),
    .A2(\hash/_0553_ ),
    .B1(\hash/_0569_ ),
    .Y(\hash/_0570_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3349_  (.A(\hash/_0570_ ),
    .B_N(\hash/_0567_ ),
    .Y(\hash/_0571_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3350_  (.A1(\hash/_0550_ ),
    .A2(\hash/_0568_ ),
    .B1(\hash/_0571_ ),
    .Y(\hash/_0572_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3351_  (.A(\hash/_1622_ ),
    .B(\hash/_0572_ ),
    .X(\hash/_0063_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3353_  (.A(\hash/_1618_ ),
    .B(\hash/_1620_ ),
    .C(\hash/_1622_ ),
    .Y(\hash/_0574_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3354_  (.A1(\hash/_1622_ ),
    .A2(\hash/_1619_ ),
    .B1(\hash/_1621_ ),
    .X(\hash/_0575_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3355_  (.A1(\hash/_1620_ ),
    .A2(\hash/_1622_ ),
    .A3(\hash/_1617_ ),
    .B1(\hash/_0575_ ),
    .Y(\hash/_0576_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3356_  (.A1(\hash/_0563_ ),
    .A2(\hash/_0574_ ),
    .B1(\hash/_0576_ ),
    .Y(\hash/_0577_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3357_  (.A(\hash/_1624_ ),
    .B(\hash/_0577_ ),
    .X(\hash/_0064_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3358_  (.A1(\hash/_1624_ ),
    .A2(\hash/_1621_ ),
    .B1(\hash/_1623_ ),
    .Y(\hash/_0578_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3359_  (.A(\hash/_0578_ ),
    .Y(\hash/_0579_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3360_  (.A1(\hash/_1622_ ),
    .A2(\hash/_1624_ ),
    .A3(\hash/_0572_ ),
    .B1(\hash/_0579_ ),
    .Y(\hash/_0580_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3361_  (.A(\hash/_1628_ ),
    .B(\hash/_0580_ ),
    .Y(\hash/_0065_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3362_  (.A(\hash/_1620_ ),
    .B(\hash/_1622_ ),
    .C(\hash/_1624_ ),
    .Y(\hash/_0581_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3363_  (.A1(\hash/_1624_ ),
    .A2(\hash/_0575_ ),
    .B1(\hash/_1623_ ),
    .Y(\hash/_0582_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3364_  (.A1(\hash/_0565_ ),
    .A2(\hash/_0581_ ),
    .B1(\hash/_0582_ ),
    .Y(\hash/_0583_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3365_  (.A1(\hash/_1628_ ),
    .A2(\hash/_0583_ ),
    .B1(\hash/_1627_ ),
    .Y(\hash/_0584_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3366_  (.A(\hash/_1626_ ),
    .B(\hash/_0584_ ),
    .Y(\hash/_0066_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3367_  (.A(\hash/_1628_ ),
    .Y(\hash/_0585_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3368_  (.A1(\hash/_0585_ ),
    .A2(\hash/_0580_ ),
    .B1_N(\hash/_1627_ ),
    .Y(\hash/_0586_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3369_  (.A1(\hash/_1626_ ),
    .A2(\hash/_0586_ ),
    .B1(\hash/_1625_ ),
    .Y(\hash/_0587_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3370_  (.A(\hash/_1630_ ),
    .B(\hash/_0587_ ),
    .Y(\hash/_0067_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3372_  (.A(\hash/_1626_ ),
    .B(\hash/_1630_ ),
    .Y(\hash/_0589_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3373_  (.A1(\hash/_1628_ ),
    .A2(\hash/_1623_ ),
    .B1(\hash/_1627_ ),
    .Y(\hash/_0590_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3374_  (.A1(\hash/_1630_ ),
    .A2(\hash/_1625_ ),
    .B1(\hash/_1629_ ),
    .Y(\hash/_0591_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3375_  (.A1(\hash/_0589_ ),
    .A2(\hash/_0590_ ),
    .B1(\hash/_0591_ ),
    .Y(\hash/_0592_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3376_  (.A(\hash/_0585_ ),
    .B(\hash/_0589_ ),
    .Y(\hash/_0593_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3377_  (.A(\hash/_1624_ ),
    .B(\hash/_0593_ ),
    .Y(\hash/_0594_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3378_  (.A(\hash/_0594_ ),
    .B_N(\hash/_0577_ ),
    .Y(\hash/_0595_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3379_  (.A(\hash/_0592_ ),
    .B(\hash/_0595_ ),
    .Y(\hash/_0596_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3380_  (.A(\hash/_1632_ ),
    .B(\hash/_0596_ ),
    .Y(\hash/_0068_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3381_  (.A(\hash/_1634_ ),
    .Y(\hash/_0597_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3382_  (.A(\hash/_1622_ ),
    .B(\hash/_1624_ ),
    .C(\hash/_1632_ ),
    .D(\hash/_0593_ ),
    .Y(\hash/_0598_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3383_  (.A1(\hash/_0550_ ),
    .A2(\hash/_0568_ ),
    .B1(\hash/_0571_ ),
    .C1(\hash/_0598_ ),
    .Y(\hash/_0599_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3384_  (.A1(\hash/_1626_ ),
    .A2(\hash/_1627_ ),
    .B1(\hash/_1625_ ),
    .X(\hash/_0600_ ));
 sky130_fd_sc_hd__a221o_1 \hash/_3385_  (.A1(\hash/_0579_ ),
    .A2(\hash/_0593_ ),
    .B1(\hash/_0600_ ),
    .B2(\hash/_1630_ ),
    .C1(\hash/_1629_ ),
    .X(\hash/_0601_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3386_  (.A1(\hash/_1632_ ),
    .A2(\hash/_0601_ ),
    .B1(\hash/_1631_ ),
    .Y(\hash/_0602_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3387_  (.A_N(\hash/_0599_ ),
    .B(\hash/_0602_ ),
    .Y(\hash/_0603_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3388_  (.A(\hash/_0597_ ),
    .B(\hash/_0603_ ),
    .Y(\hash/_0069_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3389_  (.A1(\hash/_0592_ ),
    .A2(\hash/_0595_ ),
    .B1(\hash/_1632_ ),
    .Y(\hash/_0604_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3390_  (.A(\hash/_1636_ ),
    .Y(\hash/_0605_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3391_  (.A(\hash/_0605_ ),
    .B(\hash/_1631_ ),
    .C(\hash/_1633_ ),
    .Y(\hash/_0606_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3392_  (.A(\hash/_0604_ ),
    .B(\hash/_0606_ ),
    .Y(\hash/_0607_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3393_  (.A(\hash/_0597_ ),
    .B(\hash/_1636_ ),
    .Y(\hash/_0608_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3394_  (.A(\hash/_1634_ ),
    .B(\hash/_0605_ ),
    .C(\hash/_1633_ ),
    .Y(\hash/_0609_ ));
 sky130_fd_sc_hd__a221oi_1 \hash/_3395_  (.A1(\hash/_0605_ ),
    .A2(\hash/_1633_ ),
    .B1(\hash/_0608_ ),
    .B2(\hash/_1631_ ),
    .C1(\hash/_0609_ ),
    .Y(\hash/_0610_ ));
 sky130_fd_sc_hd__o311ai_1 \hash/_3396_  (.A1(\hash/_0597_ ),
    .A2(\hash/_1636_ ),
    .A3(\hash/_0604_ ),
    .B1(\hash/_0607_ ),
    .C1(\hash/_0610_ ),
    .Y(\hash/_0070_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3397_  (.A1(\hash/_1634_ ),
    .A2(\hash/_0603_ ),
    .B1(\hash/_1633_ ),
    .X(\hash/_0611_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3398_  (.A1(\hash/_1636_ ),
    .A2(\hash/_0611_ ),
    .B1(\hash/_1635_ ),
    .Y(\hash/_0612_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3399_  (.A(\hash/_1638_ ),
    .B(\hash/_0612_ ),
    .Y(\hash/_0071_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3400_  (.A(\hash/_1634_ ),
    .B(\hash/_1636_ ),
    .C(\hash/_1638_ ),
    .X(\hash/_0613_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3401_  (.A1(\hash/_1632_ ),
    .A2(\hash/_0592_ ),
    .B1(\hash/_1631_ ),
    .X(\hash/_0614_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3402_  (.A1(\hash/_1634_ ),
    .A2(\hash/_0614_ ),
    .B1(\hash/_1633_ ),
    .Y(\hash/_0615_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3403_  (.A(\hash/_1636_ ),
    .B(\hash/_1638_ ),
    .Y(\hash/_0616_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3404_  (.A1(\hash/_1638_ ),
    .A2(\hash/_1635_ ),
    .B1(\hash/_1637_ ),
    .Y(\hash/_0617_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3405_  (.A1(\hash/_0615_ ),
    .A2(\hash/_0616_ ),
    .B1(\hash/_0617_ ),
    .Y(\hash/_0618_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3406_  (.A1(\hash/_1632_ ),
    .A2(\hash/_0595_ ),
    .A3(\hash/_0613_ ),
    .B1(\hash/_0618_ ),
    .Y(\hash/_0619_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3407_  (.A(\hash/_1640_ ),
    .B(\hash/_0619_ ),
    .Y(\hash/_0072_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3408_  (.A1(\hash/_1636_ ),
    .A2(\hash/_1633_ ),
    .B1(\hash/_1635_ ),
    .X(\hash/_0620_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3409_  (.A1(\hash/_1638_ ),
    .A2(\hash/_1640_ ),
    .A3(\hash/_0620_ ),
    .B1(\hash/_1639_ ),
    .Y(\hash/_0621_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3410_  (.A(\hash/_1634_ ),
    .B(\hash/_1636_ ),
    .C(\hash/_1638_ ),
    .Y(\hash/_0622_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3411_  (.A(\hash/_0602_ ),
    .B(\hash/_0622_ ),
    .Y(\hash/_0623_ ));
 sky130_fd_sc_hd__or3_1 \hash/_3412_  (.A(\hash/_0571_ ),
    .B(\hash/_0598_ ),
    .C(\hash/_0622_ ),
    .X(\hash/_0624_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3413_  (.A1(\hash/_0550_ ),
    .A2(\hash/_0568_ ),
    .B1(\hash/_0624_ ),
    .Y(\hash/_0625_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_3414_  (.A1(\hash/_1637_ ),
    .A2(\hash/_0623_ ),
    .A3(\hash/_0625_ ),
    .B1(\hash/_1640_ ),
    .Y(\hash/_0626_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3415_  (.A(\hash/_0621_ ),
    .B(\hash/_0626_ ),
    .Y(\hash/_0627_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3416_  (.A(\hash/_1642_ ),
    .B(\hash/_0627_ ),
    .X(\hash/_0073_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3417_  (.A(\hash/_1644_ ),
    .Y(\hash/_0628_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3418_  (.A1(\hash/_1642_ ),
    .A2(\hash/_1639_ ),
    .B1(\hash/_1641_ ),
    .Y(\hash/_0629_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3419_  (.A(\hash/_1632_ ),
    .B(\hash/_1640_ ),
    .C(\hash/_1642_ ),
    .Y(\hash/_0630_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3420_  (.A(\hash/_0594_ ),
    .B(\hash/_0622_ ),
    .C(\hash/_0630_ ),
    .Y(\hash/_0631_ ));
 sky130_fd_sc_hd__a32oi_1 \hash/_3421_  (.A1(\hash/_1640_ ),
    .A2(\hash/_1642_ ),
    .A3(\hash/_0618_ ),
    .B1(\hash/_0631_ ),
    .B2(\hash/_0577_ ),
    .Y(\hash/_0632_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3422_  (.A(\hash/_0629_ ),
    .B(\hash/_0632_ ),
    .Y(\hash/_0633_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3423_  (.A(\hash/_0628_ ),
    .B(\hash/_0633_ ),
    .Y(\hash/_0074_ ));
 sky130_fd_sc_hd__nor4b_2 \hash/_3424_  (.A(\hash/_1637_ ),
    .B(\hash/_0623_ ),
    .C(\hash/_0625_ ),
    .D_N(\hash/_0621_ ),
    .Y(\hash/_0634_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3425_  (.A1(\hash/_1640_ ),
    .A2(\hash/_1639_ ),
    .B1(\hash/_1642_ ),
    .Y(\hash/_0635_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3426_  (.A1(\hash/_0634_ ),
    .A2(\hash/_0635_ ),
    .B1_N(\hash/_1641_ ),
    .Y(\hash/_0636_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3427_  (.A1(\hash/_1644_ ),
    .A2(\hash/_0636_ ),
    .B1(\hash/_1643_ ),
    .Y(\hash/_0637_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3428_  (.A(\hash/_1646_ ),
    .B(\hash/_0637_ ),
    .Y(\hash/_0075_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3429_  (.A(\hash/_1648_ ),
    .Y(\hash/_0638_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3430_  (.A(\hash/_1644_ ),
    .B(\hash/_1646_ ),
    .Y(\hash/_0639_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3431_  (.A1(\hash/_0628_ ),
    .A2(\hash/_0629_ ),
    .B1_N(\hash/_1643_ ),
    .Y(\hash/_0640_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3432_  (.A1(\hash/_1646_ ),
    .A2(\hash/_0640_ ),
    .B1(\hash/_1645_ ),
    .Y(\hash/_0641_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3433_  (.A1(\hash/_0632_ ),
    .A2(\hash/_0639_ ),
    .B1(\hash/_0641_ ),
    .Y(\hash/_0642_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3434_  (.A(\hash/_0638_ ),
    .B(\hash/_0642_ ),
    .Y(\hash/_0076_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3435_  (.A1(\hash/_1644_ ),
    .A2(\hash/_1641_ ),
    .B1(\hash/_1643_ ),
    .X(\hash/_0643_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3436_  (.A1(\hash/_1646_ ),
    .A2(\hash/_0643_ ),
    .B1(\hash/_1645_ ),
    .Y(\hash/_0644_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3437_  (.A1(\hash/_0638_ ),
    .A2(\hash/_0644_ ),
    .B1_N(\hash/_1647_ ),
    .Y(\hash/_0645_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3438_  (.A(\hash/_1644_ ),
    .B(\hash/_1646_ ),
    .C(\hash/_1648_ ),
    .Y(\hash/_0646_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3439_  (.A(\hash/_0634_ ),
    .B(\hash/_0635_ ),
    .C(\hash/_0646_ ),
    .Y(\hash/_0647_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3440_  (.A(\hash/_0645_ ),
    .B(\hash/_0647_ ),
    .Y(\hash/_0648_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3441_  (.A(\hash/_1650_ ),
    .B(\hash/_0648_ ),
    .Y(\hash/_0077_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3442_  (.A1(\hash/_1646_ ),
    .A2(\hash/_1643_ ),
    .B1(\hash/_1645_ ),
    .Y(\hash/_0649_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3443_  (.A(\hash/_1647_ ),
    .B(\hash/_1649_ ),
    .Y(\hash/_0650_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3444_  (.A1(\hash/_0638_ ),
    .A2(\hash/_0649_ ),
    .B1(\hash/_0650_ ),
    .Y(\hash/_0651_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3445_  (.A1(\hash/_0629_ ),
    .A2(\hash/_0632_ ),
    .B1(\hash/_0646_ ),
    .Y(\hash/_0652_ ));
 sky130_fd_sc_hd__o22ai_1 \hash/_3446_  (.A1(\hash/_1650_ ),
    .A2(\hash/_1649_ ),
    .B1(\hash/_0651_ ),
    .B2(\hash/_0652_ ),
    .Y(\hash/_0653_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3447_  (.A(\hash/_1652_ ),
    .B(\hash/_0653_ ),
    .Y(\hash/_0078_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3448_  (.A1(\hash/_1650_ ),
    .A2(\hash/_1649_ ),
    .B1(\hash/_1652_ ),
    .Y(\hash/_0654_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3449_  (.A_N(\hash/_1651_ ),
    .B(\hash/_0654_ ),
    .Y(\hash/_0655_ ));
 sky130_fd_sc_hd__o41ai_1 \hash/_3450_  (.A1(\hash/_1649_ ),
    .A2(\hash/_1651_ ),
    .A3(\hash/_0645_ ),
    .A4(\hash/_0647_ ),
    .B1(\hash/_0655_ ),
    .Y(\hash/_0656_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3451_  (.A(\hash/_1654_ ),
    .B(\hash/_0656_ ),
    .Y(\hash/_0079_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3452_  (.A(\hash/_1650_ ),
    .B(\hash/_1652_ ),
    .C(\hash/_1654_ ),
    .Y(\hash/_0657_ ));
 sky130_fd_sc_hd__or2_2 \hash/_3453_  (.A(\hash/_0646_ ),
    .B(\hash/_0657_ ),
    .X(\hash/_0658_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3454_  (.A1(\hash/_1652_ ),
    .A2(\hash/_1649_ ),
    .B1(\hash/_1651_ ),
    .C1(\hash/_1647_ ),
    .Y(\hash/_0659_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3455_  (.A1(\hash/_0638_ ),
    .A2(\hash/_0641_ ),
    .B1(\hash/_0659_ ),
    .Y(\hash/_0660_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3456_  (.A1(\hash/_1654_ ),
    .A2(\hash/_0655_ ),
    .A3(\hash/_0660_ ),
    .B1(\hash/_1653_ ),
    .Y(\hash/_0661_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3457_  (.A1(\hash/_0632_ ),
    .A2(\hash/_0658_ ),
    .B1(\hash/_0661_ ),
    .Y(\hash/_0662_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3458_  (.A(\hash/_1656_ ),
    .B(\hash/_0662_ ),
    .X(\hash/_0081_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_3460_  (.A0(\hash/a_cap[31] ),
    .A1(_09578_),
    .S(reset_hash_dash),
    .X(\hash/c[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3461_  (.A(_09578_),
    .B(\hash/a_cap[31] ),
    .Y(\hash/_0664_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3462_  (.A(reset_hash_dash),
    .B(\hash/_0664_ ),
    .Y(\hash/_0665_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3463_  (.A1(\hash/_1650_ ),
    .A2(\hash/_0645_ ),
    .B1(\hash/_1649_ ),
    .X(\hash/_0666_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3464_  (.A1(\hash/_1652_ ),
    .A2(\hash/_0666_ ),
    .B1(\hash/_1651_ ),
    .X(\hash/_0667_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3465_  (.A1(\hash/_1654_ ),
    .A2(\hash/_0667_ ),
    .B1(\hash/_1653_ ),
    .Y(\hash/_0668_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_3466_  (.A1(\hash/_0634_ ),
    .A2(\hash/_0635_ ),
    .A3(\hash/_0658_ ),
    .B1(\hash/_0668_ ),
    .Y(\hash/_0669_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3467_  (.A1(\hash/_1656_ ),
    .A2(\hash/_0669_ ),
    .B1(\hash/_1655_ ),
    .Y(\hash/_0670_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3468_  (.A(\hash/_0665_ ),
    .B(\hash/_0670_ ),
    .Y(\hash/_0082_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3469_  (.A(\hash/_1468_ ),
    .B(\hash/_1662_ ),
    .X(\hash/_0110_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3470_  (.A1(\hash/_1467_ ),
    .A2(\hash/_1658_ ),
    .B1(\hash/_1657_ ),
    .X(\hash/_0671_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3471_  (.A1(\hash/_1662_ ),
    .A2(\hash/_0671_ ),
    .B1(\hash/_1661_ ),
    .Y(\hash/_0672_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3472_  (.A(\hash/_1660_ ),
    .B(\hash/_0672_ ),
    .Y(\hash/_0113_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3473_  (.A1(\hash/_1468_ ),
    .A2(\hash/_1662_ ),
    .B1(\hash/_1659_ ),
    .C1(\hash/_1661_ ),
    .Y(\hash/_0673_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3474_  (.A1(\hash/_1660_ ),
    .A2(\hash/_1659_ ),
    .B1(\hash/_1664_ ),
    .Y(\hash/_0674_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3475_  (.A(\hash/_0673_ ),
    .B(\hash/_0674_ ),
    .Y(\hash/_0675_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3476_  (.A1(\hash/_1468_ ),
    .A2(\hash/_1662_ ),
    .B1(\hash/_1661_ ),
    .X(\hash/_0676_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3477_  (.A1(\hash/_1660_ ),
    .A2(\hash/_0676_ ),
    .B1(\hash/_1659_ ),
    .C1(\hash/_1664_ ),
    .Y(\hash/_0677_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3478_  (.A(\hash/_0675_ ),
    .B(\hash/_0677_ ),
    .Y(\hash/_0114_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3480_  (.A(\hash/_0672_ ),
    .B_N(\hash/_1660_ ),
    .Y(\hash/_0679_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3481_  (.A1(\hash/_1659_ ),
    .A2(\hash/_0679_ ),
    .B1(\hash/_1664_ ),
    .X(\hash/_0680_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3482_  (.A(\hash/_1663_ ),
    .B(\hash/_0680_ ),
    .Y(\hash/_0681_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3483_  (.A(\hash/_1666_ ),
    .B(\hash/_0681_ ),
    .Y(\hash/_0115_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3484_  (.A1(\hash/_1663_ ),
    .A2(\hash/_0675_ ),
    .B1(\hash/_1666_ ),
    .X(\hash/_0682_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3485_  (.A(\hash/_1665_ ),
    .B(\hash/_0682_ ),
    .Y(\hash/_0683_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3486_  (.A(\hash/_1668_ ),
    .B(\hash/_0683_ ),
    .Y(\hash/_0116_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3487_  (.A(\hash/_1666_ ),
    .Y(\hash/_0684_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3488_  (.A1(\hash/_0684_ ),
    .A2(\hash/_0681_ ),
    .B1_N(\hash/_1665_ ),
    .Y(\hash/_0685_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3489_  (.A1(\hash/_1668_ ),
    .A2(\hash/_0685_ ),
    .B1(\hash/_1667_ ),
    .Y(\hash/_0686_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3490_  (.A(\hash/_1670_ ),
    .B(\hash/_0686_ ),
    .Y(\hash/_0117_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3491_  (.A(\hash/_1668_ ),
    .Y(\hash/_0687_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3492_  (.A1(\hash/_0687_ ),
    .A2(\hash/_0683_ ),
    .B1_N(\hash/_1667_ ),
    .Y(\hash/_0688_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3493_  (.A1(\hash/_1670_ ),
    .A2(\hash/_0688_ ),
    .B1(\hash/_1669_ ),
    .Y(\hash/_0689_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3494_  (.A(\hash/_1672_ ),
    .B(\hash/_0689_ ),
    .Y(\hash/_0118_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3495_  (.A(\hash/_1668_ ),
    .B(\hash/_1670_ ),
    .C(\hash/_1672_ ),
    .Y(\hash/_0690_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3496_  (.A(\hash/_1664_ ),
    .B(\hash/_1666_ ),
    .Y(\hash/_0691_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3497_  (.A(\hash/_0690_ ),
    .B(\hash/_0691_ ),
    .Y(\hash/_0692_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3498_  (.A(\hash/_1666_ ),
    .B(\hash/_1663_ ),
    .Y(\hash/_0693_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3499_  (.A(\hash/_1664_ ),
    .B(\hash/_1666_ ),
    .C(\hash/_1659_ ),
    .Y(\hash/_0694_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3500_  (.A1(\hash/_0693_ ),
    .A2(\hash/_0694_ ),
    .B1(\hash/_0690_ ),
    .Y(\hash/_0695_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3501_  (.A1(\hash/_0679_ ),
    .A2(\hash/_0692_ ),
    .B1(\hash/_0695_ ),
    .Y(\hash/_0696_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3502_  (.A1(\hash/_1668_ ),
    .A2(\hash/_1665_ ),
    .B1(\hash/_1667_ ),
    .X(\hash/_0697_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3503_  (.A1(\hash/_1670_ ),
    .A2(\hash/_0697_ ),
    .B1(\hash/_1669_ ),
    .X(\hash/_0698_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3504_  (.A1(\hash/_1672_ ),
    .A2(\hash/_0698_ ),
    .B1(\hash/_1671_ ),
    .Y(\hash/_0699_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3505_  (.A(\hash/_0696_ ),
    .B(\hash/_0699_ ),
    .Y(\hash/_0700_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3506_  (.A(\hash/_1674_ ),
    .B(\hash/_0700_ ),
    .X(\hash/_0119_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3507_  (.A(\hash/_1672_ ),
    .Y(\hash/_0701_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3508_  (.A1(\hash/_0701_ ),
    .A2(\hash/_0689_ ),
    .B1_N(\hash/_1671_ ),
    .Y(\hash/_0702_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3509_  (.A1(\hash/_1674_ ),
    .A2(\hash/_0702_ ),
    .B1(\hash/_1673_ ),
    .Y(\hash/_0703_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3510_  (.A(\hash/_1676_ ),
    .B(\hash/_0703_ ),
    .Y(\hash/_0090_ ));
 sky130_fd_sc_hd__nor3b_1 \hash/_3511_  (.A(\hash/_1673_ ),
    .B(\hash/_1675_ ),
    .C_N(\hash/_0699_ ),
    .Y(\hash/_0704_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3512_  (.A1(\hash/_1674_ ),
    .A2(\hash/_1673_ ),
    .B1(\hash/_1676_ ),
    .X(\hash/_0705_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3513_  (.A(\hash/_1675_ ),
    .B(\hash/_0705_ ),
    .Y(\hash/_0706_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3514_  (.A(\hash/_1678_ ),
    .Y(\hash/_0707_ ));
 sky130_fd_sc_hd__a211oi_2 \hash/_3515_  (.A1(\hash/_0696_ ),
    .A2(\hash/_0704_ ),
    .B1(\hash/_0706_ ),
    .C1(\hash/_0707_ ),
    .Y(\hash/_0708_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3516_  (.A1(\hash/_0696_ ),
    .A2(\hash/_0704_ ),
    .B1(\hash/_0706_ ),
    .Y(\hash/_0709_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3517_  (.A(\hash/_1678_ ),
    .B(\hash/_0709_ ),
    .Y(\hash/_0710_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3518_  (.A(\hash/_0708_ ),
    .B(\hash/_0710_ ),
    .Y(\hash/_0091_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3519_  (.A(\hash/_1674_ ),
    .B(\hash/_1676_ ),
    .Y(\hash/_0711_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3520_  (.A(\hash/_1666_ ),
    .B(\hash/_1665_ ),
    .Y(\hash/_0712_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3521_  (.A(\hash/_0690_ ),
    .B(\hash/_0711_ ),
    .C(\hash/_0712_ ),
    .Y(\hash/_0713_ ));
 sky130_fd_sc_hd__o31ai_1 \hash/_3522_  (.A1(\hash/_1663_ ),
    .A2(\hash/_1665_ ),
    .A3(\hash/_0675_ ),
    .B1(\hash/_0713_ ),
    .Y(\hash/_0714_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3523_  (.A1(\hash/_1670_ ),
    .A2(\hash/_1667_ ),
    .B1(\hash/_1669_ ),
    .X(\hash/_0715_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3524_  (.A1(\hash/_1672_ ),
    .A2(\hash/_0715_ ),
    .B1(\hash/_1671_ ),
    .Y(\hash/_0716_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3525_  (.A1(\hash/_1676_ ),
    .A2(\hash/_1673_ ),
    .B1(\hash/_1675_ ),
    .Y(\hash/_0717_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3526_  (.A1(\hash/_0711_ ),
    .A2(\hash/_0716_ ),
    .B1(\hash/_0717_ ),
    .X(\hash/_0718_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3527_  (.A1(\hash/_0714_ ),
    .A2(\hash/_0718_ ),
    .B1(\hash/_0707_ ),
    .Y(\hash/_0719_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3528_  (.A(\hash/_1677_ ),
    .B(\hash/_0719_ ),
    .Y(\hash/_0720_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3529_  (.A(\hash/_1680_ ),
    .B(\hash/_0720_ ),
    .Y(\hash/_0092_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3530_  (.A1(\hash/_1677_ ),
    .A2(\hash/_0708_ ),
    .B1(\hash/_1680_ ),
    .X(\hash/_0721_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3531_  (.A(\hash/_1679_ ),
    .B(\hash/_0721_ ),
    .Y(\hash/_0722_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3532_  (.A(\hash/_1682_ ),
    .B(\hash/_0722_ ),
    .Y(\hash/_0093_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3533_  (.A(\hash/_1677_ ),
    .B(\hash/_1679_ ),
    .Y(\hash/_0723_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3534_  (.A1(\hash/_1678_ ),
    .A2(\hash/_1677_ ),
    .B1(\hash/_1680_ ),
    .X(\hash/_0724_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3535_  (.A1(\hash/_1679_ ),
    .A2(\hash/_0724_ ),
    .B1(\hash/_1682_ ),
    .Y(\hash/_0725_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3536_  (.A1(\hash/_0714_ ),
    .A2(\hash/_0718_ ),
    .A3(\hash/_0723_ ),
    .B1(\hash/_0725_ ),
    .Y(\hash/_0726_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3537_  (.A(\hash/_1681_ ),
    .B(\hash/_0726_ ),
    .Y(\hash/_0727_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3538_  (.A(\hash/_1684_ ),
    .B(\hash/_0727_ ),
    .Y(\hash/_0094_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3539_  (.A1(\hash/_1680_ ),
    .A2(\hash/_1677_ ),
    .B1(\hash/_1679_ ),
    .X(\hash/_0728_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3540_  (.A(\hash/_1682_ ),
    .B(\hash/_0728_ ),
    .Y(\hash/_0729_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3541_  (.A(\hash/_0729_ ),
    .Y(\hash/_0730_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3542_  (.A1(\hash/_1680_ ),
    .A2(\hash/_1682_ ),
    .A3(\hash/_0708_ ),
    .B1(\hash/_0730_ ),
    .Y(\hash/_0731_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3543_  (.A_N(\hash/_1681_ ),
    .B(\hash/_0731_ ),
    .Y(\hash/_0732_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3544_  (.A1(\hash/_1684_ ),
    .A2(\hash/_0732_ ),
    .B1(\hash/_1683_ ),
    .Y(\hash/_0733_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3545_  (.A(\hash/_1688_ ),
    .B(\hash/_0733_ ),
    .Y(\hash/_0095_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3546_  (.A1(\hash/_1684_ ),
    .A2(\hash/_1683_ ),
    .B1(\hash/_1688_ ),
    .Y(\hash/_0734_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3547_  (.A(\hash/_0734_ ),
    .Y(\hash/_0735_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3548_  (.A(\hash/_1681_ ),
    .B(\hash/_1683_ ),
    .Y(\hash/_0736_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3549_  (.A_N(\hash/_0726_ ),
    .B(\hash/_0736_ ),
    .Y(\hash/_0737_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3550_  (.A1(\hash/_0735_ ),
    .A2(\hash/_0737_ ),
    .B1(\hash/_1687_ ),
    .Y(\hash/_0738_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3551_  (.A(\hash/_1686_ ),
    .B(\hash/_0738_ ),
    .Y(\hash/_0096_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3552_  (.A1(\hash/_1688_ ),
    .A2(\hash/_1683_ ),
    .B1(\hash/_1687_ ),
    .X(\hash/_0739_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3553_  (.A1(\hash/_1686_ ),
    .A2(\hash/_0739_ ),
    .B1(\hash/_1685_ ),
    .X(\hash/_0740_ ));
 sky130_fd_sc_hd__a41oi_1 \hash/_3554_  (.A1(\hash/_1684_ ),
    .A2(\hash/_1688_ ),
    .A3(\hash/_1686_ ),
    .A4(\hash/_0732_ ),
    .B1(\hash/_0740_ ),
    .Y(\hash/_0741_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3555_  (.A(\hash/_1690_ ),
    .B(\hash/_0741_ ),
    .Y(\hash/_0097_ ));
 sky130_fd_sc_hd__and4_1 \hash/_3556_  (.A(\hash/_1684_ ),
    .B(\hash/_1688_ ),
    .C(\hash/_1686_ ),
    .D(\hash/_1690_ ),
    .X(\hash/_0742_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3557_  (.A1(\hash/_1681_ ),
    .A2(\hash/_0726_ ),
    .B1(\hash/_0742_ ),
    .Y(\hash/_0743_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3558_  (.A1(\hash/_1690_ ),
    .A2(\hash/_0740_ ),
    .B1(\hash/_1689_ ),
    .Y(\hash/_0744_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3559_  (.A(\hash/_0743_ ),
    .B(\hash/_0744_ ),
    .Y(\hash/_0745_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3560_  (.A(\hash/_1692_ ),
    .B(\hash/_0745_ ),
    .X(\hash/_0098_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3561_  (.A1(\hash/_1686_ ),
    .A2(\hash/_1687_ ),
    .B1(\hash/_1685_ ),
    .X(\hash/_0746_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3562_  (.A1(\hash/_1690_ ),
    .A2(\hash/_0746_ ),
    .B1(\hash/_1689_ ),
    .X(\hash/_0747_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3563_  (.A1(\hash/_1692_ ),
    .A2(\hash/_0747_ ),
    .B1(\hash/_1691_ ),
    .Y(\hash/_0748_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3564_  (.A(\hash/_1686_ ),
    .B(\hash/_1690_ ),
    .C(\hash/_1692_ ),
    .D(\hash/_0735_ ),
    .Y(\hash/_0749_ ));
 sky130_fd_sc_hd__and2_1 \hash/_3565_  (.A(\hash/_0748_ ),
    .B(\hash/_0749_ ),
    .X(\hash/_0750_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3566_  (.A(\hash/_0729_ ),
    .B(\hash/_0736_ ),
    .C(\hash/_0748_ ),
    .Y(\hash/_0751_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3567_  (.A1(\hash/_1680_ ),
    .A2(\hash/_1682_ ),
    .A3(\hash/_0708_ ),
    .B1(\hash/_0751_ ),
    .Y(\hash/_0752_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3568_  (.A(\hash/_0750_ ),
    .B(\hash/_0752_ ),
    .Y(\hash/_0753_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3569_  (.A(\hash/_1694_ ),
    .B(\hash/_0753_ ),
    .X(\hash/_0099_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3570_  (.A1(\hash/_1692_ ),
    .A2(\hash/_0745_ ),
    .B1(\hash/_1691_ ),
    .X(\hash/_0754_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3571_  (.A1(\hash/_1694_ ),
    .A2(\hash/_0754_ ),
    .B1(\hash/_1693_ ),
    .Y(\hash/_0755_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3572_  (.A(\hash/_1696_ ),
    .B(\hash/_0755_ ),
    .Y(\hash/_0100_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3573_  (.A1(\hash/_1696_ ),
    .A2(\hash/_1693_ ),
    .B1(\hash/_1695_ ),
    .Y(\hash/_0756_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3574_  (.A1(\hash/_1696_ ),
    .A2(\hash/_1693_ ),
    .B1(\hash/_1695_ ),
    .X(\hash/_0757_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3575_  (.A1(\hash/_1694_ ),
    .A2(\hash/_1696_ ),
    .B1(\hash/_0757_ ),
    .Y(\hash/_0758_ ));
 sky130_fd_sc_hd__a31o_1 \hash/_3576_  (.A1(\hash/_0748_ ),
    .A2(\hash/_0749_ ),
    .A3(\hash/_0756_ ),
    .B1(\hash/_0758_ ),
    .X(\hash/_0759_ ));
 sky130_fd_sc_hd__a41o_1 \hash/_3577_  (.A1(\hash/_0731_ ),
    .A2(\hash/_0736_ ),
    .A3(\hash/_0748_ ),
    .A4(\hash/_0756_ ),
    .B1(\hash/_0759_ ),
    .X(\hash/_0760_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3578_  (.A(\hash/_1698_ ),
    .B(\hash/_0760_ ),
    .Y(\hash/_0101_ ));
 sky130_fd_sc_hd__and3_1 \hash/_3579_  (.A(\hash/_1692_ ),
    .B(\hash/_1694_ ),
    .C(\hash/_1696_ ),
    .X(\hash/_0761_ ));
 sky130_fd_sc_hd__o211ai_1 \hash/_3580_  (.A1(\hash/_1681_ ),
    .A2(\hash/_0726_ ),
    .B1(\hash/_0742_ ),
    .C1(\hash/_0761_ ),
    .Y(\hash/_0762_ ));
 sky130_fd_sc_hd__nand2b_1 \hash/_3581_  (.A_N(\hash/_0744_ ),
    .B(\hash/_1692_ ),
    .Y(\hash/_0763_ ));
 sky130_fd_sc_hd__nor3_1 \hash/_3582_  (.A(\hash/_1691_ ),
    .B(\hash/_1693_ ),
    .C(\hash/_1695_ ),
    .Y(\hash/_0764_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3583_  (.A1(\hash/_0763_ ),
    .A2(\hash/_0764_ ),
    .B1(\hash/_0758_ ),
    .X(\hash/_0765_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3584_  (.A(\hash/_0762_ ),
    .B(\hash/_0765_ ),
    .Y(\hash/_0766_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3585_  (.A1(\hash/_1698_ ),
    .A2(\hash/_0766_ ),
    .B1(\hash/_1697_ ),
    .X(\hash/_0767_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3586_  (.A(\hash/_1700_ ),
    .B(\hash/_0767_ ),
    .X(\hash/_0102_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3587_  (.A(\hash/_1694_ ),
    .B(\hash/_1696_ ),
    .Y(\hash/_0768_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3588_  (.A(\hash/_1698_ ),
    .B(\hash/_1700_ ),
    .Y(\hash/_0769_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3589_  (.A1(\hash/_1698_ ),
    .A2(\hash/_0757_ ),
    .B1(\hash/_1697_ ),
    .X(\hash/_0770_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3590_  (.A1(\hash/_1700_ ),
    .A2(\hash/_0770_ ),
    .B1(\hash/_1699_ ),
    .Y(\hash/_0771_ ));
 sky130_fd_sc_hd__o41a_1 \hash/_3591_  (.A1(\hash/_0750_ ),
    .A2(\hash/_0752_ ),
    .A3(\hash/_0768_ ),
    .A4(\hash/_0769_ ),
    .B1(\hash/_0771_ ),
    .X(\hash/_0772_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3592_  (.A(\hash/_1702_ ),
    .B(\hash/_0772_ ),
    .Y(\hash/_0103_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3594_  (.A1(\hash/_1702_ ),
    .A2(\hash/_1699_ ),
    .B1(\hash/_1701_ ),
    .X(\hash/_0774_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3595_  (.A(\hash/_1697_ ),
    .B(\hash/_0774_ ),
    .Y(\hash/_0775_ ));
 sky130_fd_sc_hd__and2_1 \hash/_3596_  (.A(\hash/_1700_ ),
    .B(\hash/_1702_ ),
    .X(\hash/_0776_ ));
 sky130_fd_sc_hd__or2_2 \hash/_3597_  (.A(\hash/_1698_ ),
    .B(\hash/_1697_ ),
    .X(\hash/_0777_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3598_  (.A1(\hash/_0776_ ),
    .A2(\hash/_0777_ ),
    .B1(\hash/_0774_ ),
    .Y(\hash/_0778_ ));
 sky130_fd_sc_hd__a31o_1 \hash/_3599_  (.A1(\hash/_0762_ ),
    .A2(\hash/_0765_ ),
    .A3(\hash/_0775_ ),
    .B1(\hash/_0778_ ),
    .X(\hash/_0779_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3600_  (.A(\hash/_1704_ ),
    .B(\hash/_0779_ ),
    .Y(\hash/_0104_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3601_  (.A(\hash/_1706_ ),
    .Y(\hash/_0780_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3602_  (.A(\hash/_1702_ ),
    .B(\hash/_1704_ ),
    .Y(\hash/_0781_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3603_  (.A1(\hash/_1704_ ),
    .A2(\hash/_1701_ ),
    .B1(\hash/_1703_ ),
    .Y(\hash/_0782_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3604_  (.A1(\hash/_0772_ ),
    .A2(\hash/_0781_ ),
    .B1(\hash/_0782_ ),
    .Y(\hash/_0783_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3605_  (.A(\hash/_0780_ ),
    .B(\hash/_0783_ ),
    .Y(\hash/_0105_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3607_  (.A1(\hash/_1704_ ),
    .A2(\hash/_0774_ ),
    .B1(\hash/_1703_ ),
    .Y(\hash/_0785_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3608_  (.A1(\hash/_0780_ ),
    .A2(\hash/_0785_ ),
    .B1_N(\hash/_1705_ ),
    .Y(\hash/_0786_ ));
 sky130_fd_sc_hd__a41o_1 \hash/_3609_  (.A1(\hash/_1704_ ),
    .A2(\hash/_1706_ ),
    .A3(\hash/_0767_ ),
    .A4(\hash/_0776_ ),
    .B1(\hash/_0786_ ),
    .X(\hash/_0787_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3610_  (.A(\hash/_1708_ ),
    .B(\hash/_0787_ ),
    .X(\hash/_0106_ ));
 sky130_fd_sc_hd__nand4_1 \hash/_3611_  (.A(\hash/_1702_ ),
    .B(\hash/_1704_ ),
    .C(\hash/_1706_ ),
    .D(\hash/_1708_ ),
    .Y(\hash/_0788_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3612_  (.A1(\hash/_0780_ ),
    .A2(\hash/_0782_ ),
    .B1_N(\hash/_1705_ ),
    .Y(\hash/_0789_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3613_  (.A1(\hash/_1708_ ),
    .A2(\hash/_0789_ ),
    .B1(\hash/_1707_ ),
    .Y(\hash/_0790_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3614_  (.A1(\hash/_0772_ ),
    .A2(\hash/_0788_ ),
    .B1(\hash/_0790_ ),
    .Y(\hash/_0791_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3615_  (.A(\hash/_1710_ ),
    .B(\hash/_0791_ ),
    .X(\hash/_0107_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3616_  (.A(\hash/_1704_ ),
    .B(\hash/_1706_ ),
    .C(\hash/_1708_ ),
    .Y(\hash/_0792_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3617_  (.A1(\hash/_1706_ ),
    .A2(\hash/_1703_ ),
    .B1(\hash/_1705_ ),
    .X(\hash/_0793_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3618_  (.A1(\hash/_1708_ ),
    .A2(\hash/_0793_ ),
    .B1(\hash/_1709_ ),
    .C1(\hash/_1707_ ),
    .Y(\hash/_0794_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3619_  (.A1(\hash/_0779_ ),
    .A2(\hash/_0792_ ),
    .B1(\hash/_0794_ ),
    .Y(\hash/_0795_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3620_  (.A1(\hash/_1710_ ),
    .A2(\hash/_1709_ ),
    .B1(\hash/_0795_ ),
    .Y(\hash/_0796_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3621_  (.A(\hash/_1712_ ),
    .B(\hash/_0796_ ),
    .Y(\hash/_0108_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3622_  (.A(\hash/_1710_ ),
    .B(\hash/_1712_ ),
    .Y(\hash/_0797_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3623_  (.A1(\hash/_1712_ ),
    .A2(\hash/_1709_ ),
    .B1(\hash/_1711_ ),
    .X(\hash/_0798_ ));
 sky130_fd_sc_hd__a41o_1 \hash/_3624_  (.A1(\hash/_1704_ ),
    .A2(\hash/_1706_ ),
    .A3(\hash/_1697_ ),
    .A4(\hash/_0776_ ),
    .B1(\hash/_0786_ ),
    .X(\hash/_0799_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3625_  (.A1(\hash/_1708_ ),
    .A2(\hash/_0799_ ),
    .B1(\hash/_1707_ ),
    .Y(\hash/_0800_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3626_  (.A(\hash/_0800_ ),
    .B(\hash/_0797_ ),
    .Y(\hash/_0801_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3627_  (.A(\hash/_0798_ ),
    .B(\hash/_0801_ ),
    .Y(\hash/_0802_ ));
 sky130_fd_sc_hd__o41ai_1 \hash/_3628_  (.A1(\hash/_0760_ ),
    .A2(\hash/_0769_ ),
    .A3(\hash/_0788_ ),
    .A4(\hash/_0797_ ),
    .B1(\hash/_0802_ ),
    .Y(\hash/_0803_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3629_  (.A(\hash/_1714_ ),
    .B(\hash/_0803_ ),
    .X(\hash/_0109_ ));
 sky130_fd_sc_hd__nand3_1 \hash/_3630_  (.A(\hash/_1710_ ),
    .B(\hash/_1712_ ),
    .C(\hash/_1714_ ),
    .Y(\hash/_0804_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3631_  (.A(\hash/_0792_ ),
    .B(\hash/_0804_ ),
    .Y(\hash/_0805_ ));
 sky130_fd_sc_hd__a211oi_1 \hash/_3632_  (.A1(\hash/_1708_ ),
    .A2(\hash/_0786_ ),
    .B1(\hash/_0798_ ),
    .C1(\hash/_1707_ ),
    .Y(\hash/_0806_ ));
 sky130_fd_sc_hd__o21a_1 \hash/_3633_  (.A1(\hash/_1710_ ),
    .A2(\hash/_1709_ ),
    .B1(\hash/_1712_ ),
    .X(\hash/_0807_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3634_  (.A1(\hash/_1711_ ),
    .A2(\hash/_0807_ ),
    .B1(\hash/_1714_ ),
    .Y(\hash/_0808_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3635_  (.A1(\hash/_0806_ ),
    .A2(\hash/_0808_ ),
    .B1_N(\hash/_1713_ ),
    .Y(\hash/_0809_ ));
 sky130_fd_sc_hd__a31oi_1 \hash/_3636_  (.A1(\hash/_0767_ ),
    .A2(\hash/_0776_ ),
    .A3(\hash/_0805_ ),
    .B1(\hash/_0809_ ),
    .Y(\hash/_0810_ ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3637_  (.A(\hash/_1716_ ),
    .B(\hash/_0810_ ),
    .Y(\hash/_0111_ ));
 sky130_fd_sc_hd__mux2_2 \hash/_3638_  (.A0(\hash/b_cap[31] ),
    .A1(_09577_),
    .S(reset_hash_dash),
    .X(\hash/d[31] ));
 sky130_fd_sc_hd__xnor2_1 \hash/_3639_  (.A(_09577_),
    .B(\hash/b_cap[31] ),
    .Y(\hash/_0811_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3640_  (.A(reset_hash_dash),
    .B(\hash/_0811_ ),
    .Y(\hash/_0812_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3641_  (.A(\hash/_1716_ ),
    .Y(\hash/_0813_ ));
 sky130_fd_sc_hd__o21bai_1 \hash/_3642_  (.A1(\hash/_0790_ ),
    .A2(\hash/_0797_ ),
    .B1_N(\hash/_0798_ ),
    .Y(\hash/_0814_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3643_  (.A1(\hash/_1714_ ),
    .A2(\hash/_0814_ ),
    .B1(\hash/_1713_ ),
    .Y(\hash/_0815_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3644_  (.A(\hash/_0813_ ),
    .B(\hash/_0815_ ),
    .Y(\hash/_0816_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3645_  (.A(\hash/_1715_ ),
    .B(\hash/_0816_ ),
    .Y(\hash/_0817_ ));
 sky130_fd_sc_hd__o41ai_2 \hash/_3646_  (.A1(\hash/_0813_ ),
    .A2(\hash/_0772_ ),
    .A3(\hash/_0788_ ),
    .A4(\hash/_0804_ ),
    .B1(\hash/_0817_ ),
    .Y(\hash/_0818_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3647_  (.A(\hash/_0812_ ),
    .B(\hash/_0818_ ),
    .X(\hash/_0112_ ));
 sky130_fd_sc_hd__xor2_1 \hash/_3648_  (.A(\hash/_1470_ ),
    .B(\hash/_1722_ ),
    .X(\hash/_0140_ ));
 sky130_fd_sc_hd__a21oi_1 \hash/_3649_  (.A1(\hash/_1469_ ),
    .A2(\hash/_1718_ ),
    .B1(\hash/_1717_ ),
    .Y(\hash/_0819_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3650_  (.A(\hash/_1722_ ),
    .B(\hash/_1720_ ),
    .Y(\hash/_0820_ ));
 sky130_fd_sc_hd__nand2_1 \hash/_3651_  (.A(\hash/_1720_ ),
    .B(\hash/_1721_ ),
    .Y(\hash/_0821_ ));
 sky130_fd_sc_hd__o21ai_1 \hash/_3652_  (.A1(\hash/_0819_ ),
    .A2(\hash/_0820_ ),
    .B1(\hash/_0821_ ),
    .Y(\hash/_0822_ ));
 sky130_fd_sc_hd__inv_1 \hash/_3653_  (.A(\hash/_1722_ ),
    .Y(\hash/_0823_ ));
 sky130_fd_sc_hd__nor2_1 \hash/_3654_  (.A(\hash/_1720_ ),
    .B(\hash/_1721_ ),
    .Y(\hash/_0824_ ));
 sky130_fd_sc_hd__o21ai_0 \hash/_3655_  (.A1(\hash/_0823_ ),
    .A2(\hash/_0819_ ),
    .B1(\hash/_0824_ ),
    .Y(\hash/_0825_ ));
 sky130_fd_sc_hd__nor2b_1 \hash/_3656_  (.A(\hash/_0822_ ),
    .B_N(\hash/_0825_ ),
    .Y(\hash/_0143_ ));
 sky130_fd_sc_hd__a21o_1 \hash/_3657_  (.A1(\hash/_1470_ ),
    .A2(\hash/_1722_ ),
    .B1(\hash/_1721_ ),
    .X(\hash/_0826_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3658_  (.A(\hash/a[1] ),
    .B(_09577_),
    .CIN(\hash/_1461_ ),
    .COUT(\hash/_1462_ ),
    .SUM(\hash/_1446_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3659_  (.A(\hash/b[1] ),
    .B(_09578_),
    .CIN(\hash/_1463_ ),
    .COUT(\hash/_1464_ ),
    .SUM(\hash/_1448_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3660_  (.A(\hash/c[1] ),
    .B(_09577_),
    .CIN(\hash/_1465_ ),
    .COUT(\hash/_1466_ ),
    .SUM(\hash/_1450_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3661_  (.A(\hash/d[1] ),
    .B(_09577_),
    .CIN(\hash/_1467_ ),
    .COUT(\hash/_1468_ ),
    .SUM(\hash/_1452_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3662_  (.A(\hash/e[1] ),
    .B(_09577_),
    .CIN(\hash/_1469_ ),
    .COUT(\hash/_1470_ ),
    .SUM(\hash/_1454_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3663_  (.A(\hash/f[1] ),
    .B(_09578_),
    .CIN(\hash/_1471_ ),
    .COUT(\hash/_1472_ ),
    .SUM(\hash/_1456_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3664_  (.A(\hash/g[1] ),
    .B(_09577_),
    .CIN(\hash/_1473_ ),
    .COUT(\hash/_1474_ ),
    .SUM(\hash/_1458_ ));
 sky130_fd_sc_hd__fa_1 \hash/_3665_  (.A(\hash/h[1] ),
    .B(_09578_),
    .CIN(\hash/_1475_ ),
    .COUT(\hash/_1476_ ),
    .SUM(\hash/_1460_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3666_  (.A(\hash/a[0] ),
    .B(_09577_),
    .COUT(\hash/_1461_ ),
    .SUM(\hash/_1445_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3667_  (.A(\hash/a[1] ),
    .B(_09577_),
    .COUT(\hash/_1477_ ),
    .SUM(\hash/_1478_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3668_  (.A(\hash/a[3] ),
    .B(_09578_),
    .COUT(\hash/_1479_ ),
    .SUM(\hash/_1480_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3669_  (.A(\hash/a[2] ),
    .B(_09577_),
    .COUT(\hash/_1481_ ),
    .SUM(\hash/_1482_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3670_  (.A(\hash/a[4] ),
    .B(_09578_),
    .COUT(\hash/_1483_ ),
    .SUM(\hash/_1484_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3671_  (.A(\hash/a[5] ),
    .B(_09577_),
    .COUT(\hash/_1485_ ),
    .SUM(\hash/_1486_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3672_  (.A(\hash/a[6] ),
    .B(_09577_),
    .COUT(\hash/_1487_ ),
    .SUM(\hash/_1488_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3673_  (.A(\hash/a[7] ),
    .B(_09578_),
    .COUT(\hash/_1489_ ),
    .SUM(\hash/_1490_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3674_  (.A(\hash/a[8] ),
    .B(_09578_),
    .COUT(\hash/_1491_ ),
    .SUM(\hash/_1492_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3675_  (.A(\hash/a[9] ),
    .B(_09577_),
    .COUT(\hash/_1493_ ),
    .SUM(\hash/_1494_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3676_  (.A(\hash/a[10] ),
    .B(_09577_),
    .COUT(\hash/_1495_ ),
    .SUM(\hash/_1496_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3677_  (.A(\hash/a[11] ),
    .B(_09578_),
    .COUT(\hash/_1497_ ),
    .SUM(\hash/_1498_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3678_  (.A(\hash/a[12] ),
    .B(_09578_),
    .COUT(\hash/_1499_ ),
    .SUM(\hash/_1500_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3679_  (.A(\hash/a[13] ),
    .B(_09577_),
    .COUT(\hash/_1501_ ),
    .SUM(\hash/_1502_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3680_  (.A(\hash/a[14] ),
    .B(_09577_),
    .COUT(\hash/_1503_ ),
    .SUM(\hash/_1504_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3681_  (.A(\hash/a[16] ),
    .B(_09577_),
    .COUT(\hash/_1505_ ),
    .SUM(\hash/_1506_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3682_  (.A(\hash/a[15] ),
    .B(_09577_),
    .COUT(\hash/_1507_ ),
    .SUM(\hash/_1508_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3683_  (.A(\hash/a[17] ),
    .B(_09578_),
    .COUT(\hash/_1509_ ),
    .SUM(\hash/_1510_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3684_  (.A(\hash/a[18] ),
    .B(_09578_),
    .COUT(\hash/_1511_ ),
    .SUM(\hash/_1512_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3685_  (.A(\hash/a[19] ),
    .B(_09577_),
    .COUT(\hash/_1513_ ),
    .SUM(\hash/_1514_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3686_  (.A(\hash/a[20] ),
    .B(_09578_),
    .COUT(\hash/_1515_ ),
    .SUM(\hash/_1516_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3687_  (.A(\hash/a[21] ),
    .B(_09578_),
    .COUT(\hash/_1517_ ),
    .SUM(\hash/_1518_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3688_  (.A(\hash/a[22] ),
    .B(_09578_),
    .COUT(\hash/_1519_ ),
    .SUM(\hash/_1520_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3689_  (.A(\hash/a[23] ),
    .B(_09578_),
    .COUT(\hash/_1521_ ),
    .SUM(\hash/_1522_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3690_  (.A(\hash/a[24] ),
    .B(_09578_),
    .COUT(\hash/_1523_ ),
    .SUM(\hash/_1524_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3691_  (.A(\hash/a[25] ),
    .B(_09577_),
    .COUT(\hash/_1525_ ),
    .SUM(\hash/_1526_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3692_  (.A(\hash/a[26] ),
    .B(_09578_),
    .COUT(\hash/_1527_ ),
    .SUM(\hash/_1528_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3693_  (.A(\hash/a[27] ),
    .B(_09577_),
    .COUT(\hash/_1529_ ),
    .SUM(\hash/_1530_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3694_  (.A(\hash/a[28] ),
    .B(_09578_),
    .COUT(\hash/_1531_ ),
    .SUM(\hash/_1532_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3695_  (.A(\hash/a[29] ),
    .B(_09577_),
    .COUT(\hash/_1533_ ),
    .SUM(\hash/_1534_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3696_  (.A(\hash/a[30] ),
    .B(_09577_),
    .COUT(\hash/_1535_ ),
    .SUM(\hash/_1536_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3697_  (.A(\hash/b[0] ),
    .B(_09577_),
    .COUT(\hash/_1463_ ),
    .SUM(\hash/_1447_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3698_  (.A(\hash/b[1] ),
    .B(_09578_),
    .COUT(\hash/_1537_ ),
    .SUM(\hash/_1538_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3699_  (.A(\hash/b[3] ),
    .B(_09578_),
    .COUT(\hash/_1539_ ),
    .SUM(\hash/_1540_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3700_  (.A(\hash/b[2] ),
    .B(_09577_),
    .COUT(\hash/_1541_ ),
    .SUM(\hash/_1542_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3701_  (.A(\hash/b[4] ),
    .B(_09578_),
    .COUT(\hash/_1543_ ),
    .SUM(\hash/_1544_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3702_  (.A(\hash/b[5] ),
    .B(_09578_),
    .COUT(\hash/_1545_ ),
    .SUM(\hash/_1546_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3703_  (.A(\hash/b[6] ),
    .B(_09578_),
    .COUT(\hash/_1547_ ),
    .SUM(\hash/_1548_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3704_  (.A(\hash/b[7] ),
    .B(_09577_),
    .COUT(\hash/_1549_ ),
    .SUM(\hash/_1550_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3705_  (.A(\hash/b[8] ),
    .B(_09578_),
    .COUT(\hash/_1551_ ),
    .SUM(\hash/_1552_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3706_  (.A(\hash/b[9] ),
    .B(_09577_),
    .COUT(\hash/_1553_ ),
    .SUM(\hash/_1554_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3707_  (.A(\hash/b[10] ),
    .B(_09577_),
    .COUT(\hash/_1555_ ),
    .SUM(\hash/_1556_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3708_  (.A(\hash/b[11] ),
    .B(_09577_),
    .COUT(\hash/_1557_ ),
    .SUM(\hash/_1558_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3709_  (.A(\hash/b[12] ),
    .B(_09578_),
    .COUT(\hash/_1559_ ),
    .SUM(\hash/_1560_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3710_  (.A(\hash/b[13] ),
    .B(_09577_),
    .COUT(\hash/_1561_ ),
    .SUM(\hash/_1562_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3711_  (.A(\hash/b[14] ),
    .B(_09578_),
    .COUT(\hash/_1563_ ),
    .SUM(\hash/_1564_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3712_  (.A(\hash/b[16] ),
    .B(_09577_),
    .COUT(\hash/_1565_ ),
    .SUM(\hash/_1566_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3713_  (.A(\hash/b[15] ),
    .B(_09577_),
    .COUT(\hash/_1567_ ),
    .SUM(\hash/_1568_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3714_  (.A(\hash/b[17] ),
    .B(_09577_),
    .COUT(\hash/_1569_ ),
    .SUM(\hash/_1570_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3715_  (.A(\hash/b[18] ),
    .B(_09577_),
    .COUT(\hash/_1571_ ),
    .SUM(\hash/_1572_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3716_  (.A(\hash/b[19] ),
    .B(_09578_),
    .COUT(\hash/_1573_ ),
    .SUM(\hash/_1574_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3717_  (.A(\hash/b[20] ),
    .B(_09578_),
    .COUT(\hash/_1575_ ),
    .SUM(\hash/_1576_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3718_  (.A(\hash/b[21] ),
    .B(_09577_),
    .COUT(\hash/_1577_ ),
    .SUM(\hash/_1578_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3719_  (.A(\hash/b[22] ),
    .B(_09577_),
    .COUT(\hash/_1579_ ),
    .SUM(\hash/_1580_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3720_  (.A(\hash/b[23] ),
    .B(_09578_),
    .COUT(\hash/_1581_ ),
    .SUM(\hash/_1582_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3721_  (.A(\hash/b[24] ),
    .B(_09577_),
    .COUT(\hash/_1583_ ),
    .SUM(\hash/_1584_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3722_  (.A(\hash/b[25] ),
    .B(_09577_),
    .COUT(\hash/_1585_ ),
    .SUM(\hash/_1586_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3723_  (.A(\hash/b[26] ),
    .B(_09578_),
    .COUT(\hash/_1587_ ),
    .SUM(\hash/_1588_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3724_  (.A(\hash/b[27] ),
    .B(_09577_),
    .COUT(\hash/_1589_ ),
    .SUM(\hash/_1590_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3725_  (.A(\hash/b[28] ),
    .B(_09577_),
    .COUT(\hash/_1591_ ),
    .SUM(\hash/_1592_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3726_  (.A(\hash/b[29] ),
    .B(_09577_),
    .COUT(\hash/_1593_ ),
    .SUM(\hash/_1594_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3727_  (.A(\hash/b[30] ),
    .B(_09578_),
    .COUT(\hash/_1595_ ),
    .SUM(\hash/_1596_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3728_  (.A(\hash/c[0] ),
    .B(_09578_),
    .COUT(\hash/_1465_ ),
    .SUM(\hash/_1449_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3729_  (.A(\hash/c[1] ),
    .B(_09577_),
    .COUT(\hash/_1597_ ),
    .SUM(\hash/_1598_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3730_  (.A(\hash/c[3] ),
    .B(_09578_),
    .COUT(\hash/_1599_ ),
    .SUM(\hash/_1600_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3731_  (.A(\hash/c[2] ),
    .B(_09578_),
    .COUT(\hash/_1601_ ),
    .SUM(\hash/_1602_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3732_  (.A(\hash/c[4] ),
    .B(_09577_),
    .COUT(\hash/_1603_ ),
    .SUM(\hash/_1604_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3733_  (.A(\hash/c[5] ),
    .B(_09577_),
    .COUT(\hash/_1605_ ),
    .SUM(\hash/_1606_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3734_  (.A(\hash/c[6] ),
    .B(_09577_),
    .COUT(\hash/_1607_ ),
    .SUM(\hash/_1608_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3735_  (.A(\hash/c[7] ),
    .B(_09578_),
    .COUT(\hash/_1609_ ),
    .SUM(\hash/_1610_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3736_  (.A(\hash/c[8] ),
    .B(_09577_),
    .COUT(\hash/_1611_ ),
    .SUM(\hash/_1612_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3737_  (.A(\hash/c[9] ),
    .B(_09577_),
    .COUT(\hash/_1613_ ),
    .SUM(\hash/_1614_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3738_  (.A(\hash/c[10] ),
    .B(_09578_),
    .COUT(\hash/_1615_ ),
    .SUM(\hash/_1616_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3739_  (.A(\hash/c[11] ),
    .B(_09578_),
    .COUT(\hash/_1617_ ),
    .SUM(\hash/_1618_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3740_  (.A(\hash/c[12] ),
    .B(_09577_),
    .COUT(\hash/_1619_ ),
    .SUM(\hash/_1620_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3741_  (.A(\hash/c[13] ),
    .B(_09577_),
    .COUT(\hash/_1621_ ),
    .SUM(\hash/_1622_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3742_  (.A(\hash/c[14] ),
    .B(_09577_),
    .COUT(\hash/_1623_ ),
    .SUM(\hash/_1624_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3743_  (.A(\hash/c[16] ),
    .B(_09578_),
    .COUT(\hash/_1625_ ),
    .SUM(\hash/_1626_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3744_  (.A(\hash/c[15] ),
    .B(_09577_),
    .COUT(\hash/_1627_ ),
    .SUM(\hash/_1628_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3745_  (.A(\hash/c[17] ),
    .B(_09577_),
    .COUT(\hash/_1629_ ),
    .SUM(\hash/_1630_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3746_  (.A(\hash/c[18] ),
    .B(_09577_),
    .COUT(\hash/_1631_ ),
    .SUM(\hash/_1632_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3747_  (.A(\hash/c[19] ),
    .B(_09577_),
    .COUT(\hash/_1633_ ),
    .SUM(\hash/_1634_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3748_  (.A(\hash/c[20] ),
    .B(_09578_),
    .COUT(\hash/_1635_ ),
    .SUM(\hash/_1636_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3749_  (.A(\hash/c[21] ),
    .B(_09577_),
    .COUT(\hash/_1637_ ),
    .SUM(\hash/_1638_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3750_  (.A(\hash/c[22] ),
    .B(_09577_),
    .COUT(\hash/_1639_ ),
    .SUM(\hash/_1640_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3751_  (.A(\hash/c[23] ),
    .B(_09578_),
    .COUT(\hash/_1641_ ),
    .SUM(\hash/_1642_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3752_  (.A(\hash/c[24] ),
    .B(_09578_),
    .COUT(\hash/_1643_ ),
    .SUM(\hash/_1644_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3753_  (.A(\hash/c[25] ),
    .B(_09578_),
    .COUT(\hash/_1645_ ),
    .SUM(\hash/_1646_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3754_  (.A(\hash/c[26] ),
    .B(_09577_),
    .COUT(\hash/_1647_ ),
    .SUM(\hash/_1648_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3755_  (.A(\hash/c[27] ),
    .B(_09577_),
    .COUT(\hash/_1649_ ),
    .SUM(\hash/_1650_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3756_  (.A(\hash/c[28] ),
    .B(_09577_),
    .COUT(\hash/_1651_ ),
    .SUM(\hash/_1652_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3757_  (.A(\hash/c[29] ),
    .B(_09577_),
    .COUT(\hash/_1653_ ),
    .SUM(\hash/_1654_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3758_  (.A(\hash/c[30] ),
    .B(_09578_),
    .COUT(\hash/_1655_ ),
    .SUM(\hash/_1656_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3759_  (.A(\hash/d[0] ),
    .B(_09578_),
    .COUT(\hash/_1467_ ),
    .SUM(\hash/_1451_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3760_  (.A(\hash/d[1] ),
    .B(_09577_),
    .COUT(\hash/_1657_ ),
    .SUM(\hash/_1658_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3761_  (.A(\hash/d[3] ),
    .B(_09577_),
    .COUT(\hash/_1659_ ),
    .SUM(\hash/_1660_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3762_  (.A(\hash/d[2] ),
    .B(_09578_),
    .COUT(\hash/_1661_ ),
    .SUM(\hash/_1662_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3763_  (.A(\hash/d[4] ),
    .B(_09577_),
    .COUT(\hash/_1663_ ),
    .SUM(\hash/_1664_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3764_  (.A(\hash/d[5] ),
    .B(_09577_),
    .COUT(\hash/_1665_ ),
    .SUM(\hash/_1666_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3765_  (.A(\hash/d[6] ),
    .B(_09578_),
    .COUT(\hash/_1667_ ),
    .SUM(\hash/_1668_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3766_  (.A(\hash/d[7] ),
    .B(_09578_),
    .COUT(\hash/_1669_ ),
    .SUM(\hash/_1670_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3767_  (.A(\hash/d[8] ),
    .B(_09577_),
    .COUT(\hash/_1671_ ),
    .SUM(\hash/_1672_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3768_  (.A(\hash/d[9] ),
    .B(_09578_),
    .COUT(\hash/_1673_ ),
    .SUM(\hash/_1674_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3769_  (.A(\hash/d[10] ),
    .B(_09577_),
    .COUT(\hash/_1675_ ),
    .SUM(\hash/_1676_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3770_  (.A(\hash/d[11] ),
    .B(_09578_),
    .COUT(\hash/_1677_ ),
    .SUM(\hash/_1678_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3771_  (.A(\hash/d[12] ),
    .B(_09577_),
    .COUT(\hash/_1679_ ),
    .SUM(\hash/_1680_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3772_  (.A(\hash/d[13] ),
    .B(_09577_),
    .COUT(\hash/_1681_ ),
    .SUM(\hash/_1682_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3773_  (.A(\hash/d[14] ),
    .B(_09577_),
    .COUT(\hash/_1683_ ),
    .SUM(\hash/_1684_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3774_  (.A(\hash/d[16] ),
    .B(_09577_),
    .COUT(\hash/_1685_ ),
    .SUM(\hash/_1686_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3775_  (.A(\hash/d[15] ),
    .B(_09577_),
    .COUT(\hash/_1687_ ),
    .SUM(\hash/_1688_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3776_  (.A(\hash/d[17] ),
    .B(_09577_),
    .COUT(\hash/_1689_ ),
    .SUM(\hash/_1690_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3777_  (.A(\hash/d[18] ),
    .B(_09577_),
    .COUT(\hash/_1691_ ),
    .SUM(\hash/_1692_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3778_  (.A(\hash/d[19] ),
    .B(_09577_),
    .COUT(\hash/_1693_ ),
    .SUM(\hash/_1694_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3779_  (.A(\hash/d[20] ),
    .B(_09578_),
    .COUT(\hash/_1695_ ),
    .SUM(\hash/_1696_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3780_  (.A(\hash/d[21] ),
    .B(_09578_),
    .COUT(\hash/_1697_ ),
    .SUM(\hash/_1698_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3781_  (.A(\hash/d[22] ),
    .B(_09577_),
    .COUT(\hash/_1699_ ),
    .SUM(\hash/_1700_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3782_  (.A(\hash/d[23] ),
    .B(_09578_),
    .COUT(\hash/_1701_ ),
    .SUM(\hash/_1702_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3783_  (.A(\hash/d[24] ),
    .B(_09577_),
    .COUT(\hash/_1703_ ),
    .SUM(\hash/_1704_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3784_  (.A(\hash/d[25] ),
    .B(_09578_),
    .COUT(\hash/_1705_ ),
    .SUM(\hash/_1706_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3785_  (.A(\hash/d[26] ),
    .B(_09577_),
    .COUT(\hash/_1707_ ),
    .SUM(\hash/_1708_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3786_  (.A(\hash/d[27] ),
    .B(_09578_),
    .COUT(\hash/_1709_ ),
    .SUM(\hash/_1710_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3787_  (.A(\hash/d[28] ),
    .B(_09578_),
    .COUT(\hash/_1711_ ),
    .SUM(\hash/_1712_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3788_  (.A(\hash/d[29] ),
    .B(_09577_),
    .COUT(\hash/_1713_ ),
    .SUM(\hash/_1714_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3789_  (.A(\hash/d[30] ),
    .B(_09578_),
    .COUT(\hash/_1715_ ),
    .SUM(\hash/_1716_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3790_  (.A(\hash/e[0] ),
    .B(_09577_),
    .COUT(\hash/_1469_ ),
    .SUM(\hash/_1453_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3791_  (.A(\hash/e[1] ),
    .B(_09577_),
    .COUT(\hash/_1717_ ),
    .SUM(\hash/_1718_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3792_  (.A(\hash/e[3] ),
    .B(_09577_),
    .COUT(\hash/_1719_ ),
    .SUM(\hash/_1720_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3793_  (.A(\hash/e[2] ),
    .B(_09577_),
    .COUT(\hash/_1721_ ),
    .SUM(\hash/_1722_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3794_  (.A(\hash/e[4] ),
    .B(_09577_),
    .COUT(\hash/_1723_ ),
    .SUM(\hash/_1724_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3795_  (.A(\hash/e[5] ),
    .B(_09577_),
    .COUT(\hash/_1725_ ),
    .SUM(\hash/_1726_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3796_  (.A(\hash/e[6] ),
    .B(_09577_),
    .COUT(\hash/_1727_ ),
    .SUM(\hash/_1728_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3797_  (.A(\hash/e[7] ),
    .B(_09578_),
    .COUT(\hash/_1729_ ),
    .SUM(\hash/_1730_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3798_  (.A(\hash/e[8] ),
    .B(_09578_),
    .COUT(\hash/_1731_ ),
    .SUM(\hash/_1732_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3799_  (.A(\hash/e[9] ),
    .B(_09577_),
    .COUT(\hash/_1733_ ),
    .SUM(\hash/_1734_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3800_  (.A(\hash/e[10] ),
    .B(_09578_),
    .COUT(\hash/_1735_ ),
    .SUM(\hash/_1736_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3801_  (.A(\hash/e[11] ),
    .B(_09578_),
    .COUT(\hash/_1737_ ),
    .SUM(\hash/_1738_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3802_  (.A(\hash/e[12] ),
    .B(_09577_),
    .COUT(\hash/_1739_ ),
    .SUM(\hash/_1740_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3803_  (.A(\hash/e[13] ),
    .B(_09578_),
    .COUT(\hash/_1741_ ),
    .SUM(\hash/_1742_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3804_  (.A(\hash/e[14] ),
    .B(_09577_),
    .COUT(\hash/_1743_ ),
    .SUM(\hash/_1744_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3805_  (.A(\hash/e[16] ),
    .B(_09578_),
    .COUT(\hash/_1745_ ),
    .SUM(\hash/_1746_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3806_  (.A(\hash/e[15] ),
    .B(_09578_),
    .COUT(\hash/_1747_ ),
    .SUM(\hash/_1748_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3807_  (.A(\hash/e[17] ),
    .B(_09577_),
    .COUT(\hash/_1749_ ),
    .SUM(\hash/_1750_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3808_  (.A(\hash/e[18] ),
    .B(_09577_),
    .COUT(\hash/_1751_ ),
    .SUM(\hash/_1752_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3809_  (.A(\hash/e[19] ),
    .B(_09577_),
    .COUT(\hash/_1753_ ),
    .SUM(\hash/_1754_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3810_  (.A(\hash/e[20] ),
    .B(_09578_),
    .COUT(\hash/_1755_ ),
    .SUM(\hash/_1756_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3811_  (.A(\hash/e[21] ),
    .B(_09578_),
    .COUT(\hash/_1757_ ),
    .SUM(\hash/_1758_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3812_  (.A(\hash/e[22] ),
    .B(_09578_),
    .COUT(\hash/_1759_ ),
    .SUM(\hash/_1760_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3813_  (.A(\hash/e[23] ),
    .B(_09578_),
    .COUT(\hash/_1761_ ),
    .SUM(\hash/_1762_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3814_  (.A(\hash/e[24] ),
    .B(_09577_),
    .COUT(\hash/_1763_ ),
    .SUM(\hash/_1764_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3815_  (.A(\hash/e[25] ),
    .B(_09578_),
    .COUT(\hash/_1765_ ),
    .SUM(\hash/_1766_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3816_  (.A(\hash/e[26] ),
    .B(_09578_),
    .COUT(\hash/_1767_ ),
    .SUM(\hash/_1768_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3817_  (.A(\hash/e[27] ),
    .B(_09578_),
    .COUT(\hash/_1769_ ),
    .SUM(\hash/_1770_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3818_  (.A(\hash/e[28] ),
    .B(_09577_),
    .COUT(\hash/_1771_ ),
    .SUM(\hash/_1772_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3819_  (.A(\hash/e[29] ),
    .B(_09578_),
    .COUT(\hash/_1773_ ),
    .SUM(\hash/_1774_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3820_  (.A(\hash/e[30] ),
    .B(_09577_),
    .COUT(\hash/_1775_ ),
    .SUM(\hash/_1776_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3821_  (.A(\hash/f[0] ),
    .B(_09578_),
    .COUT(\hash/_1471_ ),
    .SUM(\hash/_1455_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3822_  (.A(\hash/f[1] ),
    .B(_09578_),
    .COUT(\hash/_1777_ ),
    .SUM(\hash/_1778_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3823_  (.A(\hash/f[3] ),
    .B(_09577_),
    .COUT(\hash/_1779_ ),
    .SUM(\hash/_1780_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3824_  (.A(\hash/f[2] ),
    .B(_09577_),
    .COUT(\hash/_1781_ ),
    .SUM(\hash/_1782_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3825_  (.A(\hash/f[4] ),
    .B(_09578_),
    .COUT(\hash/_1783_ ),
    .SUM(\hash/_1784_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3826_  (.A(\hash/f[5] ),
    .B(_09578_),
    .COUT(\hash/_1785_ ),
    .SUM(\hash/_1786_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3827_  (.A(\hash/f[6] ),
    .B(_09578_),
    .COUT(\hash/_1787_ ),
    .SUM(\hash/_1788_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3828_  (.A(\hash/f[7] ),
    .B(_09577_),
    .COUT(\hash/_1789_ ),
    .SUM(\hash/_1790_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3829_  (.A(\hash/f[8] ),
    .B(_09578_),
    .COUT(\hash/_1791_ ),
    .SUM(\hash/_1792_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3830_  (.A(\hash/f[9] ),
    .B(_09578_),
    .COUT(\hash/_1793_ ),
    .SUM(\hash/_1794_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3831_  (.A(\hash/f[10] ),
    .B(_09578_),
    .COUT(\hash/_1795_ ),
    .SUM(\hash/_1796_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3832_  (.A(\hash/f[11] ),
    .B(_09577_),
    .COUT(\hash/_1797_ ),
    .SUM(\hash/_1798_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3833_  (.A(\hash/f[12] ),
    .B(_09578_),
    .COUT(\hash/_1799_ ),
    .SUM(\hash/_1800_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3834_  (.A(\hash/f[13] ),
    .B(_09577_),
    .COUT(\hash/_1801_ ),
    .SUM(\hash/_1802_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3835_  (.A(\hash/f[14] ),
    .B(_09577_),
    .COUT(\hash/_1803_ ),
    .SUM(\hash/_1804_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3836_  (.A(\hash/f[16] ),
    .B(_09577_),
    .COUT(\hash/_1805_ ),
    .SUM(\hash/_1806_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3837_  (.A(\hash/f[15] ),
    .B(_09578_),
    .COUT(\hash/_1807_ ),
    .SUM(\hash/_1808_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3838_  (.A(\hash/f[17] ),
    .B(_09578_),
    .COUT(\hash/_1809_ ),
    .SUM(\hash/_1810_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3839_  (.A(\hash/f[18] ),
    .B(_09577_),
    .COUT(\hash/_1811_ ),
    .SUM(\hash/_1812_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3840_  (.A(\hash/f[19] ),
    .B(_09578_),
    .COUT(\hash/_1813_ ),
    .SUM(\hash/_1814_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3841_  (.A(\hash/f[20] ),
    .B(_09578_),
    .COUT(\hash/_1815_ ),
    .SUM(\hash/_1816_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3842_  (.A(\hash/f[21] ),
    .B(_09578_),
    .COUT(\hash/_1817_ ),
    .SUM(\hash/_1818_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3843_  (.A(\hash/f[22] ),
    .B(_09578_),
    .COUT(\hash/_1819_ ),
    .SUM(\hash/_1820_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3844_  (.A(\hash/f[23] ),
    .B(_09578_),
    .COUT(\hash/_1821_ ),
    .SUM(\hash/_1822_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3845_  (.A(\hash/f[24] ),
    .B(_09577_),
    .COUT(\hash/_1823_ ),
    .SUM(\hash/_1824_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3846_  (.A(\hash/f[25] ),
    .B(_09577_),
    .COUT(\hash/_1825_ ),
    .SUM(\hash/_1826_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3847_  (.A(\hash/f[26] ),
    .B(_09578_),
    .COUT(\hash/_1827_ ),
    .SUM(\hash/_1828_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3848_  (.A(\hash/f[27] ),
    .B(_09577_),
    .COUT(\hash/_1829_ ),
    .SUM(\hash/_1830_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3849_  (.A(\hash/f[28] ),
    .B(_09577_),
    .COUT(\hash/_1831_ ),
    .SUM(\hash/_1832_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3850_  (.A(\hash/f[29] ),
    .B(_09578_),
    .COUT(\hash/_1833_ ),
    .SUM(\hash/_1834_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3851_  (.A(\hash/f[30] ),
    .B(_09578_),
    .COUT(\hash/_1835_ ),
    .SUM(\hash/_1836_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3852_  (.A(\hash/g[0] ),
    .B(_09577_),
    .COUT(\hash/_1473_ ),
    .SUM(\hash/_1457_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3853_  (.A(\hash/g[1] ),
    .B(_09577_),
    .COUT(\hash/_1837_ ),
    .SUM(\hash/_1838_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3854_  (.A(\hash/g[3] ),
    .B(_09577_),
    .COUT(\hash/_1839_ ),
    .SUM(\hash/_1840_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3855_  (.A(\hash/g[2] ),
    .B(_09578_),
    .COUT(\hash/_1841_ ),
    .SUM(\hash/_1842_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3856_  (.A(\hash/g[4] ),
    .B(_09578_),
    .COUT(\hash/_1843_ ),
    .SUM(\hash/_1844_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3857_  (.A(\hash/g[5] ),
    .B(_09577_),
    .COUT(\hash/_1845_ ),
    .SUM(\hash/_1846_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3858_  (.A(\hash/g[6] ),
    .B(_09578_),
    .COUT(\hash/_1847_ ),
    .SUM(\hash/_1848_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3859_  (.A(\hash/g[7] ),
    .B(_09577_),
    .COUT(\hash/_1849_ ),
    .SUM(\hash/_1850_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3860_  (.A(\hash/g[8] ),
    .B(_09577_),
    .COUT(\hash/_1851_ ),
    .SUM(\hash/_1852_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3861_  (.A(\hash/g[9] ),
    .B(_09578_),
    .COUT(\hash/_1853_ ),
    .SUM(\hash/_1854_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3862_  (.A(\hash/g[10] ),
    .B(_09578_),
    .COUT(\hash/_1855_ ),
    .SUM(\hash/_1856_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3863_  (.A(\hash/g[11] ),
    .B(_09577_),
    .COUT(\hash/_1857_ ),
    .SUM(\hash/_1858_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3864_  (.A(\hash/g[12] ),
    .B(_09577_),
    .COUT(\hash/_1859_ ),
    .SUM(\hash/_1860_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3865_  (.A(\hash/g[13] ),
    .B(_09578_),
    .COUT(\hash/_1861_ ),
    .SUM(\hash/_1862_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3866_  (.A(\hash/g[14] ),
    .B(_09577_),
    .COUT(\hash/_1863_ ),
    .SUM(\hash/_1864_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3867_  (.A(\hash/g[16] ),
    .B(_09577_),
    .COUT(\hash/_1865_ ),
    .SUM(\hash/_1866_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3868_  (.A(\hash/g[15] ),
    .B(_09577_),
    .COUT(\hash/_1867_ ),
    .SUM(\hash/_1868_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3869_  (.A(\hash/g[17] ),
    .B(_09577_),
    .COUT(\hash/_1869_ ),
    .SUM(\hash/_1870_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3870_  (.A(\hash/g[18] ),
    .B(_09578_),
    .COUT(\hash/_1871_ ),
    .SUM(\hash/_1872_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3871_  (.A(\hash/g[19] ),
    .B(_09578_),
    .COUT(\hash/_1873_ ),
    .SUM(\hash/_1874_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3872_  (.A(\hash/g[20] ),
    .B(_09578_),
    .COUT(\hash/_1875_ ),
    .SUM(\hash/_1876_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3873_  (.A(\hash/g[21] ),
    .B(_09578_),
    .COUT(\hash/_1877_ ),
    .SUM(\hash/_1878_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3874_  (.A(\hash/g[22] ),
    .B(_09578_),
    .COUT(\hash/_1879_ ),
    .SUM(\hash/_1880_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3875_  (.A(\hash/g[23] ),
    .B(_09577_),
    .COUT(\hash/_1881_ ),
    .SUM(\hash/_1882_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3876_  (.A(\hash/g[24] ),
    .B(_09577_),
    .COUT(\hash/_1883_ ),
    .SUM(\hash/_1884_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3877_  (.A(\hash/g[25] ),
    .B(_09577_),
    .COUT(\hash/_1885_ ),
    .SUM(\hash/_1886_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3878_  (.A(\hash/g[26] ),
    .B(_09577_),
    .COUT(\hash/_1887_ ),
    .SUM(\hash/_1888_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3879_  (.A(\hash/g[27] ),
    .B(_09577_),
    .COUT(\hash/_1889_ ),
    .SUM(\hash/_1890_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3880_  (.A(\hash/g[28] ),
    .B(_09577_),
    .COUT(\hash/_1891_ ),
    .SUM(\hash/_1892_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3881_  (.A(\hash/g[29] ),
    .B(_09578_),
    .COUT(\hash/_1893_ ),
    .SUM(\hash/_1894_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3882_  (.A(\hash/g[30] ),
    .B(_09578_),
    .COUT(\hash/_1895_ ),
    .SUM(\hash/_1896_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3883_  (.A(\hash/h[0] ),
    .B(_09577_),
    .COUT(\hash/_1475_ ),
    .SUM(\hash/_1459_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3884_  (.A(\hash/h[1] ),
    .B(_09578_),
    .COUT(\hash/_1897_ ),
    .SUM(\hash/_1898_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3885_  (.A(\hash/h[3] ),
    .B(_09577_),
    .COUT(\hash/_1899_ ),
    .SUM(\hash/_1900_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3886_  (.A(\hash/h[2] ),
    .B(_09578_),
    .COUT(\hash/_1901_ ),
    .SUM(\hash/_1902_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3887_  (.A(\hash/h[4] ),
    .B(_09577_),
    .COUT(\hash/_1903_ ),
    .SUM(\hash/_1904_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3888_  (.A(\hash/h[5] ),
    .B(_09578_),
    .COUT(\hash/_1905_ ),
    .SUM(\hash/_1906_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3889_  (.A(\hash/h[6] ),
    .B(_09578_),
    .COUT(\hash/_1907_ ),
    .SUM(\hash/_1908_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3890_  (.A(\hash/h[7] ),
    .B(_09578_),
    .COUT(\hash/_1909_ ),
    .SUM(\hash/_1910_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3891_  (.A(\hash/h[8] ),
    .B(_09577_),
    .COUT(\hash/_1911_ ),
    .SUM(\hash/_1912_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3892_  (.A(\hash/h[9] ),
    .B(_09578_),
    .COUT(\hash/_1913_ ),
    .SUM(\hash/_1914_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3893_  (.A(\hash/h[10] ),
    .B(_09577_),
    .COUT(\hash/_1915_ ),
    .SUM(\hash/_1916_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3894_  (.A(\hash/h[11] ),
    .B(_09577_),
    .COUT(\hash/_1917_ ),
    .SUM(\hash/_1918_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3895_  (.A(\hash/h[12] ),
    .B(_09578_),
    .COUT(\hash/_1919_ ),
    .SUM(\hash/_1920_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3896_  (.A(\hash/h[13] ),
    .B(_09578_),
    .COUT(\hash/_1921_ ),
    .SUM(\hash/_1922_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3897_  (.A(\hash/h[14] ),
    .B(_09577_),
    .COUT(\hash/_1923_ ),
    .SUM(\hash/_1924_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3898_  (.A(\hash/h[16] ),
    .B(_09578_),
    .COUT(\hash/_1925_ ),
    .SUM(\hash/_1926_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3899_  (.A(\hash/h[15] ),
    .B(_09577_),
    .COUT(\hash/_1927_ ),
    .SUM(\hash/_1928_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3900_  (.A(\hash/h[17] ),
    .B(_09578_),
    .COUT(\hash/_1929_ ),
    .SUM(\hash/_1930_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3901_  (.A(\hash/h[18] ),
    .B(_09578_),
    .COUT(\hash/_1931_ ),
    .SUM(\hash/_1932_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3902_  (.A(\hash/h[19] ),
    .B(_09578_),
    .COUT(\hash/_1933_ ),
    .SUM(\hash/_1934_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3903_  (.A(\hash/h[20] ),
    .B(_09578_),
    .COUT(\hash/_1935_ ),
    .SUM(\hash/_1936_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3904_  (.A(\hash/h[21] ),
    .B(_09577_),
    .COUT(\hash/_1937_ ),
    .SUM(\hash/_1938_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3905_  (.A(\hash/h[22] ),
    .B(_09577_),
    .COUT(\hash/_1939_ ),
    .SUM(\hash/_1940_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3906_  (.A(\hash/h[23] ),
    .B(_09577_),
    .COUT(\hash/_1941_ ),
    .SUM(\hash/_1942_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3907_  (.A(\hash/h[24] ),
    .B(_09577_),
    .COUT(\hash/_1943_ ),
    .SUM(\hash/_1944_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3908_  (.A(\hash/h[25] ),
    .B(_09577_),
    .COUT(\hash/_1945_ ),
    .SUM(\hash/_1946_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3909_  (.A(\hash/h[26] ),
    .B(_09578_),
    .COUT(\hash/_1947_ ),
    .SUM(\hash/_1948_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3910_  (.A(\hash/h[27] ),
    .B(_09577_),
    .COUT(\hash/_1949_ ),
    .SUM(\hash/_1950_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3911_  (.A(\hash/h[28] ),
    .B(_09577_),
    .COUT(\hash/_1951_ ),
    .SUM(\hash/_1952_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3912_  (.A(\hash/h[29] ),
    .B(_09578_),
    .COUT(\hash/_1953_ ),
    .SUM(\hash/_1954_ ));
 sky130_fd_sc_hd__ha_1 \hash/_3913_  (.A(\hash/h[30] ),
    .B(_09577_),
    .COUT(\hash/_1955_ ),
    .SUM(\hash/_1956_ ));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[0]$_DFF_P_  (.D(\hash/a[0] ),
    .Q(\hash/a_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[10]$_DFF_P_  (.D(\hash/a[10] ),
    .Q(\hash/a_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[11]$_DFF_P_  (.D(\hash/a[11] ),
    .Q(\hash/a_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[12]$_DFF_P_  (.D(\hash/a[12] ),
    .Q(\hash/a_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[13]$_DFF_P_  (.D(\hash/a[13] ),
    .Q(\hash/a_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[14]$_DFF_P_  (.D(\hash/a[14] ),
    .Q(\hash/a_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[15]$_DFF_P_  (.D(\hash/a[15] ),
    .Q(\hash/a_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[16]$_DFF_P_  (.D(\hash/a[16] ),
    .Q(\hash/a_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[17]$_DFF_P_  (.D(\hash/a[17] ),
    .Q(\hash/a_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[18]$_DFF_P_  (.D(\hash/a[18] ),
    .Q(\hash/a_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[19]$_DFF_P_  (.D(\hash/a[19] ),
    .Q(\hash/a_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[1]$_DFF_P_  (.D(\hash/a[1] ),
    .Q(\hash/a_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[20]$_DFF_P_  (.D(\hash/a[20] ),
    .Q(\hash/a_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[21]$_DFF_P_  (.D(\hash/a[21] ),
    .Q(\hash/a_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[22]$_DFF_P_  (.D(\hash/a[22] ),
    .Q(\hash/a_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[23]$_DFF_P_  (.D(\hash/a[23] ),
    .Q(\hash/a_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[24]$_DFF_P_  (.D(\hash/a[24] ),
    .Q(\hash/a_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[25]$_DFF_P_  (.D(\hash/a[25] ),
    .Q(\hash/a_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[26]$_DFF_P_  (.D(\hash/a[26] ),
    .Q(\hash/a_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[27]$_DFF_P_  (.D(\hash/a[27] ),
    .Q(\hash/a_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[28]$_DFF_P_  (.D(\hash/a[28] ),
    .Q(\hash/a_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[29]$_DFF_P_  (.D(\hash/a[29] ),
    .Q(\hash/a_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[2]$_DFF_P_  (.D(\hash/a[2] ),
    .Q(\hash/a_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[30]$_DFF_P_  (.D(\hash/a[30] ),
    .Q(\hash/a_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[31]$_DFF_P_  (.D(\hash/a[31] ),
    .Q(\hash/a_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[3]$_DFF_P_  (.D(\hash/a[3] ),
    .Q(\hash/a_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[4]$_DFF_P_  (.D(\hash/a[4] ),
    .Q(\hash/a_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[5]$_DFF_P_  (.D(\hash/a[5] ),
    .Q(\hash/a_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[6]$_DFF_P_  (.D(\hash/a[6] ),
    .Q(\hash/a_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[7]$_DFF_P_  (.D(\hash/a[7] ),
    .Q(\hash/a_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[8]$_DFF_P_  (.D(\hash/a[8] ),
    .Q(\hash/a_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/a_cap[9]$_DFF_P_  (.D(\hash/a[9] ),
    .Q(\hash/a_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[0]$_DFF_P_  (.D(\hash/b[0] ),
    .Q(\hash/b_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[10]$_DFF_P_  (.D(\hash/b[10] ),
    .Q(\hash/b_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[11]$_DFF_P_  (.D(\hash/b[11] ),
    .Q(\hash/b_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[12]$_DFF_P_  (.D(\hash/b[12] ),
    .Q(\hash/b_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[13]$_DFF_P_  (.D(\hash/b[13] ),
    .Q(\hash/b_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[14]$_DFF_P_  (.D(\hash/b[14] ),
    .Q(\hash/b_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[15]$_DFF_P_  (.D(\hash/b[15] ),
    .Q(\hash/b_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[16]$_DFF_P_  (.D(\hash/b[16] ),
    .Q(\hash/b_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[17]$_DFF_P_  (.D(\hash/b[17] ),
    .Q(\hash/b_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[18]$_DFF_P_  (.D(\hash/b[18] ),
    .Q(\hash/b_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[19]$_DFF_P_  (.D(\hash/b[19] ),
    .Q(\hash/b_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[1]$_DFF_P_  (.D(\hash/b[1] ),
    .Q(\hash/b_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[20]$_DFF_P_  (.D(\hash/b[20] ),
    .Q(\hash/b_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[21]$_DFF_P_  (.D(\hash/b[21] ),
    .Q(\hash/b_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[22]$_DFF_P_  (.D(\hash/b[22] ),
    .Q(\hash/b_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[23]$_DFF_P_  (.D(\hash/b[23] ),
    .Q(\hash/b_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[24]$_DFF_P_  (.D(\hash/b[24] ),
    .Q(\hash/b_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[25]$_DFF_P_  (.D(\hash/b[25] ),
    .Q(\hash/b_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[26]$_DFF_P_  (.D(\hash/b[26] ),
    .Q(\hash/b_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[27]$_DFF_P_  (.D(\hash/b[27] ),
    .Q(\hash/b_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[28]$_DFF_P_  (.D(\hash/b[28] ),
    .Q(\hash/b_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[29]$_DFF_P_  (.D(\hash/b[29] ),
    .Q(\hash/b_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[2]$_DFF_P_  (.D(\hash/b[2] ),
    .Q(\hash/b_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[30]$_DFF_P_  (.D(\hash/b[30] ),
    .Q(\hash/b_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[31]$_DFF_P_  (.D(\hash/b[31] ),
    .Q(\hash/b_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[3]$_DFF_P_  (.D(\hash/b[3] ),
    .Q(\hash/b_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[4]$_DFF_P_  (.D(\hash/b[4] ),
    .Q(\hash/b_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[5]$_DFF_P_  (.D(\hash/b[5] ),
    .Q(\hash/b_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[6]$_DFF_P_  (.D(\hash/b[6] ),
    .Q(\hash/b_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[7]$_DFF_P_  (.D(\hash/b[7] ),
    .Q(\hash/b_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[8]$_DFF_P_  (.D(\hash/b[8] ),
    .Q(\hash/b_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/b_cap[9]$_DFF_P_  (.D(\hash/b[9] ),
    .Q(\hash/b_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[0]$_DFF_P_  (.D(\hash/e[0] ),
    .Q(\hash/e_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[10]$_DFF_P_  (.D(\hash/e[10] ),
    .Q(\hash/e_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[11]$_DFF_P_  (.D(\hash/e[11] ),
    .Q(\hash/e_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[12]$_DFF_P_  (.D(\hash/e[12] ),
    .Q(\hash/e_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[13]$_DFF_P_  (.D(\hash/e[13] ),
    .Q(\hash/e_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[14]$_DFF_P_  (.D(\hash/e[14] ),
    .Q(\hash/e_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[15]$_DFF_P_  (.D(\hash/e[15] ),
    .Q(\hash/e_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[16]$_DFF_P_  (.D(\hash/e[16] ),
    .Q(\hash/e_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[17]$_DFF_P_  (.D(\hash/e[17] ),
    .Q(\hash/e_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[18]$_DFF_P_  (.D(\hash/e[18] ),
    .Q(\hash/e_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[19]$_DFF_P_  (.D(\hash/e[19] ),
    .Q(\hash/e_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[1]$_DFF_P_  (.D(\hash/e[1] ),
    .Q(\hash/e_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[20]$_DFF_P_  (.D(\hash/e[20] ),
    .Q(\hash/e_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[21]$_DFF_P_  (.D(\hash/e[21] ),
    .Q(\hash/e_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[22]$_DFF_P_  (.D(\hash/e[22] ),
    .Q(\hash/e_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[23]$_DFF_P_  (.D(\hash/e[23] ),
    .Q(\hash/e_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[24]$_DFF_P_  (.D(\hash/e[24] ),
    .Q(\hash/e_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[25]$_DFF_P_  (.D(\hash/e[25] ),
    .Q(\hash/e_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[26]$_DFF_P_  (.D(\hash/e[26] ),
    .Q(\hash/e_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[27]$_DFF_P_  (.D(\hash/e[27] ),
    .Q(\hash/e_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[28]$_DFF_P_  (.D(\hash/e[28] ),
    .Q(\hash/e_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[29]$_DFF_P_  (.D(\hash/e[29] ),
    .Q(\hash/e_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[2]$_DFF_P_  (.D(\hash/e[2] ),
    .Q(\hash/e_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[30]$_DFF_P_  (.D(\hash/e[30] ),
    .Q(\hash/e_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[31]$_DFF_P_  (.D(\hash/e[31] ),
    .Q(\hash/e_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[3]$_DFF_P_  (.D(\hash/e[3] ),
    .Q(\hash/e_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[4]$_DFF_P_  (.D(\hash/e[4] ),
    .Q(\hash/e_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[5]$_DFF_P_  (.D(\hash/e[5] ),
    .Q(\hash/e_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[6]$_DFF_P_  (.D(\hash/e[6] ),
    .Q(\hash/e_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[7]$_DFF_P_  (.D(\hash/e[7] ),
    .Q(\hash/e_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[8]$_DFF_P_  (.D(\hash/e[8] ),
    .Q(\hash/e_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/e_cap[9]$_DFF_P_  (.D(\hash/e[9] ),
    .Q(\hash/e_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[0]$_DFF_P_  (.D(\hash/f[0] ),
    .Q(\hash/f_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[10]$_DFF_P_  (.D(\hash/f[10] ),
    .Q(\hash/f_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[11]$_DFF_P_  (.D(\hash/f[11] ),
    .Q(\hash/f_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[12]$_DFF_P_  (.D(\hash/f[12] ),
    .Q(\hash/f_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[13]$_DFF_P_  (.D(\hash/f[13] ),
    .Q(\hash/f_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[14]$_DFF_P_  (.D(\hash/f[14] ),
    .Q(\hash/f_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[15]$_DFF_P_  (.D(\hash/f[15] ),
    .Q(\hash/f_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[16]$_DFF_P_  (.D(\hash/f[16] ),
    .Q(\hash/f_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[17]$_DFF_P_  (.D(\hash/f[17] ),
    .Q(\hash/f_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[18]$_DFF_P_  (.D(\hash/f[18] ),
    .Q(\hash/f_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[19]$_DFF_P_  (.D(\hash/f[19] ),
    .Q(\hash/f_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[1]$_DFF_P_  (.D(\hash/f[1] ),
    .Q(\hash/f_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[20]$_DFF_P_  (.D(\hash/f[20] ),
    .Q(\hash/f_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[21]$_DFF_P_  (.D(\hash/f[21] ),
    .Q(\hash/f_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[22]$_DFF_P_  (.D(\hash/f[22] ),
    .Q(\hash/f_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[23]$_DFF_P_  (.D(\hash/f[23] ),
    .Q(\hash/f_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[24]$_DFF_P_  (.D(\hash/f[24] ),
    .Q(\hash/f_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[25]$_DFF_P_  (.D(\hash/f[25] ),
    .Q(\hash/f_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[26]$_DFF_P_  (.D(\hash/f[26] ),
    .Q(\hash/f_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[27]$_DFF_P_  (.D(\hash/f[27] ),
    .Q(\hash/f_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[28]$_DFF_P_  (.D(\hash/f[28] ),
    .Q(\hash/f_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[29]$_DFF_P_  (.D(\hash/f[29] ),
    .Q(\hash/f_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[2]$_DFF_P_  (.D(\hash/f[2] ),
    .Q(\hash/f_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[30]$_DFF_P_  (.D(\hash/f[30] ),
    .Q(\hash/f_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[31]$_DFF_P_  (.D(\hash/f[31] ),
    .Q(\hash/f_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[3]$_DFF_P_  (.D(\hash/f[3] ),
    .Q(\hash/f_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[4]$_DFF_P_  (.D(\hash/f[4] ),
    .Q(\hash/f_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[5]$_DFF_P_  (.D(\hash/f[5] ),
    .Q(\hash/f_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[6]$_DFF_P_  (.D(\hash/f[6] ),
    .Q(\hash/f_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[7]$_DFF_P_  (.D(\hash/f[7] ),
    .Q(\hash/f_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[8]$_DFF_P_  (.D(\hash/f[8] ),
    .Q(\hash/f_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/f_cap[9]$_DFF_P_  (.D(\hash/f[9] ),
    .Q(\hash/f_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[0]$_DFFE_PP_  (.D(\hash/_1445_ ),
    .DE(select),
    .Q(hashvalue[224]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[10]$_DFFE_PP_  (.D(\hash/_0000_ ),
    .DE(select),
    .Q(hashvalue[234]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[11]$_DFFE_PP_  (.D(\hash/_0001_ ),
    .DE(select),
    .Q(hashvalue[235]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[12]$_DFFE_PP_  (.D(\hash/_0002_ ),
    .DE(select),
    .Q(hashvalue[236]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[13]$_DFFE_PP_  (.D(\hash/_0003_ ),
    .DE(select),
    .Q(hashvalue[237]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[14]$_DFFE_PP_  (.D(\hash/_0004_ ),
    .DE(select),
    .Q(hashvalue[238]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[15]$_DFFE_PP_  (.D(\hash/_0005_ ),
    .DE(select),
    .Q(hashvalue[239]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[16]$_DFFE_PP_  (.D(\hash/_0006_ ),
    .DE(select),
    .Q(hashvalue[240]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[17]$_DFFE_PP_  (.D(\hash/_0007_ ),
    .DE(select),
    .Q(hashvalue[241]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[18]$_DFFE_PP_  (.D(\hash/_0008_ ),
    .DE(select),
    .Q(hashvalue[242]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[19]$_DFFE_PP_  (.D(\hash/_0009_ ),
    .DE(select),
    .Q(hashvalue[243]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[1]$_DFFE_PP_  (.D(\hash/_1446_ ),
    .DE(select),
    .Q(hashvalue[225]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[20]$_DFFE_PP_  (.D(\hash/_0010_ ),
    .DE(select),
    .Q(hashvalue[244]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[21]$_DFFE_PP_  (.D(\hash/_0011_ ),
    .DE(select),
    .Q(hashvalue[245]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[22]$_DFFE_PP_  (.D(\hash/_0012_ ),
    .DE(select),
    .Q(hashvalue[246]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[23]$_DFFE_PP_  (.D(\hash/_0013_ ),
    .DE(select),
    .Q(hashvalue[247]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[24]$_DFFE_PP_  (.D(\hash/_0014_ ),
    .DE(select),
    .Q(hashvalue[248]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[25]$_DFFE_PP_  (.D(\hash/_0015_ ),
    .DE(select),
    .Q(hashvalue[249]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[26]$_DFFE_PP_  (.D(\hash/_0016_ ),
    .DE(select),
    .Q(hashvalue[250]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[27]$_DFFE_PP_  (.D(\hash/_0017_ ),
    .DE(select),
    .Q(hashvalue[251]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[28]$_DFFE_PP_  (.D(\hash/_0018_ ),
    .DE(select),
    .Q(hashvalue[252]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[29]$_DFFE_PP_  (.D(\hash/_0019_ ),
    .DE(select),
    .Q(hashvalue[253]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[2]$_DFFE_PP_  (.D(\hash/_0020_ ),
    .DE(select),
    .Q(hashvalue[226]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[30]$_DFFE_PP_  (.D(\hash/_0021_ ),
    .DE(select),
    .Q(hashvalue[254]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[31]$_DFFE_PP_  (.D(\hash/_0022_ ),
    .DE(select),
    .Q(hashvalue[255]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[3]$_DFFE_PP_  (.D(\hash/_0023_ ),
    .DE(select),
    .Q(hashvalue[227]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[4]$_DFFE_PP_  (.D(\hash/_0024_ ),
    .DE(select),
    .Q(hashvalue[228]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[5]$_DFFE_PP_  (.D(\hash/_0025_ ),
    .DE(select),
    .Q(hashvalue[229]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[6]$_DFFE_PP_  (.D(\hash/_0026_ ),
    .DE(select),
    .Q(hashvalue[230]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[7]$_DFFE_PP_  (.D(\hash/_0027_ ),
    .DE(select),
    .Q(hashvalue[231]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[8]$_DFFE_PP_  (.D(\hash/_0028_ ),
    .DE(select),
    .Q(hashvalue[232]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h0_out[9]$_DFFE_PP_  (.D(\hash/_0029_ ),
    .DE(select),
    .Q(hashvalue[233]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[0]$_DFFE_PP_  (.D(\hash/_1447_ ),
    .DE(select),
    .Q(hashvalue[192]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[10]$_DFFE_PP_  (.D(\hash/_0030_ ),
    .DE(select),
    .Q(hashvalue[202]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[11]$_DFFE_PP_  (.D(\hash/_0031_ ),
    .DE(select),
    .Q(hashvalue[203]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[12]$_DFFE_PP_  (.D(\hash/_0032_ ),
    .DE(select),
    .Q(hashvalue[204]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[13]$_DFFE_PP_  (.D(\hash/_0033_ ),
    .DE(select),
    .Q(hashvalue[205]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[14]$_DFFE_PP_  (.D(\hash/_0034_ ),
    .DE(select),
    .Q(hashvalue[206]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[15]$_DFFE_PP_  (.D(\hash/_0035_ ),
    .DE(select),
    .Q(hashvalue[207]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[16]$_DFFE_PP_  (.D(\hash/_0036_ ),
    .DE(select),
    .Q(hashvalue[208]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[17]$_DFFE_PP_  (.D(\hash/_0037_ ),
    .DE(select),
    .Q(hashvalue[209]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[18]$_DFFE_PP_  (.D(\hash/_0038_ ),
    .DE(select),
    .Q(hashvalue[210]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[19]$_DFFE_PP_  (.D(\hash/_0039_ ),
    .DE(select),
    .Q(hashvalue[211]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[1]$_DFFE_PP_  (.D(\hash/_1448_ ),
    .DE(select),
    .Q(hashvalue[193]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[20]$_DFFE_PP_  (.D(\hash/_0040_ ),
    .DE(select),
    .Q(hashvalue[212]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[21]$_DFFE_PP_  (.D(\hash/_0041_ ),
    .DE(select),
    .Q(hashvalue[213]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[22]$_DFFE_PP_  (.D(\hash/_0042_ ),
    .DE(select),
    .Q(hashvalue[214]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[23]$_DFFE_PP_  (.D(\hash/_0043_ ),
    .DE(select),
    .Q(hashvalue[215]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[24]$_DFFE_PP_  (.D(\hash/_0044_ ),
    .DE(select),
    .Q(hashvalue[216]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[25]$_DFFE_PP_  (.D(\hash/_0045_ ),
    .DE(select),
    .Q(hashvalue[217]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[26]$_DFFE_PP_  (.D(\hash/_0046_ ),
    .DE(select),
    .Q(hashvalue[218]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[27]$_DFFE_PP_  (.D(\hash/_0047_ ),
    .DE(select),
    .Q(hashvalue[219]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[28]$_DFFE_PP_  (.D(\hash/_0048_ ),
    .DE(select),
    .Q(hashvalue[220]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[29]$_DFFE_PP_  (.D(\hash/_0049_ ),
    .DE(select),
    .Q(hashvalue[221]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[2]$_DFFE_PP_  (.D(\hash/_0050_ ),
    .DE(select),
    .Q(hashvalue[194]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[30]$_DFFE_PP_  (.D(\hash/_0051_ ),
    .DE(select),
    .Q(hashvalue[222]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[31]$_DFFE_PP_  (.D(\hash/_0052_ ),
    .DE(select),
    .Q(hashvalue[223]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[3]$_DFFE_PP_  (.D(\hash/_0053_ ),
    .DE(select),
    .Q(hashvalue[195]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[4]$_DFFE_PP_  (.D(\hash/_0054_ ),
    .DE(select),
    .Q(hashvalue[196]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[5]$_DFFE_PP_  (.D(\hash/_0055_ ),
    .DE(select),
    .Q(hashvalue[197]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[6]$_DFFE_PP_  (.D(\hash/_0056_ ),
    .DE(select),
    .Q(hashvalue[198]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[7]$_DFFE_PP_  (.D(\hash/_0057_ ),
    .DE(select),
    .Q(hashvalue[199]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[8]$_DFFE_PP_  (.D(\hash/_0058_ ),
    .DE(select),
    .Q(hashvalue[200]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h1_out[9]$_DFFE_PP_  (.D(\hash/_0059_ ),
    .DE(select),
    .Q(hashvalue[201]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[0]$_DFFE_PP_  (.D(\hash/_1449_ ),
    .DE(select),
    .Q(hashvalue[160]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[10]$_DFFE_PP_  (.D(\hash/_0060_ ),
    .DE(select),
    .Q(hashvalue[170]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[11]$_DFFE_PP_  (.D(\hash/_0061_ ),
    .DE(select),
    .Q(hashvalue[171]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[12]$_DFFE_PP_  (.D(\hash/_0062_ ),
    .DE(select),
    .Q(hashvalue[172]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[13]$_DFFE_PP_  (.D(\hash/_0063_ ),
    .DE(select),
    .Q(hashvalue[173]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[14]$_DFFE_PP_  (.D(\hash/_0064_ ),
    .DE(select),
    .Q(hashvalue[174]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[15]$_DFFE_PP_  (.D(\hash/_0065_ ),
    .DE(select),
    .Q(hashvalue[175]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[16]$_DFFE_PP_  (.D(\hash/_0066_ ),
    .DE(select),
    .Q(hashvalue[176]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[17]$_DFFE_PP_  (.D(\hash/_0067_ ),
    .DE(select),
    .Q(hashvalue[177]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[18]$_DFFE_PP_  (.D(\hash/_0068_ ),
    .DE(select),
    .Q(hashvalue[178]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[19]$_DFFE_PP_  (.D(\hash/_0069_ ),
    .DE(select),
    .Q(hashvalue[179]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[1]$_DFFE_PP_  (.D(\hash/_1450_ ),
    .DE(select),
    .Q(hashvalue[161]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[20]$_DFFE_PP_  (.D(\hash/_0070_ ),
    .DE(select),
    .Q(hashvalue[180]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[21]$_DFFE_PP_  (.D(\hash/_0071_ ),
    .DE(select),
    .Q(hashvalue[181]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[22]$_DFFE_PP_  (.D(\hash/_0072_ ),
    .DE(select),
    .Q(hashvalue[182]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[23]$_DFFE_PP_  (.D(\hash/_0073_ ),
    .DE(select),
    .Q(hashvalue[183]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[24]$_DFFE_PP_  (.D(\hash/_0074_ ),
    .DE(select),
    .Q(hashvalue[184]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[25]$_DFFE_PP_  (.D(\hash/_0075_ ),
    .DE(select),
    .Q(hashvalue[185]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[26]$_DFFE_PP_  (.D(\hash/_0076_ ),
    .DE(select),
    .Q(hashvalue[186]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[27]$_DFFE_PP_  (.D(\hash/_0077_ ),
    .DE(select),
    .Q(hashvalue[187]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[28]$_DFFE_PP_  (.D(\hash/_0078_ ),
    .DE(select),
    .Q(hashvalue[188]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[29]$_DFFE_PP_  (.D(\hash/_0079_ ),
    .DE(select),
    .Q(hashvalue[189]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[2]$_DFFE_PP_  (.D(\hash/_0080_ ),
    .DE(select),
    .Q(hashvalue[162]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[30]$_DFFE_PP_  (.D(\hash/_0081_ ),
    .DE(select),
    .Q(hashvalue[190]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[31]$_DFFE_PP_  (.D(\hash/_0082_ ),
    .DE(select),
    .Q(hashvalue[191]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[3]$_DFFE_PP_  (.D(\hash/_0083_ ),
    .DE(select),
    .Q(hashvalue[163]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[4]$_DFFE_PP_  (.D(\hash/_0084_ ),
    .DE(select),
    .Q(hashvalue[164]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[5]$_DFFE_PP_  (.D(\hash/_0085_ ),
    .DE(select),
    .Q(hashvalue[165]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[6]$_DFFE_PP_  (.D(\hash/_0086_ ),
    .DE(select),
    .Q(hashvalue[166]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[7]$_DFFE_PP_  (.D(\hash/_0087_ ),
    .DE(select),
    .Q(hashvalue[167]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[8]$_DFFE_PP_  (.D(\hash/_0088_ ),
    .DE(select),
    .Q(hashvalue[168]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h2_out[9]$_DFFE_PP_  (.D(\hash/_0089_ ),
    .DE(select),
    .Q(hashvalue[169]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[0]$_DFFE_PP_  (.D(\hash/_1451_ ),
    .DE(select),
    .Q(hashvalue[128]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[10]$_DFFE_PP_  (.D(\hash/_0090_ ),
    .DE(select),
    .Q(hashvalue[138]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[11]$_DFFE_PP_  (.D(\hash/_0091_ ),
    .DE(select),
    .Q(hashvalue[139]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[12]$_DFFE_PP_  (.D(\hash/_0092_ ),
    .DE(select),
    .Q(hashvalue[140]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[13]$_DFFE_PP_  (.D(\hash/_0093_ ),
    .DE(select),
    .Q(hashvalue[141]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[14]$_DFFE_PP_  (.D(\hash/_0094_ ),
    .DE(select),
    .Q(hashvalue[142]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[15]$_DFFE_PP_  (.D(\hash/_0095_ ),
    .DE(select),
    .Q(hashvalue[143]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[16]$_DFFE_PP_  (.D(\hash/_0096_ ),
    .DE(select),
    .Q(hashvalue[144]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[17]$_DFFE_PP_  (.D(\hash/_0097_ ),
    .DE(select),
    .Q(hashvalue[145]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[18]$_DFFE_PP_  (.D(\hash/_0098_ ),
    .DE(select),
    .Q(hashvalue[146]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[19]$_DFFE_PP_  (.D(\hash/_0099_ ),
    .DE(select),
    .Q(hashvalue[147]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[1]$_DFFE_PP_  (.D(\hash/_1452_ ),
    .DE(select),
    .Q(hashvalue[129]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[20]$_DFFE_PP_  (.D(\hash/_0100_ ),
    .DE(select),
    .Q(hashvalue[148]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[21]$_DFFE_PP_  (.D(\hash/_0101_ ),
    .DE(select),
    .Q(hashvalue[149]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[22]$_DFFE_PP_  (.D(\hash/_0102_ ),
    .DE(select),
    .Q(hashvalue[150]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[23]$_DFFE_PP_  (.D(\hash/_0103_ ),
    .DE(select),
    .Q(hashvalue[151]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[24]$_DFFE_PP_  (.D(\hash/_0104_ ),
    .DE(select),
    .Q(hashvalue[152]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[25]$_DFFE_PP_  (.D(\hash/_0105_ ),
    .DE(select),
    .Q(hashvalue[153]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[26]$_DFFE_PP_  (.D(\hash/_0106_ ),
    .DE(select),
    .Q(hashvalue[154]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[27]$_DFFE_PP_  (.D(\hash/_0107_ ),
    .DE(select),
    .Q(hashvalue[155]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[28]$_DFFE_PP_  (.D(\hash/_0108_ ),
    .DE(select),
    .Q(hashvalue[156]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[29]$_DFFE_PP_  (.D(\hash/_0109_ ),
    .DE(select),
    .Q(hashvalue[157]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[2]$_DFFE_PP_  (.D(\hash/_0110_ ),
    .DE(select),
    .Q(hashvalue[130]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[30]$_DFFE_PP_  (.D(\hash/_0111_ ),
    .DE(select),
    .Q(hashvalue[158]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[31]$_DFFE_PP_  (.D(\hash/_0112_ ),
    .DE(select),
    .Q(hashvalue[159]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[3]$_DFFE_PP_  (.D(\hash/_0113_ ),
    .DE(select),
    .Q(hashvalue[131]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[4]$_DFFE_PP_  (.D(\hash/_0114_ ),
    .DE(select),
    .Q(hashvalue[132]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[5]$_DFFE_PP_  (.D(\hash/_0115_ ),
    .DE(select),
    .Q(hashvalue[133]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[6]$_DFFE_PP_  (.D(\hash/_0116_ ),
    .DE(select),
    .Q(hashvalue[134]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[7]$_DFFE_PP_  (.D(\hash/_0117_ ),
    .DE(select),
    .Q(hashvalue[135]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[8]$_DFFE_PP_  (.D(\hash/_0118_ ),
    .DE(select),
    .Q(hashvalue[136]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h3_out[9]$_DFFE_PP_  (.D(\hash/_0119_ ),
    .DE(select),
    .Q(hashvalue[137]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[0]$_DFFE_PP_  (.D(\hash/_1453_ ),
    .DE(select),
    .Q(hashvalue[96]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[10]$_DFFE_PP_  (.D(\hash/_0120_ ),
    .DE(select),
    .Q(hashvalue[106]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[11]$_DFFE_PP_  (.D(\hash/_0121_ ),
    .DE(select),
    .Q(hashvalue[107]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[12]$_DFFE_PP_  (.D(\hash/_0122_ ),
    .DE(select),
    .Q(hashvalue[108]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[13]$_DFFE_PP_  (.D(\hash/_0123_ ),
    .DE(select),
    .Q(hashvalue[109]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[14]$_DFFE_PP_  (.D(\hash/_0124_ ),
    .DE(select),
    .Q(hashvalue[110]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[15]$_DFFE_PP_  (.D(\hash/_0125_ ),
    .DE(select),
    .Q(hashvalue[111]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[16]$_DFFE_PP_  (.D(\hash/_0126_ ),
    .DE(select),
    .Q(hashvalue[112]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[17]$_DFFE_PP_  (.D(\hash/_0127_ ),
    .DE(select),
    .Q(hashvalue[113]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[18]$_DFFE_PP_  (.D(\hash/_0128_ ),
    .DE(select),
    .Q(hashvalue[114]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[19]$_DFFE_PP_  (.D(\hash/_0129_ ),
    .DE(select),
    .Q(hashvalue[115]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[1]$_DFFE_PP_  (.D(\hash/_1454_ ),
    .DE(select),
    .Q(hashvalue[97]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[20]$_DFFE_PP_  (.D(\hash/_0130_ ),
    .DE(select),
    .Q(hashvalue[116]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[21]$_DFFE_PP_  (.D(\hash/_0131_ ),
    .DE(select),
    .Q(hashvalue[117]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[22]$_DFFE_PP_  (.D(\hash/_0132_ ),
    .DE(select),
    .Q(hashvalue[118]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[23]$_DFFE_PP_  (.D(\hash/_0133_ ),
    .DE(select),
    .Q(hashvalue[119]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[24]$_DFFE_PP_  (.D(\hash/_0134_ ),
    .DE(select),
    .Q(hashvalue[120]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[25]$_DFFE_PP_  (.D(\hash/_0135_ ),
    .DE(select),
    .Q(hashvalue[121]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[26]$_DFFE_PP_  (.D(\hash/_0136_ ),
    .DE(select),
    .Q(hashvalue[122]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[27]$_DFFE_PP_  (.D(\hash/_0137_ ),
    .DE(select),
    .Q(hashvalue[123]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[28]$_DFFE_PP_  (.D(\hash/_0138_ ),
    .DE(select),
    .Q(hashvalue[124]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[29]$_DFFE_PP_  (.D(\hash/_0139_ ),
    .DE(select),
    .Q(hashvalue[125]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[2]$_DFFE_PP_  (.D(\hash/_0140_ ),
    .DE(select),
    .Q(hashvalue[98]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[30]$_DFFE_PP_  (.D(\hash/_0141_ ),
    .DE(select),
    .Q(hashvalue[126]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[31]$_DFFE_PP_  (.D(\hash/_0142_ ),
    .DE(select),
    .Q(hashvalue[127]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[3]$_DFFE_PP_  (.D(\hash/_0143_ ),
    .DE(select),
    .Q(hashvalue[99]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[4]$_DFFE_PP_  (.D(\hash/_0144_ ),
    .DE(select),
    .Q(hashvalue[100]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[5]$_DFFE_PP_  (.D(\hash/_0145_ ),
    .DE(select),
    .Q(hashvalue[101]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[6]$_DFFE_PP_  (.D(\hash/_0146_ ),
    .DE(select),
    .Q(hashvalue[102]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[7]$_DFFE_PP_  (.D(\hash/_0147_ ),
    .DE(select),
    .Q(hashvalue[103]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[8]$_DFFE_PP_  (.D(\hash/_0148_ ),
    .DE(select),
    .Q(hashvalue[104]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h4_out[9]$_DFFE_PP_  (.D(\hash/_0149_ ),
    .DE(select),
    .Q(hashvalue[105]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[0]$_DFFE_PP_  (.D(\hash/_1455_ ),
    .DE(select),
    .Q(hashvalue[64]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[10]$_DFFE_PP_  (.D(\hash/_0150_ ),
    .DE(select),
    .Q(hashvalue[74]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[11]$_DFFE_PP_  (.D(\hash/_0151_ ),
    .DE(select),
    .Q(hashvalue[75]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[12]$_DFFE_PP_  (.D(\hash/_0152_ ),
    .DE(select),
    .Q(hashvalue[76]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[13]$_DFFE_PP_  (.D(\hash/_0153_ ),
    .DE(select),
    .Q(hashvalue[77]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[14]$_DFFE_PP_  (.D(\hash/_0154_ ),
    .DE(select),
    .Q(hashvalue[78]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[15]$_DFFE_PP_  (.D(\hash/_0155_ ),
    .DE(select),
    .Q(hashvalue[79]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[16]$_DFFE_PP_  (.D(\hash/_0156_ ),
    .DE(select),
    .Q(hashvalue[80]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[17]$_DFFE_PP_  (.D(\hash/_0157_ ),
    .DE(select),
    .Q(hashvalue[81]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[18]$_DFFE_PP_  (.D(\hash/_0158_ ),
    .DE(select),
    .Q(hashvalue[82]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[19]$_DFFE_PP_  (.D(\hash/_0159_ ),
    .DE(select),
    .Q(hashvalue[83]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[1]$_DFFE_PP_  (.D(\hash/_1456_ ),
    .DE(select),
    .Q(hashvalue[65]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[20]$_DFFE_PP_  (.D(\hash/_0160_ ),
    .DE(select),
    .Q(hashvalue[84]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[21]$_DFFE_PP_  (.D(\hash/_0161_ ),
    .DE(select),
    .Q(hashvalue[85]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[22]$_DFFE_PP_  (.D(\hash/_0162_ ),
    .DE(select),
    .Q(hashvalue[86]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[23]$_DFFE_PP_  (.D(\hash/_0163_ ),
    .DE(select),
    .Q(hashvalue[87]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[24]$_DFFE_PP_  (.D(\hash/_0164_ ),
    .DE(select),
    .Q(hashvalue[88]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[25]$_DFFE_PP_  (.D(\hash/_0165_ ),
    .DE(select),
    .Q(hashvalue[89]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[26]$_DFFE_PP_  (.D(\hash/_0166_ ),
    .DE(select),
    .Q(hashvalue[90]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[27]$_DFFE_PP_  (.D(\hash/_0167_ ),
    .DE(select),
    .Q(hashvalue[91]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[28]$_DFFE_PP_  (.D(\hash/_0168_ ),
    .DE(select),
    .Q(hashvalue[92]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[29]$_DFFE_PP_  (.D(\hash/_0169_ ),
    .DE(select),
    .Q(hashvalue[93]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[2]$_DFFE_PP_  (.D(\hash/_0170_ ),
    .DE(select),
    .Q(hashvalue[66]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[30]$_DFFE_PP_  (.D(\hash/_0171_ ),
    .DE(select),
    .Q(hashvalue[94]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[31]$_DFFE_PP_  (.D(\hash/_0172_ ),
    .DE(select),
    .Q(hashvalue[95]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[3]$_DFFE_PP_  (.D(\hash/_0173_ ),
    .DE(select),
    .Q(hashvalue[67]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[4]$_DFFE_PP_  (.D(\hash/_0174_ ),
    .DE(select),
    .Q(hashvalue[68]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[5]$_DFFE_PP_  (.D(\hash/_0175_ ),
    .DE(select),
    .Q(hashvalue[69]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[6]$_DFFE_PP_  (.D(\hash/_0176_ ),
    .DE(select),
    .Q(hashvalue[70]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[7]$_DFFE_PP_  (.D(\hash/_0177_ ),
    .DE(select),
    .Q(hashvalue[71]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[8]$_DFFE_PP_  (.D(\hash/_0178_ ),
    .DE(select),
    .Q(hashvalue[72]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h5_out[9]$_DFFE_PP_  (.D(\hash/_0179_ ),
    .DE(select),
    .Q(hashvalue[73]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[0]$_DFFE_PP_  (.D(\hash/_1457_ ),
    .DE(select),
    .Q(hashvalue[32]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[10]$_DFFE_PP_  (.D(\hash/_0180_ ),
    .DE(select),
    .Q(hashvalue[42]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[11]$_DFFE_PP_  (.D(\hash/_0181_ ),
    .DE(select),
    .Q(hashvalue[43]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[12]$_DFFE_PP_  (.D(\hash/_0182_ ),
    .DE(select),
    .Q(hashvalue[44]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[13]$_DFFE_PP_  (.D(\hash/_0183_ ),
    .DE(select),
    .Q(hashvalue[45]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[14]$_DFFE_PP_  (.D(\hash/_0184_ ),
    .DE(select),
    .Q(hashvalue[46]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[15]$_DFFE_PP_  (.D(\hash/_0185_ ),
    .DE(select),
    .Q(hashvalue[47]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[16]$_DFFE_PP_  (.D(\hash/_0186_ ),
    .DE(select),
    .Q(hashvalue[48]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[17]$_DFFE_PP_  (.D(\hash/_0187_ ),
    .DE(select),
    .Q(hashvalue[49]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[18]$_DFFE_PP_  (.D(\hash/_0188_ ),
    .DE(select),
    .Q(hashvalue[50]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[19]$_DFFE_PP_  (.D(\hash/_0189_ ),
    .DE(select),
    .Q(hashvalue[51]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[1]$_DFFE_PP_  (.D(\hash/_1458_ ),
    .DE(select),
    .Q(hashvalue[33]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[20]$_DFFE_PP_  (.D(\hash/_0190_ ),
    .DE(select),
    .Q(hashvalue[52]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[21]$_DFFE_PP_  (.D(\hash/_0191_ ),
    .DE(select),
    .Q(hashvalue[53]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[22]$_DFFE_PP_  (.D(\hash/_0192_ ),
    .DE(select),
    .Q(hashvalue[54]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[23]$_DFFE_PP_  (.D(\hash/_0193_ ),
    .DE(select),
    .Q(hashvalue[55]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[24]$_DFFE_PP_  (.D(\hash/_0194_ ),
    .DE(select),
    .Q(hashvalue[56]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[25]$_DFFE_PP_  (.D(\hash/_0195_ ),
    .DE(select),
    .Q(hashvalue[57]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[26]$_DFFE_PP_  (.D(\hash/_0196_ ),
    .DE(select),
    .Q(hashvalue[58]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[27]$_DFFE_PP_  (.D(\hash/_0197_ ),
    .DE(select),
    .Q(hashvalue[59]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[28]$_DFFE_PP_  (.D(\hash/_0198_ ),
    .DE(select),
    .Q(hashvalue[60]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[29]$_DFFE_PP_  (.D(\hash/_0199_ ),
    .DE(select),
    .Q(hashvalue[61]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[2]$_DFFE_PP_  (.D(\hash/_0200_ ),
    .DE(select),
    .Q(hashvalue[34]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[30]$_DFFE_PP_  (.D(\hash/_0201_ ),
    .DE(select),
    .Q(hashvalue[62]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[31]$_DFFE_PP_  (.D(\hash/_0202_ ),
    .DE(select),
    .Q(hashvalue[63]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[3]$_DFFE_PP_  (.D(\hash/_0203_ ),
    .DE(select),
    .Q(hashvalue[35]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[4]$_DFFE_PP_  (.D(\hash/_0204_ ),
    .DE(select),
    .Q(hashvalue[36]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[5]$_DFFE_PP_  (.D(\hash/_0205_ ),
    .DE(select),
    .Q(hashvalue[37]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[6]$_DFFE_PP_  (.D(\hash/_0206_ ),
    .DE(select),
    .Q(hashvalue[38]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[7]$_DFFE_PP_  (.D(\hash/_0207_ ),
    .DE(select),
    .Q(hashvalue[39]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[8]$_DFFE_PP_  (.D(\hash/_0208_ ),
    .DE(select),
    .Q(hashvalue[40]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h6_out[9]$_DFFE_PP_  (.D(\hash/_0209_ ),
    .DE(select),
    .Q(hashvalue[41]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[0]$_DFFE_PP_  (.D(\hash/_1459_ ),
    .DE(select),
    .Q(hashvalue[0]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[10]$_DFFE_PP_  (.D(\hash/_0210_ ),
    .DE(select),
    .Q(hashvalue[10]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[11]$_DFFE_PP_  (.D(\hash/_0211_ ),
    .DE(select),
    .Q(hashvalue[11]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[12]$_DFFE_PP_  (.D(\hash/_0212_ ),
    .DE(select),
    .Q(hashvalue[12]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[13]$_DFFE_PP_  (.D(\hash/_0213_ ),
    .DE(select),
    .Q(hashvalue[13]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[14]$_DFFE_PP_  (.D(\hash/_0214_ ),
    .DE(select),
    .Q(hashvalue[14]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[15]$_DFFE_PP_  (.D(\hash/_0215_ ),
    .DE(select),
    .Q(hashvalue[15]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[16]$_DFFE_PP_  (.D(\hash/_0216_ ),
    .DE(select),
    .Q(hashvalue[16]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[17]$_DFFE_PP_  (.D(\hash/_0217_ ),
    .DE(select),
    .Q(hashvalue[17]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[18]$_DFFE_PP_  (.D(\hash/_0218_ ),
    .DE(select),
    .Q(hashvalue[18]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[19]$_DFFE_PP_  (.D(\hash/_0219_ ),
    .DE(select),
    .Q(hashvalue[19]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[1]$_DFFE_PP_  (.D(\hash/_1460_ ),
    .DE(select),
    .Q(hashvalue[1]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[20]$_DFFE_PP_  (.D(\hash/_0220_ ),
    .DE(select),
    .Q(hashvalue[20]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[21]$_DFFE_PP_  (.D(\hash/_0221_ ),
    .DE(select),
    .Q(hashvalue[21]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[22]$_DFFE_PP_  (.D(\hash/_0222_ ),
    .DE(select),
    .Q(hashvalue[22]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[23]$_DFFE_PP_  (.D(\hash/_0223_ ),
    .DE(select),
    .Q(hashvalue[23]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[24]$_DFFE_PP_  (.D(\hash/_0224_ ),
    .DE(select),
    .Q(hashvalue[24]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[25]$_DFFE_PP_  (.D(\hash/_0225_ ),
    .DE(select),
    .Q(hashvalue[25]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[26]$_DFFE_PP_  (.D(\hash/_0226_ ),
    .DE(select),
    .Q(hashvalue[26]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[27]$_DFFE_PP_  (.D(\hash/_0227_ ),
    .DE(select),
    .Q(hashvalue[27]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[28]$_DFFE_PP_  (.D(\hash/_0228_ ),
    .DE(select),
    .Q(hashvalue[28]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[29]$_DFFE_PP_  (.D(\hash/_0229_ ),
    .DE(select),
    .Q(hashvalue[29]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[2]$_DFFE_PP_  (.D(\hash/_0230_ ),
    .DE(select),
    .Q(hashvalue[2]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[30]$_DFFE_PP_  (.D(\hash/_0231_ ),
    .DE(select),
    .Q(hashvalue[30]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[31]$_DFFE_PP_  (.D(\hash/_0232_ ),
    .DE(select),
    .Q(hashvalue[31]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[3]$_DFFE_PP_  (.D(\hash/_0233_ ),
    .DE(select),
    .Q(hashvalue[3]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[4]$_DFFE_PP_  (.D(\hash/_0234_ ),
    .DE(select),
    .Q(hashvalue[4]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[5]$_DFFE_PP_  (.D(\hash/_0235_ ),
    .DE(select),
    .Q(hashvalue[5]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[6]$_DFFE_PP_  (.D(\hash/_0236_ ),
    .DE(select),
    .Q(hashvalue[6]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[7]$_DFFE_PP_  (.D(\hash/_0237_ ),
    .DE(select),
    .Q(hashvalue[7]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[8]$_DFFE_PP_  (.D(\hash/_0238_ ),
    .DE(select),
    .Q(hashvalue[8]),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \hash/h7_out[9]$_DFFE_PP_  (.D(\hash/_0239_ ),
    .DE(select),
    .Q(hashvalue[9]),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[0]$_DFF_P_  (.D(\hash/p1[0] ),
    .Q(\hash/p1_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[10]$_DFF_P_  (.D(\hash/p1[10] ),
    .Q(\hash/p1_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[11]$_DFF_P_  (.D(\hash/p1[11] ),
    .Q(\hash/p1_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[12]$_DFF_P_  (.D(\hash/p1[12] ),
    .Q(\hash/p1_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[13]$_DFF_P_  (.D(\hash/p1[13] ),
    .Q(\hash/p1_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[14]$_DFF_P_  (.D(\hash/p1[14] ),
    .Q(\hash/p1_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[15]$_DFF_P_  (.D(\hash/p1[15] ),
    .Q(\hash/p1_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[16]$_DFF_P_  (.D(\hash/p1[16] ),
    .Q(\hash/p1_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[17]$_DFF_P_  (.D(\hash/p1[17] ),
    .Q(\hash/p1_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[18]$_DFF_P_  (.D(\hash/p1[18] ),
    .Q(\hash/p1_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[19]$_DFF_P_  (.D(\hash/p1[19] ),
    .Q(\hash/p1_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[1]$_DFF_P_  (.D(\hash/p1[1] ),
    .Q(\hash/p1_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[20]$_DFF_P_  (.D(\hash/p1[20] ),
    .Q(\hash/p1_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[21]$_DFF_P_  (.D(\hash/p1[21] ),
    .Q(\hash/p1_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[22]$_DFF_P_  (.D(\hash/p1[22] ),
    .Q(\hash/p1_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[23]$_DFF_P_  (.D(\hash/p1[23] ),
    .Q(\hash/p1_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[24]$_DFF_P_  (.D(\hash/p1[24] ),
    .Q(\hash/p1_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[25]$_DFF_P_  (.D(\hash/p1[25] ),
    .Q(\hash/p1_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[26]$_DFF_P_  (.D(\hash/p1[26] ),
    .Q(\hash/p1_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[27]$_DFF_P_  (.D(\hash/p1[27] ),
    .Q(\hash/p1_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[28]$_DFF_P_  (.D(\hash/p1[28] ),
    .Q(\hash/p1_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[29]$_DFF_P_  (.D(\hash/p1[29] ),
    .Q(\hash/p1_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[2]$_DFF_P_  (.D(\hash/p1[2] ),
    .Q(\hash/p1_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[30]$_DFF_P_  (.D(\hash/p1[30] ),
    .Q(\hash/p1_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[31]$_DFF_P_  (.D(\hash/p1[31] ),
    .Q(\hash/p1_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[3]$_DFF_P_  (.D(\hash/p1[3] ),
    .Q(\hash/p1_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[4]$_DFF_P_  (.D(\hash/p1[4] ),
    .Q(\hash/p1_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[5]$_DFF_P_  (.D(\hash/p1[5] ),
    .Q(\hash/p1_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[6]$_DFF_P_  (.D(\hash/p1[6] ),
    .Q(\hash/p1_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[7]$_DFF_P_  (.D(\hash/p1[7] ),
    .Q(\hash/p1_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[8]$_DFF_P_  (.D(\hash/p1[8] ),
    .Q(\hash/p1_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p1_cap[9]$_DFF_P_  (.D(\hash/p1[9] ),
    .Q(\hash/p1_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[0]$_DFF_P_  (.D(\hash/p2[0] ),
    .Q(\hash/p2_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[10]$_DFF_P_  (.D(\hash/p2[10] ),
    .Q(\hash/p2_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[11]$_DFF_P_  (.D(\hash/p2[11] ),
    .Q(\hash/p2_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[12]$_DFF_P_  (.D(\hash/p2[12] ),
    .Q(\hash/p2_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[13]$_DFF_P_  (.D(\hash/p2[13] ),
    .Q(\hash/p2_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[14]$_DFF_P_  (.D(\hash/p2[14] ),
    .Q(\hash/p2_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[15]$_DFF_P_  (.D(\hash/p2[15] ),
    .Q(\hash/p2_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[16]$_DFF_P_  (.D(\hash/p2[16] ),
    .Q(\hash/p2_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[17]$_DFF_P_  (.D(\hash/p2[17] ),
    .Q(\hash/p2_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[18]$_DFF_P_  (.D(\hash/p2[18] ),
    .Q(\hash/p2_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[19]$_DFF_P_  (.D(\hash/p2[19] ),
    .Q(\hash/p2_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[1]$_DFF_P_  (.D(\hash/p2[1] ),
    .Q(\hash/p2_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[20]$_DFF_P_  (.D(\hash/p2[20] ),
    .Q(\hash/p2_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[21]$_DFF_P_  (.D(\hash/p2[21] ),
    .Q(\hash/p2_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[22]$_DFF_P_  (.D(\hash/p2[22] ),
    .Q(\hash/p2_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[23]$_DFF_P_  (.D(\hash/p2[23] ),
    .Q(\hash/p2_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[24]$_DFF_P_  (.D(\hash/p2[24] ),
    .Q(\hash/p2_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[25]$_DFF_P_  (.D(\hash/p2[25] ),
    .Q(\hash/p2_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[26]$_DFF_P_  (.D(\hash/p2[26] ),
    .Q(\hash/p2_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[27]$_DFF_P_  (.D(\hash/p2[27] ),
    .Q(\hash/p2_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[28]$_DFF_P_  (.D(\hash/p2[28] ),
    .Q(\hash/p2_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[29]$_DFF_P_  (.D(\hash/p2[29] ),
    .Q(\hash/p2_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[2]$_DFF_P_  (.D(\hash/p2[2] ),
    .Q(\hash/p2_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[30]$_DFF_P_  (.D(\hash/p2[30] ),
    .Q(\hash/p2_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[31]$_DFF_P_  (.D(\hash/p2[31] ),
    .Q(\hash/p2_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[3]$_DFF_P_  (.D(\hash/p2[3] ),
    .Q(\hash/p2_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[4]$_DFF_P_  (.D(\hash/p2[4] ),
    .Q(\hash/p2_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[5]$_DFF_P_  (.D(\hash/p2[5] ),
    .Q(\hash/p2_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[6]$_DFF_P_  (.D(\hash/p2[6] ),
    .Q(\hash/p2_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[7]$_DFF_P_  (.D(\hash/p2[7] ),
    .Q(\hash/p2_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[8]$_DFF_P_  (.D(\hash/p2[8] ),
    .Q(\hash/p2_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p2_cap[9]$_DFF_P_  (.D(\hash/p2[9] ),
    .Q(\hash/p2_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[0]$_DFF_P_  (.D(\hash/p3[0] ),
    .Q(\hash/p3_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[10]$_DFF_P_  (.D(\hash/p3[10] ),
    .Q(\hash/p3_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[11]$_DFF_P_  (.D(\hash/p3[11] ),
    .Q(\hash/p3_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[12]$_DFF_P_  (.D(\hash/p3[12] ),
    .Q(\hash/p3_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[13]$_DFF_P_  (.D(\hash/p3[13] ),
    .Q(\hash/p3_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[14]$_DFF_P_  (.D(\hash/p3[14] ),
    .Q(\hash/p3_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[15]$_DFF_P_  (.D(\hash/p3[15] ),
    .Q(\hash/p3_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[16]$_DFF_P_  (.D(\hash/p3[16] ),
    .Q(\hash/p3_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[17]$_DFF_P_  (.D(\hash/p3[17] ),
    .Q(\hash/p3_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[18]$_DFF_P_  (.D(\hash/p3[18] ),
    .Q(\hash/p3_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[19]$_DFF_P_  (.D(\hash/p3[19] ),
    .Q(\hash/p3_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[1]$_DFF_P_  (.D(\hash/p3[1] ),
    .Q(\hash/p3_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[20]$_DFF_P_  (.D(\hash/p3[20] ),
    .Q(\hash/p3_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[21]$_DFF_P_  (.D(\hash/p3[21] ),
    .Q(\hash/p3_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[22]$_DFF_P_  (.D(\hash/p3[22] ),
    .Q(\hash/p3_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[23]$_DFF_P_  (.D(\hash/p3[23] ),
    .Q(\hash/p3_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[24]$_DFF_P_  (.D(\hash/p3[24] ),
    .Q(\hash/p3_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[25]$_DFF_P_  (.D(\hash/p3[25] ),
    .Q(\hash/p3_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[26]$_DFF_P_  (.D(\hash/p3[26] ),
    .Q(\hash/p3_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[27]$_DFF_P_  (.D(\hash/p3[27] ),
    .Q(\hash/p3_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[28]$_DFF_P_  (.D(\hash/p3[28] ),
    .Q(\hash/p3_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[29]$_DFF_P_  (.D(\hash/p3[29] ),
    .Q(\hash/p3_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[2]$_DFF_P_  (.D(\hash/p3[2] ),
    .Q(\hash/p3_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[30]$_DFF_P_  (.D(\hash/p3[30] ),
    .Q(\hash/p3_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[31]$_DFF_P_  (.D(\hash/p3[31] ),
    .Q(\hash/p3_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[3]$_DFF_P_  (.D(\hash/p3[3] ),
    .Q(\hash/p3_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[4]$_DFF_P_  (.D(\hash/p3[4] ),
    .Q(\hash/p3_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[5]$_DFF_P_  (.D(\hash/p3[5] ),
    .Q(\hash/p3_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[6]$_DFF_P_  (.D(\hash/p3[6] ),
    .Q(\hash/p3_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[7]$_DFF_P_  (.D(\hash/p3[7] ),
    .Q(\hash/p3_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[8]$_DFF_P_  (.D(\hash/p3[8] ),
    .Q(\hash/p3_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p3_cap[9]$_DFF_P_  (.D(\hash/p3[9] ),
    .Q(\hash/p3_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[0]$_DFF_P_  (.D(\hash/p4[0] ),
    .Q(\hash/p4_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[10]$_DFF_P_  (.D(\hash/p4[10] ),
    .Q(\hash/p4_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[11]$_DFF_P_  (.D(\hash/p4[11] ),
    .Q(\hash/p4_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[12]$_DFF_P_  (.D(\hash/p4[12] ),
    .Q(\hash/p4_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[13]$_DFF_P_  (.D(\hash/p4[13] ),
    .Q(\hash/p4_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[14]$_DFF_P_  (.D(\hash/p4[14] ),
    .Q(\hash/p4_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[15]$_DFF_P_  (.D(\hash/p4[15] ),
    .Q(\hash/p4_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[16]$_DFF_P_  (.D(\hash/p4[16] ),
    .Q(\hash/p4_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[17]$_DFF_P_  (.D(\hash/p4[17] ),
    .Q(\hash/p4_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[18]$_DFF_P_  (.D(\hash/p4[18] ),
    .Q(\hash/p4_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[19]$_DFF_P_  (.D(\hash/p4[19] ),
    .Q(\hash/p4_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[1]$_DFF_P_  (.D(\hash/p4[1] ),
    .Q(\hash/p4_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[20]$_DFF_P_  (.D(\hash/p4[20] ),
    .Q(\hash/p4_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[21]$_DFF_P_  (.D(\hash/p4[21] ),
    .Q(\hash/p4_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[22]$_DFF_P_  (.D(\hash/p4[22] ),
    .Q(\hash/p4_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[23]$_DFF_P_  (.D(\hash/p4[23] ),
    .Q(\hash/p4_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[24]$_DFF_P_  (.D(\hash/p4[24] ),
    .Q(\hash/p4_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[25]$_DFF_P_  (.D(\hash/p4[25] ),
    .Q(\hash/p4_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[26]$_DFF_P_  (.D(\hash/p4[26] ),
    .Q(\hash/p4_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[27]$_DFF_P_  (.D(\hash/p4[27] ),
    .Q(\hash/p4_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[28]$_DFF_P_  (.D(\hash/p4[28] ),
    .Q(\hash/p4_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[29]$_DFF_P_  (.D(\hash/p4[29] ),
    .Q(\hash/p4_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[2]$_DFF_P_  (.D(\hash/p4[2] ),
    .Q(\hash/p4_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[30]$_DFF_P_  (.D(\hash/p4[30] ),
    .Q(\hash/p4_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[31]$_DFF_P_  (.D(\hash/p4[31] ),
    .Q(\hash/p4_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[3]$_DFF_P_  (.D(\hash/p4[3] ),
    .Q(\hash/p4_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[4]$_DFF_P_  (.D(\hash/p4[4] ),
    .Q(\hash/p4_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[5]$_DFF_P_  (.D(\hash/p4[5] ),
    .Q(\hash/p4_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[6]$_DFF_P_  (.D(\hash/p4[6] ),
    .Q(\hash/p4_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[7]$_DFF_P_  (.D(\hash/p4[7] ),
    .Q(\hash/p4_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[8]$_DFF_P_  (.D(\hash/p4[8] ),
    .Q(\hash/p4_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p4_cap[9]$_DFF_P_  (.D(\hash/p4[9] ),
    .Q(\hash/p4_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[0]$_DFF_P_  (.D(\hash/p5[0] ),
    .Q(\hash/p5_cap[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[10]$_DFF_P_  (.D(\hash/p5[10] ),
    .Q(\hash/p5_cap[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[11]$_DFF_P_  (.D(\hash/p5[11] ),
    .Q(\hash/p5_cap[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[12]$_DFF_P_  (.D(\hash/p5[12] ),
    .Q(\hash/p5_cap[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[13]$_DFF_P_  (.D(\hash/p5[13] ),
    .Q(\hash/p5_cap[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[14]$_DFF_P_  (.D(\hash/p5[14] ),
    .Q(\hash/p5_cap[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[15]$_DFF_P_  (.D(\hash/p5[15] ),
    .Q(\hash/p5_cap[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[16]$_DFF_P_  (.D(\hash/p5[16] ),
    .Q(\hash/p5_cap[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[17]$_DFF_P_  (.D(\hash/p5[17] ),
    .Q(\hash/p5_cap[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[18]$_DFF_P_  (.D(\hash/p5[18] ),
    .Q(\hash/p5_cap[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[19]$_DFF_P_  (.D(\hash/p5[19] ),
    .Q(\hash/p5_cap[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[1]$_DFF_P_  (.D(\hash/p5[1] ),
    .Q(\hash/p5_cap[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[20]$_DFF_P_  (.D(\hash/p5[20] ),
    .Q(\hash/p5_cap[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[21]$_DFF_P_  (.D(\hash/p5[21] ),
    .Q(\hash/p5_cap[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[22]$_DFF_P_  (.D(\hash/p5[22] ),
    .Q(\hash/p5_cap[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[23]$_DFF_P_  (.D(\hash/p5[23] ),
    .Q(\hash/p5_cap[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[24]$_DFF_P_  (.D(\hash/p5[24] ),
    .Q(\hash/p5_cap[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[25]$_DFF_P_  (.D(\hash/p5[25] ),
    .Q(\hash/p5_cap[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[26]$_DFF_P_  (.D(\hash/p5[26] ),
    .Q(\hash/p5_cap[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[27]$_DFF_P_  (.D(\hash/p5[27] ),
    .Q(\hash/p5_cap[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[28]$_DFF_P_  (.D(\hash/p5[28] ),
    .Q(\hash/p5_cap[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[29]$_DFF_P_  (.D(\hash/p5[29] ),
    .Q(\hash/p5_cap[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[2]$_DFF_P_  (.D(\hash/p5[2] ),
    .Q(\hash/p5_cap[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[30]$_DFF_P_  (.D(\hash/p5[30] ),
    .Q(\hash/p5_cap[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[31]$_DFF_P_  (.D(\hash/p5[31] ),
    .Q(\hash/p5_cap[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[3]$_DFF_P_  (.D(\hash/p5[3] ),
    .Q(\hash/p5_cap[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[4]$_DFF_P_  (.D(\hash/p5[4] ),
    .Q(\hash/p5_cap[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[5]$_DFF_P_  (.D(\hash/p5[5] ),
    .Q(\hash/p5_cap[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[6]$_DFF_P_  (.D(\hash/p5[6] ),
    .Q(\hash/p5_cap[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[7]$_DFF_P_  (.D(\hash/p5[7] ),
    .Q(\hash/p5_cap[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[8]$_DFF_P_  (.D(\hash/p5[8] ),
    .Q(\hash/p5_cap[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \hash/p5_cap[9]$_DFF_P_  (.D(\hash/p5[9] ),
    .Q(\hash/p5_cap[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[0]$_SDFF_PP0_  (.D(_00720_),
    .Q(\k_value1[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[10]$_SDFF_PP1_  (.D(_00721_),
    .Q(\k_value1[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[11]$_SDFF_PP1_  (.D(_00722_),
    .Q(\k_value1[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[12]$_SDFF_PP0_  (.D(_00723_),
    .Q(\k_value1[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[13]$_SDFF_PP1_  (.D(_00724_),
    .Q(\k_value1[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[14]$_SDFF_PP0_  (.D(_00725_),
    .Q(\k_value1[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[15]$_SDFF_PP0_  (.D(_00726_),
    .Q(\k_value1[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[16]$_SDFF_PP0_  (.D(_00727_),
    .Q(\k_value1[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[17]$_SDFF_PP1_  (.D(_00728_),
    .Q(\k_value1[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[18]$_SDFF_PP0_  (.D(_00729_),
    .Q(\k_value1[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[19]$_SDFF_PP1_  (.D(_00730_),
    .Q(\k_value1[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[1]$_SDFF_PP0_  (.D(_00731_),
    .Q(\k_value1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[20]$_SDFF_PP0_  (.D(_00732_),
    .Q(\k_value1[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[21]$_SDFF_PP0_  (.D(_00733_),
    .Q(\k_value1[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[22]$_SDFF_PP0_  (.D(_00734_),
    .Q(\k_value1[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[23]$_SDFF_PP1_  (.D(_00735_),
    .Q(\k_value1[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[24]$_SDFF_PP0_  (.D(_00736_),
    .Q(\k_value1[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[25]$_SDFF_PP1_  (.D(_00737_),
    .Q(\k_value1[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[26]$_SDFF_PP0_  (.D(_00738_),
    .Q(\k_value1[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[27]$_SDFF_PP0_  (.D(_00739_),
    .Q(\k_value1[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[28]$_SDFF_PP0_  (.D(_00740_),
    .Q(\k_value1[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[29]$_SDFF_PP0_  (.D(_00741_),
    .Q(\k_value1[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[2]$_SDFF_PP0_  (.D(_00742_),
    .Q(\k_value1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[30]$_SDFF_PP1_  (.D(_00743_),
    .Q(\k_value1[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[31]$_SDFF_PP0_  (.D(_00744_),
    .Q(\k_value1[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[3]$_SDFF_PP1_  (.D(_00745_),
    .Q(\k_value1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[4]$_SDFF_PP1_  (.D(_00746_),
    .Q(\k_value1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[5]$_SDFF_PP0_  (.D(_00747_),
    .Q(\k_value1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[6]$_SDFF_PP0_  (.D(_00748_),
    .Q(\k_value1[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[7]$_SDFF_PP1_  (.D(_00749_),
    .Q(\k_value1[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[8]$_SDFF_PP1_  (.D(_00750_),
    .Q(\k_value1[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[9]$_SDFF_PP1_  (.D(_00751_),
    .Q(\k_value1[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[0]$_SDFF_PP1_  (.D(_00752_),
    .Q(\k_value2[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[10]$_SDFF_PP1_  (.D(_00753_),
    .Q(\k_value2[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[11]$_SDFF_PP0_  (.D(_00754_),
    .Q(\k_value2[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[12]$_SDFF_PP0_  (.D(_00755_),
    .Q(\k_value2[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[13]$_SDFF_PP0_  (.D(_00756_),
    .Q(\k_value2[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[14]$_SDFF_PP1_  (.D(_00757_),
    .Q(\k_value2[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[15]$_SDFF_PP0_  (.D(_00758_),
    .Q(\k_value2[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[16]$_SDFF_PP1_  (.D(_00759_),
    .Q(\k_value2[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[17]$_SDFF_PP1_  (.D(_00760_),
    .Q(\k_value2[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[18]$_SDFF_PP1_  (.D(_00761_),
    .Q(\k_value2[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[19]$_SDFF_PP0_  (.D(_00762_),
    .Q(\k_value2[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[1]$_SDFF_PP0_  (.D(_00763_),
    .Q(\k_value2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[20]$_SDFF_PP1_  (.D(_00764_),
    .Q(\k_value2[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[21]$_SDFF_PP1_  (.D(_00765_),
    .Q(\k_value2[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[22]$_SDFF_PP0_  (.D(_00766_),
    .Q(\k_value2[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[23]$_SDFF_PP0_  (.D(_00767_),
    .Q(\k_value2[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[24]$_SDFF_PP1_  (.D(_00768_),
    .Q(\k_value2[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[25]$_SDFF_PP0_  (.D(_00769_),
    .Q(\k_value2[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[26]$_SDFF_PP0_  (.D(_00770_),
    .Q(\k_value2[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[27]$_SDFF_PP0_  (.D(_00771_),
    .Q(\k_value2[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[28]$_SDFF_PP1_  (.D(_00772_),
    .Q(\k_value2[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[29]$_SDFF_PP1_  (.D(_00773_),
    .Q(\k_value2[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[2]$_SDFF_PP0_  (.D(_00774_),
    .Q(\k_value2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[30]$_SDFF_PP1_  (.D(_00775_),
    .Q(\k_value2[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[31]$_SDFF_PP0_  (.D(_00776_),
    .Q(\k_value2[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[3]$_SDFF_PP0_  (.D(_00777_),
    .Q(\k_value2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[4]$_SDFF_PP1_  (.D(_00778_),
    .Q(\k_value2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[5]$_SDFF_PP0_  (.D(_00779_),
    .Q(\k_value2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[6]$_SDFF_PP0_  (.D(_00780_),
    .Q(\k_value2[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[7]$_SDFF_PP1_  (.D(_00781_),
    .Q(\k_value2[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[8]$_SDFF_PP0_  (.D(_00782_),
    .Q(\k_value2[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[9]$_SDFF_PP0_  (.D(_00783_),
    .Q(\k_value2[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \ready$_DFF_P_  (.D(ready_dash),
    .Q(ready),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \ready_dash$_SDFF_PP0_  (.D(_00784_),
    .Q(ready_dash),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_2 \reset_hash$_DFF_P_  (.D(reset),
    .Q(reset_hash),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_4 \reset_hash_dash$_DFF_P_  (.D(reset_hash),
    .Q(reset_hash_dash),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][0]$_DFFE_PP_  (.D(_00129_),
    .DE(_00127_),
    .Q(\w[0][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][10]$_DFFE_PP_  (.D(_00130_),
    .DE(_00127_),
    .Q(\w[0][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][11]$_DFFE_PP_  (.D(_00131_),
    .DE(_00127_),
    .Q(\w[0][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][12]$_DFFE_PP_  (.D(_00132_),
    .DE(_00127_),
    .Q(\w[0][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][13]$_DFFE_PP_  (.D(_00133_),
    .DE(_00127_),
    .Q(\w[0][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][14]$_DFFE_PP_  (.D(_00134_),
    .DE(_00127_),
    .Q(\w[0][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][15]$_DFFE_PP_  (.D(_00135_),
    .DE(_00127_),
    .Q(\w[0][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][16]$_DFFE_PP_  (.D(_00136_),
    .DE(_00127_),
    .Q(\w[0][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][17]$_DFFE_PP_  (.D(_00137_),
    .DE(_00127_),
    .Q(\w[0][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][18]$_DFFE_PP_  (.D(_00138_),
    .DE(_00127_),
    .Q(\w[0][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][19]$_DFFE_PP_  (.D(_00139_),
    .DE(_00127_),
    .Q(\w[0][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][1]$_DFFE_PP_  (.D(_00140_),
    .DE(_00127_),
    .Q(\w[0][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][20]$_DFFE_PP_  (.D(_00141_),
    .DE(_00127_),
    .Q(\w[0][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][21]$_DFFE_PP_  (.D(_00142_),
    .DE(_00127_),
    .Q(\w[0][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][22]$_DFFE_PP_  (.D(_00143_),
    .DE(_00127_),
    .Q(\w[0][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][23]$_DFFE_PP_  (.D(_00144_),
    .DE(_00127_),
    .Q(\w[0][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][24]$_DFFE_PP_  (.D(_00145_),
    .DE(_00127_),
    .Q(\w[0][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][25]$_DFFE_PP_  (.D(_00146_),
    .DE(_00127_),
    .Q(\w[0][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][26]$_DFFE_PP_  (.D(_00147_),
    .DE(_00127_),
    .Q(\w[0][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][27]$_DFFE_PP_  (.D(_00148_),
    .DE(_00127_),
    .Q(\w[0][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][28]$_DFFE_PP_  (.D(_00149_),
    .DE(_00127_),
    .Q(\w[0][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][29]$_DFFE_PP_  (.D(_00150_),
    .DE(_00127_),
    .Q(\w[0][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][2]$_DFFE_PP_  (.D(_00151_),
    .DE(_00127_),
    .Q(\w[0][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][30]$_DFFE_PP_  (.D(_00152_),
    .DE(_00127_),
    .Q(\w[0][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][31]$_DFFE_PP_  (.D(_00153_),
    .DE(_00127_),
    .Q(\w[0][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][3]$_DFFE_PP_  (.D(_00154_),
    .DE(_00127_),
    .Q(\w[0][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][4]$_DFFE_PP_  (.D(_00155_),
    .DE(_00127_),
    .Q(\w[0][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][5]$_DFFE_PP_  (.D(_00156_),
    .DE(_00127_),
    .Q(\w[0][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][6]$_DFFE_PP_  (.D(_00157_),
    .DE(_00127_),
    .Q(\w[0][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][7]$_DFFE_PP_  (.D(_00158_),
    .DE(_00127_),
    .Q(\w[0][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][8]$_DFFE_PP_  (.D(_00159_),
    .DE(_00127_),
    .Q(\w[0][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][9]$_DFFE_PP_  (.D(_00160_),
    .DE(_00127_),
    .Q(\w[0][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][0]$_DFFE_PP_  (.D(_00161_),
    .DE(_00126_),
    .Q(\w[10][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][10]$_DFFE_PP_  (.D(_00162_),
    .DE(_00126_),
    .Q(\w[10][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][11]$_DFFE_PP_  (.D(_00163_),
    .DE(_00126_),
    .Q(\w[10][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][12]$_DFFE_PP_  (.D(_00164_),
    .DE(_00126_),
    .Q(\w[10][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][13]$_DFFE_PP_  (.D(_00165_),
    .DE(_00126_),
    .Q(\w[10][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][14]$_DFFE_PP_  (.D(_00166_),
    .DE(_00126_),
    .Q(\w[10][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][15]$_DFFE_PP_  (.D(_00167_),
    .DE(_00126_),
    .Q(\w[10][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][16]$_DFFE_PP_  (.D(_00168_),
    .DE(_00126_),
    .Q(\w[10][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][17]$_DFFE_PP_  (.D(_00169_),
    .DE(_00126_),
    .Q(\w[10][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][18]$_DFFE_PP_  (.D(_00170_),
    .DE(_00126_),
    .Q(\w[10][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][19]$_DFFE_PP_  (.D(_00171_),
    .DE(_00126_),
    .Q(\w[10][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][1]$_DFFE_PP_  (.D(_00172_),
    .DE(_00126_),
    .Q(\w[10][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][20]$_DFFE_PP_  (.D(_00173_),
    .DE(_00126_),
    .Q(\w[10][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][21]$_DFFE_PP_  (.D(_00174_),
    .DE(_00126_),
    .Q(\w[10][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][22]$_DFFE_PP_  (.D(_00175_),
    .DE(_00126_),
    .Q(\w[10][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][23]$_DFFE_PP_  (.D(_00176_),
    .DE(_00126_),
    .Q(\w[10][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][24]$_DFFE_PP_  (.D(_00177_),
    .DE(_00126_),
    .Q(\w[10][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][25]$_DFFE_PP_  (.D(_00178_),
    .DE(_00126_),
    .Q(\w[10][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][26]$_DFFE_PP_  (.D(_00179_),
    .DE(_00126_),
    .Q(\w[10][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][27]$_DFFE_PP_  (.D(_00180_),
    .DE(_00126_),
    .Q(\w[10][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][28]$_DFFE_PP_  (.D(_00181_),
    .DE(_00126_),
    .Q(\w[10][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][29]$_DFFE_PP_  (.D(_00182_),
    .DE(_00126_),
    .Q(\w[10][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][2]$_DFFE_PP_  (.D(_00183_),
    .DE(_00126_),
    .Q(\w[10][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][30]$_DFFE_PP_  (.D(_00184_),
    .DE(_00126_),
    .Q(\w[10][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][31]$_DFFE_PP_  (.D(_00185_),
    .DE(_00126_),
    .Q(\w[10][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][3]$_DFFE_PP_  (.D(_00186_),
    .DE(_00126_),
    .Q(\w[10][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][4]$_DFFE_PP_  (.D(_00187_),
    .DE(_00126_),
    .Q(\w[10][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][5]$_DFFE_PP_  (.D(_00188_),
    .DE(_00126_),
    .Q(\w[10][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][6]$_DFFE_PP_  (.D(_00189_),
    .DE(_00126_),
    .Q(\w[10][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][7]$_DFFE_PP_  (.D(_00190_),
    .DE(_00126_),
    .Q(\w[10][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][8]$_DFFE_PP_  (.D(_00191_),
    .DE(_00126_),
    .Q(\w[10][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][9]$_DFFE_PP_  (.D(_00192_),
    .DE(_00126_),
    .Q(\w[10][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][0]$_DFFE_PP_  (.D(_00193_),
    .DE(_00095_),
    .Q(\w[11][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][10]$_DFFE_PP_  (.D(_00194_),
    .DE(_00095_),
    .Q(\w[11][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][11]$_DFFE_PP_  (.D(_00195_),
    .DE(_00095_),
    .Q(\w[11][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][12]$_DFFE_PP_  (.D(_00196_),
    .DE(_00095_),
    .Q(\w[11][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][13]$_DFFE_PP_  (.D(_00197_),
    .DE(_00095_),
    .Q(\w[11][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][14]$_DFFE_PP_  (.D(_00198_),
    .DE(_00095_),
    .Q(\w[11][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][15]$_DFFE_PP_  (.D(_00199_),
    .DE(_00095_),
    .Q(\w[11][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][16]$_DFFE_PP_  (.D(_00200_),
    .DE(_00095_),
    .Q(\w[11][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][17]$_DFFE_PP_  (.D(_00201_),
    .DE(_00095_),
    .Q(\w[11][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][18]$_DFFE_PP_  (.D(_00202_),
    .DE(_00095_),
    .Q(\w[11][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][19]$_DFFE_PP_  (.D(_00203_),
    .DE(_00095_),
    .Q(\w[11][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][1]$_DFFE_PP_  (.D(_00204_),
    .DE(_00095_),
    .Q(\w[11][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][20]$_DFFE_PP_  (.D(_00205_),
    .DE(_00095_),
    .Q(\w[11][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][21]$_DFFE_PP_  (.D(_00206_),
    .DE(_00095_),
    .Q(\w[11][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][22]$_DFFE_PP_  (.D(_00207_),
    .DE(_00095_),
    .Q(\w[11][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][23]$_DFFE_PP_  (.D(_00208_),
    .DE(_00095_),
    .Q(\w[11][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][24]$_DFFE_PP_  (.D(_00209_),
    .DE(_00095_),
    .Q(\w[11][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][25]$_DFFE_PP_  (.D(_00210_),
    .DE(_00095_),
    .Q(\w[11][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][26]$_DFFE_PP_  (.D(_00211_),
    .DE(_00095_),
    .Q(\w[11][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][27]$_DFFE_PP_  (.D(_00212_),
    .DE(_00095_),
    .Q(\w[11][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][28]$_DFFE_PP_  (.D(_00213_),
    .DE(_00095_),
    .Q(\w[11][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][29]$_DFFE_PP_  (.D(_00214_),
    .DE(_00095_),
    .Q(\w[11][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][2]$_DFFE_PP_  (.D(_00215_),
    .DE(_00095_),
    .Q(\w[11][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][30]$_DFFE_PP_  (.D(_00216_),
    .DE(_00095_),
    .Q(\w[11][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][31]$_DFFE_PP_  (.D(_00217_),
    .DE(_00095_),
    .Q(\w[11][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][3]$_DFFE_PP_  (.D(_00218_),
    .DE(_00095_),
    .Q(\w[11][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][4]$_DFFE_PP_  (.D(_00219_),
    .DE(_00095_),
    .Q(\w[11][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][5]$_DFFE_PP_  (.D(_00220_),
    .DE(_00095_),
    .Q(\w[11][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][6]$_DFFE_PP_  (.D(_00221_),
    .DE(_00095_),
    .Q(\w[11][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][7]$_DFFE_PP_  (.D(_00222_),
    .DE(_00095_),
    .Q(\w[11][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][8]$_DFFE_PP_  (.D(_00223_),
    .DE(_00095_),
    .Q(\w[11][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][9]$_DFFE_PP_  (.D(_00224_),
    .DE(_00095_),
    .Q(\w[11][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][0]$_DFFE_PP_  (.D(_00225_),
    .DE(_00125_),
    .Q(\w[12][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][10]$_DFFE_PP_  (.D(_00226_),
    .DE(_00125_),
    .Q(\w[12][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][11]$_DFFE_PP_  (.D(_00227_),
    .DE(_00125_),
    .Q(\w[12][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][12]$_DFFE_PP_  (.D(_00228_),
    .DE(_00125_),
    .Q(\w[12][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][13]$_DFFE_PP_  (.D(_00229_),
    .DE(_00125_),
    .Q(\w[12][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][14]$_DFFE_PP_  (.D(_00230_),
    .DE(_00125_),
    .Q(\w[12][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][15]$_DFFE_PP_  (.D(_00231_),
    .DE(_00125_),
    .Q(\w[12][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][16]$_DFFE_PP_  (.D(_00232_),
    .DE(_00125_),
    .Q(\w[12][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][17]$_DFFE_PP_  (.D(_00233_),
    .DE(_00125_),
    .Q(\w[12][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][18]$_DFFE_PP_  (.D(_00234_),
    .DE(_00125_),
    .Q(\w[12][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][19]$_DFFE_PP_  (.D(_00235_),
    .DE(_00125_),
    .Q(\w[12][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][1]$_DFFE_PP_  (.D(_00236_),
    .DE(_00125_),
    .Q(\w[12][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][20]$_DFFE_PP_  (.D(_00237_),
    .DE(_00125_),
    .Q(\w[12][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][21]$_DFFE_PP_  (.D(_00238_),
    .DE(_00125_),
    .Q(\w[12][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][22]$_DFFE_PP_  (.D(_00239_),
    .DE(_00125_),
    .Q(\w[12][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][23]$_DFFE_PP_  (.D(_00240_),
    .DE(_00125_),
    .Q(\w[12][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][24]$_DFFE_PP_  (.D(_00241_),
    .DE(_00125_),
    .Q(\w[12][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][25]$_DFFE_PP_  (.D(_00242_),
    .DE(_00125_),
    .Q(\w[12][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][26]$_DFFE_PP_  (.D(_00243_),
    .DE(_00125_),
    .Q(\w[12][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][27]$_DFFE_PP_  (.D(_00244_),
    .DE(_00125_),
    .Q(\w[12][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][28]$_DFFE_PP_  (.D(_00245_),
    .DE(_00125_),
    .Q(\w[12][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][29]$_DFFE_PP_  (.D(_00246_),
    .DE(_00125_),
    .Q(\w[12][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][2]$_DFFE_PP_  (.D(_00247_),
    .DE(_00125_),
    .Q(\w[12][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][30]$_DFFE_PP_  (.D(_00248_),
    .DE(_00125_),
    .Q(\w[12][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][31]$_DFFE_PP_  (.D(_00249_),
    .DE(_00125_),
    .Q(\w[12][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][3]$_DFFE_PP_  (.D(_00250_),
    .DE(_00125_),
    .Q(\w[12][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][4]$_DFFE_PP_  (.D(_00251_),
    .DE(_00125_),
    .Q(\w[12][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][5]$_DFFE_PP_  (.D(_00252_),
    .DE(_00125_),
    .Q(\w[12][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][6]$_DFFE_PP_  (.D(_00253_),
    .DE(_00125_),
    .Q(\w[12][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][7]$_DFFE_PP_  (.D(_00254_),
    .DE(_00125_),
    .Q(\w[12][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][8]$_DFFE_PP_  (.D(_00255_),
    .DE(_00125_),
    .Q(\w[12][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][9]$_DFFE_PP_  (.D(_00256_),
    .DE(_00125_),
    .Q(\w[12][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][0]$_DFFE_PP_  (.D(_00257_),
    .DE(_00094_),
    .Q(\w[13][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][10]$_DFFE_PP_  (.D(_00258_),
    .DE(_00094_),
    .Q(\w[13][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][11]$_DFFE_PP_  (.D(_00259_),
    .DE(_00094_),
    .Q(\w[13][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][12]$_DFFE_PP_  (.D(_00260_),
    .DE(_00094_),
    .Q(\w[13][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][13]$_DFFE_PP_  (.D(_00261_),
    .DE(_00094_),
    .Q(\w[13][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][14]$_DFFE_PP_  (.D(_00262_),
    .DE(_00094_),
    .Q(\w[13][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][15]$_DFFE_PP_  (.D(_00263_),
    .DE(_00094_),
    .Q(\w[13][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][16]$_DFFE_PP_  (.D(_00264_),
    .DE(_00094_),
    .Q(\w[13][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][17]$_DFFE_PP_  (.D(_00265_),
    .DE(_00094_),
    .Q(\w[13][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][18]$_DFFE_PP_  (.D(_00266_),
    .DE(_00094_),
    .Q(\w[13][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][19]$_DFFE_PP_  (.D(_00267_),
    .DE(_00094_),
    .Q(\w[13][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][1]$_DFFE_PP_  (.D(_00268_),
    .DE(_00094_),
    .Q(\w[13][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][20]$_DFFE_PP_  (.D(_00269_),
    .DE(_00094_),
    .Q(\w[13][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][21]$_DFFE_PP_  (.D(_00270_),
    .DE(_00094_),
    .Q(\w[13][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][22]$_DFFE_PP_  (.D(_00271_),
    .DE(_00094_),
    .Q(\w[13][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][23]$_DFFE_PP_  (.D(_00272_),
    .DE(_00094_),
    .Q(\w[13][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][24]$_DFFE_PP_  (.D(_00273_),
    .DE(_00094_),
    .Q(\w[13][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][25]$_DFFE_PP_  (.D(_00274_),
    .DE(_00094_),
    .Q(\w[13][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][26]$_DFFE_PP_  (.D(_00275_),
    .DE(_00094_),
    .Q(\w[13][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][27]$_DFFE_PP_  (.D(_00276_),
    .DE(_00094_),
    .Q(\w[13][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][28]$_DFFE_PP_  (.D(_00277_),
    .DE(_00094_),
    .Q(\w[13][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][29]$_DFFE_PP_  (.D(_00278_),
    .DE(_00094_),
    .Q(\w[13][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][2]$_DFFE_PP_  (.D(_00279_),
    .DE(_00094_),
    .Q(\w[13][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][30]$_DFFE_PP_  (.D(_00280_),
    .DE(_00094_),
    .Q(\w[13][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][31]$_DFFE_PP_  (.D(_00281_),
    .DE(_00094_),
    .Q(\w[13][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][3]$_DFFE_PP_  (.D(_00282_),
    .DE(_00094_),
    .Q(\w[13][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][4]$_DFFE_PP_  (.D(_00283_),
    .DE(_00094_),
    .Q(\w[13][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][5]$_DFFE_PP_  (.D(_00284_),
    .DE(_00094_),
    .Q(\w[13][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][6]$_DFFE_PP_  (.D(_00285_),
    .DE(_00094_),
    .Q(\w[13][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][7]$_DFFE_PP_  (.D(_00286_),
    .DE(_00094_),
    .Q(\w[13][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][8]$_DFFE_PP_  (.D(_00287_),
    .DE(_00094_),
    .Q(\w[13][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][9]$_DFFE_PP_  (.D(_00288_),
    .DE(_00094_),
    .Q(\w[13][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][0]$_DFFE_PP_  (.D(_00289_),
    .DE(_00124_),
    .Q(\w[14][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][10]$_DFFE_PP_  (.D(_00290_),
    .DE(_00124_),
    .Q(\w[14][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][11]$_DFFE_PP_  (.D(_00291_),
    .DE(_00124_),
    .Q(\w[14][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][12]$_DFFE_PP_  (.D(_00292_),
    .DE(_00124_),
    .Q(\w[14][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][13]$_DFFE_PP_  (.D(_00293_),
    .DE(_00124_),
    .Q(\w[14][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][14]$_DFFE_PP_  (.D(_00294_),
    .DE(_00124_),
    .Q(\w[14][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][15]$_DFFE_PP_  (.D(_00295_),
    .DE(_00124_),
    .Q(\w[14][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][16]$_DFFE_PP_  (.D(_00296_),
    .DE(_00124_),
    .Q(\w[14][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][17]$_DFFE_PP_  (.D(_00297_),
    .DE(_00124_),
    .Q(\w[14][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][18]$_DFFE_PP_  (.D(_00298_),
    .DE(_00124_),
    .Q(\w[14][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][19]$_DFFE_PP_  (.D(_00299_),
    .DE(_00124_),
    .Q(\w[14][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][1]$_DFFE_PP_  (.D(_00300_),
    .DE(_00124_),
    .Q(\w[14][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][20]$_DFFE_PP_  (.D(_00301_),
    .DE(_00124_),
    .Q(\w[14][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][21]$_DFFE_PP_  (.D(_00302_),
    .DE(_00124_),
    .Q(\w[14][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][22]$_DFFE_PP_  (.D(_00303_),
    .DE(_00124_),
    .Q(\w[14][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][23]$_DFFE_PP_  (.D(_00304_),
    .DE(_00124_),
    .Q(\w[14][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][24]$_DFFE_PP_  (.D(_00305_),
    .DE(_00124_),
    .Q(\w[14][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][25]$_DFFE_PP_  (.D(_00306_),
    .DE(_00124_),
    .Q(\w[14][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][26]$_DFFE_PP_  (.D(_00307_),
    .DE(_00124_),
    .Q(\w[14][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][27]$_DFFE_PP_  (.D(_00308_),
    .DE(_00124_),
    .Q(\w[14][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][28]$_DFFE_PP_  (.D(_00309_),
    .DE(_00124_),
    .Q(\w[14][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][29]$_DFFE_PP_  (.D(_00310_),
    .DE(_00124_),
    .Q(\w[14][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][2]$_DFFE_PP_  (.D(_00311_),
    .DE(_00124_),
    .Q(\w[14][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][30]$_DFFE_PP_  (.D(_00312_),
    .DE(_00124_),
    .Q(\w[14][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][31]$_DFFE_PP_  (.D(_00313_),
    .DE(_00124_),
    .Q(\w[14][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][3]$_DFFE_PP_  (.D(_00314_),
    .DE(_00124_),
    .Q(\w[14][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][4]$_DFFE_PP_  (.D(_00315_),
    .DE(_00124_),
    .Q(\w[14][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][5]$_DFFE_PP_  (.D(_00316_),
    .DE(_00124_),
    .Q(\w[14][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][6]$_DFFE_PP_  (.D(_00317_),
    .DE(_00124_),
    .Q(\w[14][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][7]$_DFFE_PP_  (.D(_00318_),
    .DE(_00124_),
    .Q(\w[14][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][8]$_DFFE_PP_  (.D(_00319_),
    .DE(_00124_),
    .Q(\w[14][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][9]$_DFFE_PP_  (.D(_00320_),
    .DE(_00124_),
    .Q(\w[14][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][0]$_DFFE_PP_  (.D(_00321_),
    .DE(_00093_),
    .Q(\w[15][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][10]$_DFFE_PP_  (.D(_00322_),
    .DE(_00093_),
    .Q(\w[15][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][11]$_DFFE_PP_  (.D(_00323_),
    .DE(_00093_),
    .Q(\w[15][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][12]$_DFFE_PP_  (.D(_00324_),
    .DE(_00093_),
    .Q(\w[15][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][13]$_DFFE_PP_  (.D(_00325_),
    .DE(_00093_),
    .Q(\w[15][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][14]$_DFFE_PP_  (.D(_00326_),
    .DE(_00093_),
    .Q(\w[15][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][15]$_DFFE_PP_  (.D(_00327_),
    .DE(_00093_),
    .Q(\w[15][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][16]$_DFFE_PP_  (.D(_00328_),
    .DE(_00093_),
    .Q(\w[15][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][17]$_DFFE_PP_  (.D(_00329_),
    .DE(_00093_),
    .Q(\w[15][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][18]$_DFFE_PP_  (.D(_00330_),
    .DE(_00093_),
    .Q(\w[15][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][19]$_DFFE_PP_  (.D(_00331_),
    .DE(_00093_),
    .Q(\w[15][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][1]$_DFFE_PP_  (.D(_00332_),
    .DE(_00093_),
    .Q(\w[15][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][20]$_DFFE_PP_  (.D(_00333_),
    .DE(_00093_),
    .Q(\w[15][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][21]$_DFFE_PP_  (.D(_00334_),
    .DE(_00093_),
    .Q(\w[15][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][22]$_DFFE_PP_  (.D(_00335_),
    .DE(_00093_),
    .Q(\w[15][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][23]$_DFFE_PP_  (.D(_00336_),
    .DE(_00093_),
    .Q(\w[15][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][24]$_DFFE_PP_  (.D(_00337_),
    .DE(_00093_),
    .Q(\w[15][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][25]$_DFFE_PP_  (.D(_00338_),
    .DE(_00093_),
    .Q(\w[15][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][26]$_DFFE_PP_  (.D(_00339_),
    .DE(_00093_),
    .Q(\w[15][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][27]$_DFFE_PP_  (.D(_00340_),
    .DE(_00093_),
    .Q(\w[15][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][28]$_DFFE_PP_  (.D(_00341_),
    .DE(_00093_),
    .Q(\w[15][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][29]$_DFFE_PP_  (.D(_00342_),
    .DE(_00093_),
    .Q(\w[15][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][2]$_DFFE_PP_  (.D(_00343_),
    .DE(_00093_),
    .Q(\w[15][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][30]$_DFFE_PP_  (.D(_00344_),
    .DE(_00093_),
    .Q(\w[15][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][31]$_DFFE_PP_  (.D(_00345_),
    .DE(_00093_),
    .Q(\w[15][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][3]$_DFFE_PP_  (.D(_00346_),
    .DE(_00093_),
    .Q(\w[15][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][4]$_DFFE_PP_  (.D(_00347_),
    .DE(_00093_),
    .Q(\w[15][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][5]$_DFFE_PP_  (.D(_00348_),
    .DE(_00093_),
    .Q(\w[15][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][6]$_DFFE_PP_  (.D(_00349_),
    .DE(_00093_),
    .Q(\w[15][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][7]$_DFFE_PP_  (.D(_00350_),
    .DE(_00093_),
    .Q(\w[15][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][8]$_DFFE_PP_  (.D(_00351_),
    .DE(_00093_),
    .Q(\w[15][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][9]$_DFFE_PP_  (.D(_00352_),
    .DE(_00093_),
    .Q(\w[15][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][0]$_SDFFCE_PN0P_  (.D(_00785_),
    .DE(_00123_),
    .Q(\w[16][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][10]$_SDFFCE_PN0P_  (.D(_00786_),
    .DE(_00123_),
    .Q(\w[16][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][11]$_SDFFCE_PN0P_  (.D(_00787_),
    .DE(_00123_),
    .Q(\w[16][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][12]$_SDFFCE_PN0P_  (.D(_00788_),
    .DE(_00123_),
    .Q(\w[16][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][13]$_SDFFCE_PN0P_  (.D(_00789_),
    .DE(_00123_),
    .Q(\w[16][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][14]$_SDFFCE_PN0P_  (.D(_00790_),
    .DE(_00123_),
    .Q(\w[16][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][15]$_SDFFCE_PN0P_  (.D(_00791_),
    .DE(_00123_),
    .Q(\w[16][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][16]$_SDFFCE_PN0P_  (.D(_00792_),
    .DE(_00123_),
    .Q(\w[16][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][17]$_SDFFCE_PN0P_  (.D(_00793_),
    .DE(_00123_),
    .Q(\w[16][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][18]$_SDFFCE_PN0P_  (.D(_00794_),
    .DE(_00123_),
    .Q(\w[16][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][19]$_SDFFCE_PN0P_  (.D(_00795_),
    .DE(_00123_),
    .Q(\w[16][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][1]$_SDFFCE_PN0P_  (.D(_00796_),
    .DE(_00123_),
    .Q(\w[16][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][20]$_SDFFCE_PN0P_  (.D(_00797_),
    .DE(_00123_),
    .Q(\w[16][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][21]$_SDFFCE_PN0P_  (.D(_00798_),
    .DE(_00123_),
    .Q(\w[16][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][22]$_SDFFCE_PN0P_  (.D(_00799_),
    .DE(_00123_),
    .Q(\w[16][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][23]$_SDFFCE_PN0P_  (.D(_00800_),
    .DE(_00123_),
    .Q(\w[16][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][24]$_SDFFCE_PN0P_  (.D(_00801_),
    .DE(_00123_),
    .Q(\w[16][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][25]$_SDFFCE_PN0P_  (.D(_00802_),
    .DE(_00123_),
    .Q(\w[16][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][26]$_SDFFCE_PN0P_  (.D(_00803_),
    .DE(_00123_),
    .Q(\w[16][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][27]$_SDFFCE_PN0P_  (.D(_00804_),
    .DE(_00123_),
    .Q(\w[16][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][28]$_SDFFCE_PN0P_  (.D(_00805_),
    .DE(_00123_),
    .Q(\w[16][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][29]$_SDFFCE_PN0P_  (.D(_00806_),
    .DE(_00123_),
    .Q(\w[16][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][2]$_SDFFCE_PN0P_  (.D(_00807_),
    .DE(_00123_),
    .Q(\w[16][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][30]$_SDFFCE_PN0P_  (.D(_00808_),
    .DE(_00123_),
    .Q(\w[16][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][31]$_SDFFCE_PN0P_  (.D(_00809_),
    .DE(_00123_),
    .Q(\w[16][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][3]$_SDFFCE_PN0P_  (.D(_00810_),
    .DE(_00123_),
    .Q(\w[16][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][4]$_SDFFCE_PN0P_  (.D(_00811_),
    .DE(_00123_),
    .Q(\w[16][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][5]$_SDFFCE_PN0P_  (.D(_00812_),
    .DE(_00123_),
    .Q(\w[16][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][6]$_SDFFCE_PN0P_  (.D(_00813_),
    .DE(_00123_),
    .Q(\w[16][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][7]$_SDFFCE_PN0P_  (.D(_00814_),
    .DE(_00123_),
    .Q(\w[16][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][8]$_SDFFCE_PN0P_  (.D(_00815_),
    .DE(_00123_),
    .Q(\w[16][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][9]$_SDFFCE_PN0P_  (.D(_00816_),
    .DE(_00123_),
    .Q(\w[16][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][0]$_SDFFCE_PN0P_  (.D(_00817_),
    .DE(_00092_),
    .Q(\w[17][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][10]$_SDFFCE_PN0P_  (.D(_00818_),
    .DE(_00092_),
    .Q(\w[17][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][11]$_SDFFCE_PN0P_  (.D(_00819_),
    .DE(_00092_),
    .Q(\w[17][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][12]$_SDFFCE_PN0P_  (.D(_00820_),
    .DE(_00092_),
    .Q(\w[17][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][13]$_SDFFCE_PN0P_  (.D(_00821_),
    .DE(_00092_),
    .Q(\w[17][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][14]$_SDFFCE_PN0P_  (.D(_00822_),
    .DE(_00092_),
    .Q(\w[17][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][15]$_SDFFCE_PN0P_  (.D(_00823_),
    .DE(_00092_),
    .Q(\w[17][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][16]$_SDFFCE_PN0P_  (.D(_00824_),
    .DE(_00092_),
    .Q(\w[17][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][17]$_SDFFCE_PN0P_  (.D(_00825_),
    .DE(_00092_),
    .Q(\w[17][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][18]$_SDFFCE_PN0P_  (.D(_00826_),
    .DE(_00092_),
    .Q(\w[17][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][19]$_SDFFCE_PN0P_  (.D(_00827_),
    .DE(_00092_),
    .Q(\w[17][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][1]$_SDFFCE_PN0P_  (.D(_00828_),
    .DE(_00092_),
    .Q(\w[17][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][20]$_SDFFCE_PN0P_  (.D(_00829_),
    .DE(_00092_),
    .Q(\w[17][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][21]$_SDFFCE_PN0P_  (.D(_00830_),
    .DE(_00092_),
    .Q(\w[17][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][22]$_SDFFCE_PN0P_  (.D(_00831_),
    .DE(_00092_),
    .Q(\w[17][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][23]$_SDFFCE_PN0P_  (.D(_00832_),
    .DE(_00092_),
    .Q(\w[17][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][24]$_SDFFCE_PN0P_  (.D(_00833_),
    .DE(_00092_),
    .Q(\w[17][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][25]$_SDFFCE_PN0P_  (.D(_00834_),
    .DE(_00092_),
    .Q(\w[17][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][26]$_SDFFCE_PN0P_  (.D(_00835_),
    .DE(_00092_),
    .Q(\w[17][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][27]$_SDFFCE_PN0P_  (.D(_00836_),
    .DE(_00092_),
    .Q(\w[17][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][28]$_SDFFCE_PN0P_  (.D(_00837_),
    .DE(_00092_),
    .Q(\w[17][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][29]$_SDFFCE_PN0P_  (.D(_00838_),
    .DE(_00092_),
    .Q(\w[17][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][2]$_SDFFCE_PN0P_  (.D(_00839_),
    .DE(_00092_),
    .Q(\w[17][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][30]$_SDFFCE_PN0P_  (.D(_00840_),
    .DE(_00092_),
    .Q(\w[17][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][31]$_SDFFCE_PN0P_  (.D(_00841_),
    .DE(_00092_),
    .Q(\w[17][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][3]$_SDFFCE_PN0P_  (.D(_00842_),
    .DE(_00092_),
    .Q(\w[17][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][4]$_SDFFCE_PN0P_  (.D(_00843_),
    .DE(_00092_),
    .Q(\w[17][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][5]$_SDFFCE_PN0P_  (.D(_00844_),
    .DE(_00092_),
    .Q(\w[17][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][6]$_SDFFCE_PN0P_  (.D(_00845_),
    .DE(_00092_),
    .Q(\w[17][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][7]$_SDFFCE_PN0P_  (.D(_00846_),
    .DE(_00092_),
    .Q(\w[17][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][8]$_SDFFCE_PN0P_  (.D(_00847_),
    .DE(_00092_),
    .Q(\w[17][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][9]$_SDFFCE_PN0P_  (.D(_00848_),
    .DE(_00092_),
    .Q(\w[17][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][0]$_SDFFCE_PN0P_  (.D(_00849_),
    .DE(_00122_),
    .Q(\w[18][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][10]$_SDFFCE_PN0P_  (.D(_00850_),
    .DE(_00122_),
    .Q(\w[18][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][11]$_SDFFCE_PN0P_  (.D(_00851_),
    .DE(_00122_),
    .Q(\w[18][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][12]$_SDFFCE_PN0P_  (.D(_00852_),
    .DE(_00122_),
    .Q(\w[18][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][13]$_SDFFCE_PN0P_  (.D(_00853_),
    .DE(_00122_),
    .Q(\w[18][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][14]$_SDFFCE_PN0P_  (.D(_00854_),
    .DE(_00122_),
    .Q(\w[18][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][15]$_SDFFCE_PN0P_  (.D(_00855_),
    .DE(_00122_),
    .Q(\w[18][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][16]$_SDFFCE_PN0P_  (.D(_00856_),
    .DE(_00122_),
    .Q(\w[18][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][17]$_SDFFCE_PN0P_  (.D(_00857_),
    .DE(_00122_),
    .Q(\w[18][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][18]$_SDFFCE_PN0P_  (.D(_00858_),
    .DE(_00122_),
    .Q(\w[18][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][19]$_SDFFCE_PN0P_  (.D(_00859_),
    .DE(_00122_),
    .Q(\w[18][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][1]$_SDFFCE_PN0P_  (.D(_00860_),
    .DE(_00122_),
    .Q(\w[18][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][20]$_SDFFCE_PN0P_  (.D(_00861_),
    .DE(_00122_),
    .Q(\w[18][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][21]$_SDFFCE_PN0P_  (.D(_00862_),
    .DE(_00122_),
    .Q(\w[18][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][22]$_SDFFCE_PN0P_  (.D(_00863_),
    .DE(_00122_),
    .Q(\w[18][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][23]$_SDFFCE_PN0P_  (.D(_00864_),
    .DE(_00122_),
    .Q(\w[18][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][24]$_SDFFCE_PN0P_  (.D(_00865_),
    .DE(_00122_),
    .Q(\w[18][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][25]$_SDFFCE_PN0P_  (.D(_00866_),
    .DE(_00122_),
    .Q(\w[18][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][26]$_SDFFCE_PN0P_  (.D(_00867_),
    .DE(_00122_),
    .Q(\w[18][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][27]$_SDFFCE_PN0P_  (.D(_00868_),
    .DE(_00122_),
    .Q(\w[18][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][28]$_SDFFCE_PN0P_  (.D(_00869_),
    .DE(_00122_),
    .Q(\w[18][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][29]$_SDFFCE_PN0P_  (.D(_00870_),
    .DE(_00122_),
    .Q(\w[18][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][2]$_SDFFCE_PN0P_  (.D(_00871_),
    .DE(_00122_),
    .Q(\w[18][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][30]$_SDFFCE_PN0P_  (.D(_00872_),
    .DE(_00122_),
    .Q(\w[18][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][31]$_SDFFCE_PN0P_  (.D(_00873_),
    .DE(_00122_),
    .Q(\w[18][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][3]$_SDFFCE_PN0P_  (.D(_00874_),
    .DE(_00122_),
    .Q(\w[18][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][4]$_SDFFCE_PN0P_  (.D(_00875_),
    .DE(_00122_),
    .Q(\w[18][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][5]$_SDFFCE_PN0P_  (.D(_00876_),
    .DE(_00122_),
    .Q(\w[18][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][6]$_SDFFCE_PN0P_  (.D(_00877_),
    .DE(_00122_),
    .Q(\w[18][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][7]$_SDFFCE_PN0P_  (.D(_00878_),
    .DE(_00122_),
    .Q(\w[18][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][8]$_SDFFCE_PN0P_  (.D(_00879_),
    .DE(_00122_),
    .Q(\w[18][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][9]$_SDFFCE_PN0P_  (.D(_00880_),
    .DE(_00122_),
    .Q(\w[18][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][0]$_SDFFCE_PN0P_  (.D(_00881_),
    .DE(_00091_),
    .Q(\w[19][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][10]$_SDFFCE_PN0P_  (.D(_00882_),
    .DE(_00091_),
    .Q(\w[19][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][11]$_SDFFCE_PN0P_  (.D(_00883_),
    .DE(_00091_),
    .Q(\w[19][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][12]$_SDFFCE_PN0P_  (.D(_00884_),
    .DE(_00091_),
    .Q(\w[19][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][13]$_SDFFCE_PN0P_  (.D(_00885_),
    .DE(_00091_),
    .Q(\w[19][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][14]$_SDFFCE_PN0P_  (.D(_00886_),
    .DE(_00091_),
    .Q(\w[19][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][15]$_SDFFCE_PN0P_  (.D(_00887_),
    .DE(_00091_),
    .Q(\w[19][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][16]$_SDFFCE_PN0P_  (.D(_00888_),
    .DE(_00091_),
    .Q(\w[19][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][17]$_SDFFCE_PN0P_  (.D(_00889_),
    .DE(_00091_),
    .Q(\w[19][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][18]$_SDFFCE_PN0P_  (.D(_00890_),
    .DE(_00091_),
    .Q(\w[19][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][19]$_SDFFCE_PN0P_  (.D(_00891_),
    .DE(_00091_),
    .Q(\w[19][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][1]$_SDFFCE_PN0P_  (.D(_00892_),
    .DE(_00091_),
    .Q(\w[19][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][20]$_SDFFCE_PN0P_  (.D(_00893_),
    .DE(_00091_),
    .Q(\w[19][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][21]$_SDFFCE_PN0P_  (.D(_00894_),
    .DE(_00091_),
    .Q(\w[19][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][22]$_SDFFCE_PN0P_  (.D(_00895_),
    .DE(_00091_),
    .Q(\w[19][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][23]$_SDFFCE_PN0P_  (.D(_00896_),
    .DE(_00091_),
    .Q(\w[19][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][24]$_SDFFCE_PN0P_  (.D(_00897_),
    .DE(_00091_),
    .Q(\w[19][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][25]$_SDFFCE_PN0P_  (.D(_00898_),
    .DE(_00091_),
    .Q(\w[19][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][26]$_SDFFCE_PN0P_  (.D(_00899_),
    .DE(_00091_),
    .Q(\w[19][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][27]$_SDFFCE_PN0P_  (.D(_00900_),
    .DE(_00091_),
    .Q(\w[19][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][28]$_SDFFCE_PN0P_  (.D(_00901_),
    .DE(_00091_),
    .Q(\w[19][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][29]$_SDFFCE_PN0P_  (.D(_00902_),
    .DE(_00091_),
    .Q(\w[19][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][2]$_SDFFCE_PN0P_  (.D(_00903_),
    .DE(_00091_),
    .Q(\w[19][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][30]$_SDFFCE_PN0P_  (.D(_00904_),
    .DE(_00091_),
    .Q(\w[19][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][31]$_SDFFCE_PN0P_  (.D(_00905_),
    .DE(_00091_),
    .Q(\w[19][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][3]$_SDFFCE_PN0P_  (.D(_00906_),
    .DE(_00091_),
    .Q(\w[19][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][4]$_SDFFCE_PN0P_  (.D(_00907_),
    .DE(_00091_),
    .Q(\w[19][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][5]$_SDFFCE_PN0P_  (.D(_00908_),
    .DE(_00091_),
    .Q(\w[19][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][6]$_SDFFCE_PN0P_  (.D(_00909_),
    .DE(_00091_),
    .Q(\w[19][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][7]$_SDFFCE_PN0P_  (.D(_00910_),
    .DE(_00091_),
    .Q(\w[19][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][8]$_SDFFCE_PN0P_  (.D(_00911_),
    .DE(_00091_),
    .Q(\w[19][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][9]$_SDFFCE_PN0P_  (.D(_00912_),
    .DE(_00091_),
    .Q(\w[19][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][0]$_DFFE_PP_  (.D(_00353_),
    .DE(_00090_),
    .Q(\w[1][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][10]$_DFFE_PP_  (.D(_00354_),
    .DE(_00090_),
    .Q(\w[1][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][11]$_DFFE_PP_  (.D(_00355_),
    .DE(_00090_),
    .Q(\w[1][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][12]$_DFFE_PP_  (.D(_00356_),
    .DE(_00090_),
    .Q(\w[1][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][13]$_DFFE_PP_  (.D(_00357_),
    .DE(_00090_),
    .Q(\w[1][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][14]$_DFFE_PP_  (.D(_00358_),
    .DE(_00090_),
    .Q(\w[1][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][15]$_DFFE_PP_  (.D(_00359_),
    .DE(_00090_),
    .Q(\w[1][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][16]$_DFFE_PP_  (.D(_00360_),
    .DE(_00090_),
    .Q(\w[1][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][17]$_DFFE_PP_  (.D(_00361_),
    .DE(_00090_),
    .Q(\w[1][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][18]$_DFFE_PP_  (.D(_00362_),
    .DE(_00090_),
    .Q(\w[1][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][19]$_DFFE_PP_  (.D(_00363_),
    .DE(_00090_),
    .Q(\w[1][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][1]$_DFFE_PP_  (.D(_00364_),
    .DE(_00090_),
    .Q(\w[1][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][20]$_DFFE_PP_  (.D(_00365_),
    .DE(_00090_),
    .Q(\w[1][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][21]$_DFFE_PP_  (.D(_00366_),
    .DE(_00090_),
    .Q(\w[1][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][22]$_DFFE_PP_  (.D(_00367_),
    .DE(_00090_),
    .Q(\w[1][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][23]$_DFFE_PP_  (.D(_00368_),
    .DE(_00090_),
    .Q(\w[1][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][24]$_DFFE_PP_  (.D(_00369_),
    .DE(_00090_),
    .Q(\w[1][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][25]$_DFFE_PP_  (.D(_00370_),
    .DE(_00090_),
    .Q(\w[1][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][26]$_DFFE_PP_  (.D(_00371_),
    .DE(_00090_),
    .Q(\w[1][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][27]$_DFFE_PP_  (.D(_00372_),
    .DE(_00090_),
    .Q(\w[1][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][28]$_DFFE_PP_  (.D(_00373_),
    .DE(_00090_),
    .Q(\w[1][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][29]$_DFFE_PP_  (.D(_00374_),
    .DE(_00090_),
    .Q(\w[1][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][2]$_DFFE_PP_  (.D(_00375_),
    .DE(_00090_),
    .Q(\w[1][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][30]$_DFFE_PP_  (.D(_00376_),
    .DE(_00090_),
    .Q(\w[1][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][31]$_DFFE_PP_  (.D(_00377_),
    .DE(_00090_),
    .Q(\w[1][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][3]$_DFFE_PP_  (.D(_00378_),
    .DE(_00090_),
    .Q(\w[1][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][4]$_DFFE_PP_  (.D(_00379_),
    .DE(_00090_),
    .Q(\w[1][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][5]$_DFFE_PP_  (.D(_00380_),
    .DE(_00090_),
    .Q(\w[1][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][6]$_DFFE_PP_  (.D(_00381_),
    .DE(_00090_),
    .Q(\w[1][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][7]$_DFFE_PP_  (.D(_00382_),
    .DE(_00090_),
    .Q(\w[1][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][8]$_DFFE_PP_  (.D(_00383_),
    .DE(_00090_),
    .Q(\w[1][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][9]$_DFFE_PP_  (.D(_00384_),
    .DE(_00090_),
    .Q(\w[1][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][0]$_SDFFCE_PN0P_  (.D(_00913_),
    .DE(_00121_),
    .Q(\w[20][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][10]$_SDFFCE_PN0P_  (.D(_00914_),
    .DE(_00121_),
    .Q(\w[20][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][11]$_SDFFCE_PN0P_  (.D(_00915_),
    .DE(_00121_),
    .Q(\w[20][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][12]$_SDFFCE_PN0P_  (.D(_00916_),
    .DE(_00121_),
    .Q(\w[20][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][13]$_SDFFCE_PN0P_  (.D(_00917_),
    .DE(_00121_),
    .Q(\w[20][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][14]$_SDFFCE_PN0P_  (.D(_00918_),
    .DE(_00121_),
    .Q(\w[20][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][15]$_SDFFCE_PN0P_  (.D(_00919_),
    .DE(_00121_),
    .Q(\w[20][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][16]$_SDFFCE_PN0P_  (.D(_00920_),
    .DE(_00121_),
    .Q(\w[20][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][17]$_SDFFCE_PN0P_  (.D(_00921_),
    .DE(_00121_),
    .Q(\w[20][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][18]$_SDFFCE_PN0P_  (.D(_00922_),
    .DE(_00121_),
    .Q(\w[20][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][19]$_SDFFCE_PN0P_  (.D(_00923_),
    .DE(_00121_),
    .Q(\w[20][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][1]$_SDFFCE_PN0P_  (.D(_00924_),
    .DE(_00121_),
    .Q(\w[20][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][20]$_SDFFCE_PN0P_  (.D(_00925_),
    .DE(_00121_),
    .Q(\w[20][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][21]$_SDFFCE_PN0P_  (.D(_00926_),
    .DE(_00121_),
    .Q(\w[20][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][22]$_SDFFCE_PN0P_  (.D(_00927_),
    .DE(_00121_),
    .Q(\w[20][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][23]$_SDFFCE_PN0P_  (.D(_00928_),
    .DE(_00121_),
    .Q(\w[20][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][24]$_SDFFCE_PN0P_  (.D(_00929_),
    .DE(_00121_),
    .Q(\w[20][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][25]$_SDFFCE_PN0P_  (.D(_00930_),
    .DE(_00121_),
    .Q(\w[20][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][26]$_SDFFCE_PN0P_  (.D(_00931_),
    .DE(_00121_),
    .Q(\w[20][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][27]$_SDFFCE_PN0P_  (.D(_00932_),
    .DE(_00121_),
    .Q(\w[20][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][28]$_SDFFCE_PN0P_  (.D(_00933_),
    .DE(_00121_),
    .Q(\w[20][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][29]$_SDFFCE_PN0P_  (.D(_00934_),
    .DE(_00121_),
    .Q(\w[20][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][2]$_SDFFCE_PN0P_  (.D(_00935_),
    .DE(_00121_),
    .Q(\w[20][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][30]$_SDFFCE_PN0P_  (.D(_00936_),
    .DE(_00121_),
    .Q(\w[20][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][31]$_SDFFCE_PN0P_  (.D(_00937_),
    .DE(_00121_),
    .Q(\w[20][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][3]$_SDFFCE_PN0P_  (.D(_00938_),
    .DE(_00121_),
    .Q(\w[20][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][4]$_SDFFCE_PN0P_  (.D(_00939_),
    .DE(_00121_),
    .Q(\w[20][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][5]$_SDFFCE_PN0P_  (.D(_00940_),
    .DE(_00121_),
    .Q(\w[20][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][6]$_SDFFCE_PN0P_  (.D(_00941_),
    .DE(_00121_),
    .Q(\w[20][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][7]$_SDFFCE_PN0P_  (.D(_00942_),
    .DE(_00121_),
    .Q(\w[20][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][8]$_SDFFCE_PN0P_  (.D(_00943_),
    .DE(_00121_),
    .Q(\w[20][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][9]$_SDFFCE_PN0P_  (.D(_00944_),
    .DE(_00121_),
    .Q(\w[20][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][0]$_SDFFCE_PN0P_  (.D(_00945_),
    .DE(_00089_),
    .Q(\w[21][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][10]$_SDFFCE_PN0P_  (.D(_00946_),
    .DE(_00089_),
    .Q(\w[21][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][11]$_SDFFCE_PN0P_  (.D(_00947_),
    .DE(_00089_),
    .Q(\w[21][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][12]$_SDFFCE_PN0P_  (.D(_00948_),
    .DE(_00089_),
    .Q(\w[21][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][13]$_SDFFCE_PN0P_  (.D(_00949_),
    .DE(_00089_),
    .Q(\w[21][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][14]$_SDFFCE_PN0P_  (.D(_00950_),
    .DE(_00089_),
    .Q(\w[21][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][15]$_SDFFCE_PN0P_  (.D(_00951_),
    .DE(_00089_),
    .Q(\w[21][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][16]$_SDFFCE_PN0P_  (.D(_00952_),
    .DE(_00089_),
    .Q(\w[21][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][17]$_SDFFCE_PN0P_  (.D(_00953_),
    .DE(_00089_),
    .Q(\w[21][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][18]$_SDFFCE_PN0P_  (.D(_00954_),
    .DE(_00089_),
    .Q(\w[21][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][19]$_SDFFCE_PN0P_  (.D(_00955_),
    .DE(_00089_),
    .Q(\w[21][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][1]$_SDFFCE_PN0P_  (.D(_00956_),
    .DE(_00089_),
    .Q(\w[21][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][20]$_SDFFCE_PN0P_  (.D(_00957_),
    .DE(_00089_),
    .Q(\w[21][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][21]$_SDFFCE_PN0P_  (.D(_00958_),
    .DE(_00089_),
    .Q(\w[21][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][22]$_SDFFCE_PN0P_  (.D(_00959_),
    .DE(_00089_),
    .Q(\w[21][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][23]$_SDFFCE_PN0P_  (.D(_00960_),
    .DE(_00089_),
    .Q(\w[21][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][24]$_SDFFCE_PN0P_  (.D(_00961_),
    .DE(_00089_),
    .Q(\w[21][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][25]$_SDFFCE_PN0P_  (.D(_00962_),
    .DE(_00089_),
    .Q(\w[21][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][26]$_SDFFCE_PN0P_  (.D(_00963_),
    .DE(_00089_),
    .Q(\w[21][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][27]$_SDFFCE_PN0P_  (.D(_00964_),
    .DE(_00089_),
    .Q(\w[21][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][28]$_SDFFCE_PN0P_  (.D(_00965_),
    .DE(_00089_),
    .Q(\w[21][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][29]$_SDFFCE_PN0P_  (.D(_00966_),
    .DE(_00089_),
    .Q(\w[21][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][2]$_SDFFCE_PN0P_  (.D(_00967_),
    .DE(_00089_),
    .Q(\w[21][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][30]$_SDFFCE_PN0P_  (.D(_00968_),
    .DE(_00089_),
    .Q(\w[21][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][31]$_SDFFCE_PN0P_  (.D(_00969_),
    .DE(_00089_),
    .Q(\w[21][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][3]$_SDFFCE_PN0P_  (.D(_00970_),
    .DE(_00089_),
    .Q(\w[21][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][4]$_SDFFCE_PN0P_  (.D(_00971_),
    .DE(_00089_),
    .Q(\w[21][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][5]$_SDFFCE_PN0P_  (.D(_00972_),
    .DE(_00089_),
    .Q(\w[21][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][6]$_SDFFCE_PN0P_  (.D(_00973_),
    .DE(_00089_),
    .Q(\w[21][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][7]$_SDFFCE_PN0P_  (.D(_00974_),
    .DE(_00089_),
    .Q(\w[21][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][8]$_SDFFCE_PN0P_  (.D(_00975_),
    .DE(_00089_),
    .Q(\w[21][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][9]$_SDFFCE_PN0P_  (.D(_00976_),
    .DE(_00089_),
    .Q(\w[21][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][0]$_SDFFCE_PN0P_  (.D(_00977_),
    .DE(_00120_),
    .Q(\w[22][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][10]$_SDFFCE_PN0P_  (.D(_00978_),
    .DE(_00120_),
    .Q(\w[22][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][11]$_SDFFCE_PN0P_  (.D(_00979_),
    .DE(_00120_),
    .Q(\w[22][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][12]$_SDFFCE_PN0P_  (.D(_00980_),
    .DE(_00120_),
    .Q(\w[22][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][13]$_SDFFCE_PN0P_  (.D(_00981_),
    .DE(_00120_),
    .Q(\w[22][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][14]$_SDFFCE_PN0P_  (.D(_00982_),
    .DE(_00120_),
    .Q(\w[22][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][15]$_SDFFCE_PN0P_  (.D(_00983_),
    .DE(_00120_),
    .Q(\w[22][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][16]$_SDFFCE_PN0P_  (.D(_00984_),
    .DE(_00120_),
    .Q(\w[22][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][17]$_SDFFCE_PN0P_  (.D(_00985_),
    .DE(_00120_),
    .Q(\w[22][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][18]$_SDFFCE_PN0P_  (.D(_00986_),
    .DE(_00120_),
    .Q(\w[22][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][19]$_SDFFCE_PN0P_  (.D(_00987_),
    .DE(_00120_),
    .Q(\w[22][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][1]$_SDFFCE_PN0P_  (.D(_00988_),
    .DE(_00120_),
    .Q(\w[22][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][20]$_SDFFCE_PN0P_  (.D(_00989_),
    .DE(_00120_),
    .Q(\w[22][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][21]$_SDFFCE_PN0P_  (.D(_00990_),
    .DE(_00120_),
    .Q(\w[22][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][22]$_SDFFCE_PN0P_  (.D(_00991_),
    .DE(_00120_),
    .Q(\w[22][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][23]$_SDFFCE_PN0P_  (.D(_00992_),
    .DE(_00120_),
    .Q(\w[22][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][24]$_SDFFCE_PN0P_  (.D(_00993_),
    .DE(_00120_),
    .Q(\w[22][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][25]$_SDFFCE_PN0P_  (.D(_00994_),
    .DE(_00120_),
    .Q(\w[22][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][26]$_SDFFCE_PN0P_  (.D(_00995_),
    .DE(_00120_),
    .Q(\w[22][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][27]$_SDFFCE_PN0P_  (.D(_00996_),
    .DE(_00120_),
    .Q(\w[22][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][28]$_SDFFCE_PN0P_  (.D(_00997_),
    .DE(_00120_),
    .Q(\w[22][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][29]$_SDFFCE_PN0P_  (.D(_00998_),
    .DE(_00120_),
    .Q(\w[22][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][2]$_SDFFCE_PN0P_  (.D(_00999_),
    .DE(_00120_),
    .Q(\w[22][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][30]$_SDFFCE_PN0P_  (.D(_01000_),
    .DE(_00120_),
    .Q(\w[22][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][31]$_SDFFCE_PN0P_  (.D(_01001_),
    .DE(_00120_),
    .Q(\w[22][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][3]$_SDFFCE_PN0P_  (.D(_01002_),
    .DE(_00120_),
    .Q(\w[22][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][4]$_SDFFCE_PN0P_  (.D(_01003_),
    .DE(_00120_),
    .Q(\w[22][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][5]$_SDFFCE_PN0P_  (.D(_01004_),
    .DE(_00120_),
    .Q(\w[22][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][6]$_SDFFCE_PN0P_  (.D(_01005_),
    .DE(_00120_),
    .Q(\w[22][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][7]$_SDFFCE_PN0P_  (.D(_01006_),
    .DE(_00120_),
    .Q(\w[22][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][8]$_SDFFCE_PN0P_  (.D(_01007_),
    .DE(_00120_),
    .Q(\w[22][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][9]$_SDFFCE_PN0P_  (.D(_01008_),
    .DE(_00120_),
    .Q(\w[22][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][0]$_SDFFCE_PN0P_  (.D(_01009_),
    .DE(_00088_),
    .Q(\w[23][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][10]$_SDFFCE_PN0P_  (.D(_01010_),
    .DE(_00088_),
    .Q(\w[23][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][11]$_SDFFCE_PN0P_  (.D(_01011_),
    .DE(_00088_),
    .Q(\w[23][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][12]$_SDFFCE_PN0P_  (.D(_01012_),
    .DE(_00088_),
    .Q(\w[23][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][13]$_SDFFCE_PN0P_  (.D(_01013_),
    .DE(_00088_),
    .Q(\w[23][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][14]$_SDFFCE_PN0P_  (.D(_01014_),
    .DE(_00088_),
    .Q(\w[23][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][15]$_SDFFCE_PN0P_  (.D(_01015_),
    .DE(_00088_),
    .Q(\w[23][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][16]$_SDFFCE_PN0P_  (.D(_01016_),
    .DE(_00088_),
    .Q(\w[23][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][17]$_SDFFCE_PN0P_  (.D(_01017_),
    .DE(_00088_),
    .Q(\w[23][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][18]$_SDFFCE_PN0P_  (.D(_01018_),
    .DE(_00088_),
    .Q(\w[23][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][19]$_SDFFCE_PN0P_  (.D(_01019_),
    .DE(_00088_),
    .Q(\w[23][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][1]$_SDFFCE_PN0P_  (.D(_01020_),
    .DE(_00088_),
    .Q(\w[23][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][20]$_SDFFCE_PN0P_  (.D(_01021_),
    .DE(_00088_),
    .Q(\w[23][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][21]$_SDFFCE_PN0P_  (.D(_01022_),
    .DE(_00088_),
    .Q(\w[23][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][22]$_SDFFCE_PN0P_  (.D(_01023_),
    .DE(_00088_),
    .Q(\w[23][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][23]$_SDFFCE_PN0P_  (.D(_01024_),
    .DE(_00088_),
    .Q(\w[23][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][24]$_SDFFCE_PN0P_  (.D(_01025_),
    .DE(_00088_),
    .Q(\w[23][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][25]$_SDFFCE_PN0P_  (.D(_01026_),
    .DE(_00088_),
    .Q(\w[23][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][26]$_SDFFCE_PN0P_  (.D(_01027_),
    .DE(_00088_),
    .Q(\w[23][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][27]$_SDFFCE_PN0P_  (.D(_01028_),
    .DE(_00088_),
    .Q(\w[23][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][28]$_SDFFCE_PN0P_  (.D(_01029_),
    .DE(_00088_),
    .Q(\w[23][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][29]$_SDFFCE_PN0P_  (.D(_01030_),
    .DE(_00088_),
    .Q(\w[23][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][2]$_SDFFCE_PN0P_  (.D(_01031_),
    .DE(_00088_),
    .Q(\w[23][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][30]$_SDFFCE_PN0P_  (.D(_01032_),
    .DE(_00088_),
    .Q(\w[23][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][31]$_SDFFCE_PN0P_  (.D(_01033_),
    .DE(_00088_),
    .Q(\w[23][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][3]$_SDFFCE_PN0P_  (.D(_01034_),
    .DE(_00088_),
    .Q(\w[23][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][4]$_SDFFCE_PN0P_  (.D(_01035_),
    .DE(_00088_),
    .Q(\w[23][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][5]$_SDFFCE_PN0P_  (.D(_01036_),
    .DE(_00088_),
    .Q(\w[23][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][6]$_SDFFCE_PN0P_  (.D(_01037_),
    .DE(_00088_),
    .Q(\w[23][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][7]$_SDFFCE_PN0P_  (.D(_01038_),
    .DE(_00088_),
    .Q(\w[23][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][8]$_SDFFCE_PN0P_  (.D(_01039_),
    .DE(_00088_),
    .Q(\w[23][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][9]$_SDFFCE_PN0P_  (.D(_01040_),
    .DE(_00088_),
    .Q(\w[23][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][0]$_SDFFCE_PN0P_  (.D(_01041_),
    .DE(_00119_),
    .Q(\w[24][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][10]$_SDFFCE_PN0P_  (.D(_01042_),
    .DE(_00119_),
    .Q(\w[24][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][11]$_SDFFCE_PN0P_  (.D(_01043_),
    .DE(_00119_),
    .Q(\w[24][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][12]$_SDFFCE_PN0P_  (.D(_01044_),
    .DE(_00119_),
    .Q(\w[24][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][13]$_SDFFCE_PN0P_  (.D(_01045_),
    .DE(_00119_),
    .Q(\w[24][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][14]$_SDFFCE_PN0P_  (.D(_01046_),
    .DE(_00119_),
    .Q(\w[24][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][15]$_SDFFCE_PN0P_  (.D(_01047_),
    .DE(_00119_),
    .Q(\w[24][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][16]$_SDFFCE_PN0P_  (.D(_01048_),
    .DE(_00119_),
    .Q(\w[24][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][17]$_SDFFCE_PN0P_  (.D(_01049_),
    .DE(_00119_),
    .Q(\w[24][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][18]$_SDFFCE_PN0P_  (.D(_01050_),
    .DE(_00119_),
    .Q(\w[24][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][19]$_SDFFCE_PN0P_  (.D(_01051_),
    .DE(_00119_),
    .Q(\w[24][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][1]$_SDFFCE_PN0P_  (.D(_01052_),
    .DE(_00119_),
    .Q(\w[24][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][20]$_SDFFCE_PN0P_  (.D(_01053_),
    .DE(_00119_),
    .Q(\w[24][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][21]$_SDFFCE_PN0P_  (.D(_01054_),
    .DE(_00119_),
    .Q(\w[24][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][22]$_SDFFCE_PN0P_  (.D(_01055_),
    .DE(_00119_),
    .Q(\w[24][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][23]$_SDFFCE_PN0P_  (.D(_01056_),
    .DE(_00119_),
    .Q(\w[24][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][24]$_SDFFCE_PN0P_  (.D(_01057_),
    .DE(_00119_),
    .Q(\w[24][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][25]$_SDFFCE_PN0P_  (.D(_01058_),
    .DE(_00119_),
    .Q(\w[24][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][26]$_SDFFCE_PN0P_  (.D(_01059_),
    .DE(_00119_),
    .Q(\w[24][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][27]$_SDFFCE_PN0P_  (.D(_01060_),
    .DE(_00119_),
    .Q(\w[24][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][28]$_SDFFCE_PN0P_  (.D(_01061_),
    .DE(_00119_),
    .Q(\w[24][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][29]$_SDFFCE_PN0P_  (.D(_01062_),
    .DE(_00119_),
    .Q(\w[24][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][2]$_SDFFCE_PN0P_  (.D(_01063_),
    .DE(_00119_),
    .Q(\w[24][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][30]$_SDFFCE_PN0P_  (.D(_01064_),
    .DE(_00119_),
    .Q(\w[24][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][31]$_SDFFCE_PN0P_  (.D(_01065_),
    .DE(_00119_),
    .Q(\w[24][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][3]$_SDFFCE_PN0P_  (.D(_01066_),
    .DE(_00119_),
    .Q(\w[24][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][4]$_SDFFCE_PN0P_  (.D(_01067_),
    .DE(_00119_),
    .Q(\w[24][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][5]$_SDFFCE_PN0P_  (.D(_01068_),
    .DE(_00119_),
    .Q(\w[24][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][6]$_SDFFCE_PN0P_  (.D(_01069_),
    .DE(_00119_),
    .Q(\w[24][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][7]$_SDFFCE_PN0P_  (.D(_01070_),
    .DE(_00119_),
    .Q(\w[24][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][8]$_SDFFCE_PN0P_  (.D(_01071_),
    .DE(_00119_),
    .Q(\w[24][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][9]$_SDFFCE_PN0P_  (.D(_01072_),
    .DE(_00119_),
    .Q(\w[24][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][0]$_SDFFCE_PN0P_  (.D(_01073_),
    .DE(_00087_),
    .Q(\w[25][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][10]$_SDFFCE_PN0P_  (.D(_01074_),
    .DE(_00087_),
    .Q(\w[25][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][11]$_SDFFCE_PN0P_  (.D(_01075_),
    .DE(_00087_),
    .Q(\w[25][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][12]$_SDFFCE_PN0P_  (.D(_01076_),
    .DE(_00087_),
    .Q(\w[25][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][13]$_SDFFCE_PN0P_  (.D(_01077_),
    .DE(_00087_),
    .Q(\w[25][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][14]$_SDFFCE_PN0P_  (.D(_01078_),
    .DE(_00087_),
    .Q(\w[25][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][15]$_SDFFCE_PN0P_  (.D(_01079_),
    .DE(_00087_),
    .Q(\w[25][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][16]$_SDFFCE_PN0P_  (.D(_01080_),
    .DE(_00087_),
    .Q(\w[25][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][17]$_SDFFCE_PN0P_  (.D(_01081_),
    .DE(_00087_),
    .Q(\w[25][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][18]$_SDFFCE_PN0P_  (.D(_01082_),
    .DE(_00087_),
    .Q(\w[25][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][19]$_SDFFCE_PN0P_  (.D(_01083_),
    .DE(_00087_),
    .Q(\w[25][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][1]$_SDFFCE_PN0P_  (.D(_01084_),
    .DE(_00087_),
    .Q(\w[25][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][20]$_SDFFCE_PN0P_  (.D(_01085_),
    .DE(_00087_),
    .Q(\w[25][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][21]$_SDFFCE_PN0P_  (.D(_01086_),
    .DE(_00087_),
    .Q(\w[25][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][22]$_SDFFCE_PN0P_  (.D(_01087_),
    .DE(_00087_),
    .Q(\w[25][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][23]$_SDFFCE_PN0P_  (.D(_01088_),
    .DE(_00087_),
    .Q(\w[25][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][24]$_SDFFCE_PN0P_  (.D(_01089_),
    .DE(_00087_),
    .Q(\w[25][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][25]$_SDFFCE_PN0P_  (.D(_01090_),
    .DE(_00087_),
    .Q(\w[25][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][26]$_SDFFCE_PN0P_  (.D(_01091_),
    .DE(_00087_),
    .Q(\w[25][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][27]$_SDFFCE_PN0P_  (.D(_01092_),
    .DE(_00087_),
    .Q(\w[25][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][28]$_SDFFCE_PN0P_  (.D(_01093_),
    .DE(_00087_),
    .Q(\w[25][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][29]$_SDFFCE_PN0P_  (.D(_01094_),
    .DE(_00087_),
    .Q(\w[25][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][2]$_SDFFCE_PN0P_  (.D(_01095_),
    .DE(_00087_),
    .Q(\w[25][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][30]$_SDFFCE_PN0P_  (.D(_01096_),
    .DE(_00087_),
    .Q(\w[25][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][31]$_SDFFCE_PN0P_  (.D(_01097_),
    .DE(_00087_),
    .Q(\w[25][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][3]$_SDFFCE_PN0P_  (.D(_01098_),
    .DE(_00087_),
    .Q(\w[25][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][4]$_SDFFCE_PN0P_  (.D(_01099_),
    .DE(_00087_),
    .Q(\w[25][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][5]$_SDFFCE_PN0P_  (.D(_01100_),
    .DE(_00087_),
    .Q(\w[25][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][6]$_SDFFCE_PN0P_  (.D(_01101_),
    .DE(_00087_),
    .Q(\w[25][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][7]$_SDFFCE_PN0P_  (.D(_01102_),
    .DE(_00087_),
    .Q(\w[25][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][8]$_SDFFCE_PN0P_  (.D(_01103_),
    .DE(_00087_),
    .Q(\w[25][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][9]$_SDFFCE_PN0P_  (.D(_01104_),
    .DE(_00087_),
    .Q(\w[25][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][0]$_SDFFCE_PN0P_  (.D(_01105_),
    .DE(_00118_),
    .Q(\w[26][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][10]$_SDFFCE_PN0P_  (.D(_01106_),
    .DE(_00118_),
    .Q(\w[26][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][11]$_SDFFCE_PN0P_  (.D(_01107_),
    .DE(_00118_),
    .Q(\w[26][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][12]$_SDFFCE_PN0P_  (.D(_01108_),
    .DE(_00118_),
    .Q(\w[26][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][13]$_SDFFCE_PN0P_  (.D(_01109_),
    .DE(_00118_),
    .Q(\w[26][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][14]$_SDFFCE_PN0P_  (.D(_01110_),
    .DE(_00118_),
    .Q(\w[26][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][15]$_SDFFCE_PN0P_  (.D(_01111_),
    .DE(_00118_),
    .Q(\w[26][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][16]$_SDFFCE_PN0P_  (.D(_01112_),
    .DE(_00118_),
    .Q(\w[26][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][17]$_SDFFCE_PN0P_  (.D(_01113_),
    .DE(_00118_),
    .Q(\w[26][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][18]$_SDFFCE_PN0P_  (.D(_01114_),
    .DE(_00118_),
    .Q(\w[26][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][19]$_SDFFCE_PN0P_  (.D(_01115_),
    .DE(_00118_),
    .Q(\w[26][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][1]$_SDFFCE_PN0P_  (.D(_01116_),
    .DE(_00118_),
    .Q(\w[26][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][20]$_SDFFCE_PN0P_  (.D(_01117_),
    .DE(_00118_),
    .Q(\w[26][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][21]$_SDFFCE_PN0P_  (.D(_01118_),
    .DE(_00118_),
    .Q(\w[26][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][22]$_SDFFCE_PN0P_  (.D(_01119_),
    .DE(_00118_),
    .Q(\w[26][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][23]$_SDFFCE_PN0P_  (.D(_01120_),
    .DE(_00118_),
    .Q(\w[26][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][24]$_SDFFCE_PN0P_  (.D(_01121_),
    .DE(_00118_),
    .Q(\w[26][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][25]$_SDFFCE_PN0P_  (.D(_01122_),
    .DE(_00118_),
    .Q(\w[26][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][26]$_SDFFCE_PN0P_  (.D(_01123_),
    .DE(_00118_),
    .Q(\w[26][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][27]$_SDFFCE_PN0P_  (.D(_01124_),
    .DE(_00118_),
    .Q(\w[26][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][28]$_SDFFCE_PN0P_  (.D(_01125_),
    .DE(_00118_),
    .Q(\w[26][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][29]$_SDFFCE_PN0P_  (.D(_01126_),
    .DE(_00118_),
    .Q(\w[26][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][2]$_SDFFCE_PN0P_  (.D(_01127_),
    .DE(_00118_),
    .Q(\w[26][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][30]$_SDFFCE_PN0P_  (.D(_01128_),
    .DE(_00118_),
    .Q(\w[26][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][31]$_SDFFCE_PN0P_  (.D(_01129_),
    .DE(_00118_),
    .Q(\w[26][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][3]$_SDFFCE_PN0P_  (.D(_01130_),
    .DE(_00118_),
    .Q(\w[26][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][4]$_SDFFCE_PN0P_  (.D(_01131_),
    .DE(_00118_),
    .Q(\w[26][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][5]$_SDFFCE_PN0P_  (.D(_01132_),
    .DE(_00118_),
    .Q(\w[26][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][6]$_SDFFCE_PN0P_  (.D(_01133_),
    .DE(_00118_),
    .Q(\w[26][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][7]$_SDFFCE_PN0P_  (.D(_01134_),
    .DE(_00118_),
    .Q(\w[26][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][8]$_SDFFCE_PN0P_  (.D(_01135_),
    .DE(_00118_),
    .Q(\w[26][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][9]$_SDFFCE_PN0P_  (.D(_01136_),
    .DE(_00118_),
    .Q(\w[26][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][0]$_SDFFCE_PN0P_  (.D(_01137_),
    .DE(_00086_),
    .Q(\w[27][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][10]$_SDFFCE_PN0P_  (.D(_01138_),
    .DE(_00086_),
    .Q(\w[27][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][11]$_SDFFCE_PN0P_  (.D(_01139_),
    .DE(_00086_),
    .Q(\w[27][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][12]$_SDFFCE_PN0P_  (.D(_01140_),
    .DE(_00086_),
    .Q(\w[27][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][13]$_SDFFCE_PN0P_  (.D(_01141_),
    .DE(_00086_),
    .Q(\w[27][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][14]$_SDFFCE_PN0P_  (.D(_01142_),
    .DE(_00086_),
    .Q(\w[27][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][15]$_SDFFCE_PN0P_  (.D(_01143_),
    .DE(_00086_),
    .Q(\w[27][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][16]$_SDFFCE_PN0P_  (.D(_01144_),
    .DE(_00086_),
    .Q(\w[27][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][17]$_SDFFCE_PN0P_  (.D(_01145_),
    .DE(_00086_),
    .Q(\w[27][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][18]$_SDFFCE_PN0P_  (.D(_01146_),
    .DE(_00086_),
    .Q(\w[27][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][19]$_SDFFCE_PN0P_  (.D(_01147_),
    .DE(_00086_),
    .Q(\w[27][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][1]$_SDFFCE_PN0P_  (.D(_01148_),
    .DE(_00086_),
    .Q(\w[27][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][20]$_SDFFCE_PN0P_  (.D(_01149_),
    .DE(_00086_),
    .Q(\w[27][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][21]$_SDFFCE_PN0P_  (.D(_01150_),
    .DE(_00086_),
    .Q(\w[27][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][22]$_SDFFCE_PN0P_  (.D(_01151_),
    .DE(_00086_),
    .Q(\w[27][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][23]$_SDFFCE_PN0P_  (.D(_01152_),
    .DE(_00086_),
    .Q(\w[27][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][24]$_SDFFCE_PN0P_  (.D(_01153_),
    .DE(_00086_),
    .Q(\w[27][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][25]$_SDFFCE_PN0P_  (.D(_01154_),
    .DE(_00086_),
    .Q(\w[27][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][26]$_SDFFCE_PN0P_  (.D(_01155_),
    .DE(_00086_),
    .Q(\w[27][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][27]$_SDFFCE_PN0P_  (.D(_01156_),
    .DE(_00086_),
    .Q(\w[27][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][28]$_SDFFCE_PN0P_  (.D(_01157_),
    .DE(_00086_),
    .Q(\w[27][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][29]$_SDFFCE_PN0P_  (.D(_01158_),
    .DE(_00086_),
    .Q(\w[27][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][2]$_SDFFCE_PN0P_  (.D(_01159_),
    .DE(_00086_),
    .Q(\w[27][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][30]$_SDFFCE_PN0P_  (.D(_01160_),
    .DE(_00086_),
    .Q(\w[27][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][31]$_SDFFCE_PN0P_  (.D(_01161_),
    .DE(_00086_),
    .Q(\w[27][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][3]$_SDFFCE_PN0P_  (.D(_01162_),
    .DE(_00086_),
    .Q(\w[27][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][4]$_SDFFCE_PN0P_  (.D(_01163_),
    .DE(_00086_),
    .Q(\w[27][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][5]$_SDFFCE_PN0P_  (.D(_01164_),
    .DE(_00086_),
    .Q(\w[27][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][6]$_SDFFCE_PN0P_  (.D(_01165_),
    .DE(_00086_),
    .Q(\w[27][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][7]$_SDFFCE_PN0P_  (.D(_01166_),
    .DE(_00086_),
    .Q(\w[27][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][8]$_SDFFCE_PN0P_  (.D(_01167_),
    .DE(_00086_),
    .Q(\w[27][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][9]$_SDFFCE_PN0P_  (.D(_01168_),
    .DE(_00086_),
    .Q(\w[27][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][0]$_SDFFCE_PN0P_  (.D(_01169_),
    .DE(_00117_),
    .Q(\w[28][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][10]$_SDFFCE_PN0P_  (.D(_01170_),
    .DE(_00117_),
    .Q(\w[28][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][11]$_SDFFCE_PN0P_  (.D(_01171_),
    .DE(_00117_),
    .Q(\w[28][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][12]$_SDFFCE_PN0P_  (.D(_01172_),
    .DE(_00117_),
    .Q(\w[28][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][13]$_SDFFCE_PN0P_  (.D(_01173_),
    .DE(_00117_),
    .Q(\w[28][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][14]$_SDFFCE_PN0P_  (.D(_01174_),
    .DE(_00117_),
    .Q(\w[28][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][15]$_SDFFCE_PN0P_  (.D(_01175_),
    .DE(_00117_),
    .Q(\w[28][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][16]$_SDFFCE_PN0P_  (.D(_01176_),
    .DE(_00117_),
    .Q(\w[28][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][17]$_SDFFCE_PN0P_  (.D(_01177_),
    .DE(_00117_),
    .Q(\w[28][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][18]$_SDFFCE_PN0P_  (.D(_01178_),
    .DE(_00117_),
    .Q(\w[28][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][19]$_SDFFCE_PN0P_  (.D(_01179_),
    .DE(_00117_),
    .Q(\w[28][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][1]$_SDFFCE_PN0P_  (.D(_01180_),
    .DE(_00117_),
    .Q(\w[28][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][20]$_SDFFCE_PN0P_  (.D(_01181_),
    .DE(_00117_),
    .Q(\w[28][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][21]$_SDFFCE_PN0P_  (.D(_01182_),
    .DE(_00117_),
    .Q(\w[28][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][22]$_SDFFCE_PN0P_  (.D(_01183_),
    .DE(_00117_),
    .Q(\w[28][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][23]$_SDFFCE_PN0P_  (.D(_01184_),
    .DE(_00117_),
    .Q(\w[28][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][24]$_SDFFCE_PN0P_  (.D(_01185_),
    .DE(_00117_),
    .Q(\w[28][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][25]$_SDFFCE_PN0P_  (.D(_01186_),
    .DE(_00117_),
    .Q(\w[28][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][26]$_SDFFCE_PN0P_  (.D(_01187_),
    .DE(_00117_),
    .Q(\w[28][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][27]$_SDFFCE_PN0P_  (.D(_01188_),
    .DE(_00117_),
    .Q(\w[28][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][28]$_SDFFCE_PN0P_  (.D(_01189_),
    .DE(_00117_),
    .Q(\w[28][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][29]$_SDFFCE_PN0P_  (.D(_01190_),
    .DE(_00117_),
    .Q(\w[28][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][2]$_SDFFCE_PN0P_  (.D(_01191_),
    .DE(_00117_),
    .Q(\w[28][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][30]$_SDFFCE_PN0P_  (.D(_01192_),
    .DE(_00117_),
    .Q(\w[28][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][31]$_SDFFCE_PN0P_  (.D(_01193_),
    .DE(_00117_),
    .Q(\w[28][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][3]$_SDFFCE_PN0P_  (.D(_01194_),
    .DE(_00117_),
    .Q(\w[28][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][4]$_SDFFCE_PN0P_  (.D(_01195_),
    .DE(_00117_),
    .Q(\w[28][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][5]$_SDFFCE_PN0P_  (.D(_01196_),
    .DE(_00117_),
    .Q(\w[28][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][6]$_SDFFCE_PN0P_  (.D(_01197_),
    .DE(_00117_),
    .Q(\w[28][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][7]$_SDFFCE_PN0P_  (.D(_01198_),
    .DE(_00117_),
    .Q(\w[28][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][8]$_SDFFCE_PN0P_  (.D(_01199_),
    .DE(_00117_),
    .Q(\w[28][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][9]$_SDFFCE_PN0P_  (.D(_01200_),
    .DE(_00117_),
    .Q(\w[28][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][0]$_SDFFCE_PN0P_  (.D(_01201_),
    .DE(_00085_),
    .Q(\w[29][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][10]$_SDFFCE_PN0P_  (.D(_01202_),
    .DE(_00085_),
    .Q(\w[29][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][11]$_SDFFCE_PN0P_  (.D(_01203_),
    .DE(_00085_),
    .Q(\w[29][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][12]$_SDFFCE_PN0P_  (.D(_01204_),
    .DE(_00085_),
    .Q(\w[29][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][13]$_SDFFCE_PN0P_  (.D(_01205_),
    .DE(_00085_),
    .Q(\w[29][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][14]$_SDFFCE_PN0P_  (.D(_01206_),
    .DE(_00085_),
    .Q(\w[29][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][15]$_SDFFCE_PN0P_  (.D(_01207_),
    .DE(_00085_),
    .Q(\w[29][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][16]$_SDFFCE_PN0P_  (.D(_01208_),
    .DE(_00085_),
    .Q(\w[29][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][17]$_SDFFCE_PN0P_  (.D(_01209_),
    .DE(_00085_),
    .Q(\w[29][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][18]$_SDFFCE_PN0P_  (.D(_01210_),
    .DE(_00085_),
    .Q(\w[29][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][19]$_SDFFCE_PN0P_  (.D(_01211_),
    .DE(_00085_),
    .Q(\w[29][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][1]$_SDFFCE_PN0P_  (.D(_01212_),
    .DE(_00085_),
    .Q(\w[29][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][20]$_SDFFCE_PN0P_  (.D(_01213_),
    .DE(_00085_),
    .Q(\w[29][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][21]$_SDFFCE_PN0P_  (.D(_01214_),
    .DE(_00085_),
    .Q(\w[29][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][22]$_SDFFCE_PN0P_  (.D(_01215_),
    .DE(_00085_),
    .Q(\w[29][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][23]$_SDFFCE_PN0P_  (.D(_01216_),
    .DE(_00085_),
    .Q(\w[29][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][24]$_SDFFCE_PN0P_  (.D(_01217_),
    .DE(_00085_),
    .Q(\w[29][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][25]$_SDFFCE_PN0P_  (.D(_01218_),
    .DE(_00085_),
    .Q(\w[29][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][26]$_SDFFCE_PN0P_  (.D(_01219_),
    .DE(_00085_),
    .Q(\w[29][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][27]$_SDFFCE_PN0P_  (.D(_01220_),
    .DE(_00085_),
    .Q(\w[29][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][28]$_SDFFCE_PN0P_  (.D(_01221_),
    .DE(_00085_),
    .Q(\w[29][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][29]$_SDFFCE_PN0P_  (.D(_01222_),
    .DE(_00085_),
    .Q(\w[29][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][2]$_SDFFCE_PN0P_  (.D(_01223_),
    .DE(_00085_),
    .Q(\w[29][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][30]$_SDFFCE_PN0P_  (.D(_01224_),
    .DE(_00085_),
    .Q(\w[29][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][31]$_SDFFCE_PN0P_  (.D(_01225_),
    .DE(_00085_),
    .Q(\w[29][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][3]$_SDFFCE_PN0P_  (.D(_01226_),
    .DE(_00085_),
    .Q(\w[29][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][4]$_SDFFCE_PN0P_  (.D(_01227_),
    .DE(_00085_),
    .Q(\w[29][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][5]$_SDFFCE_PN0P_  (.D(_01228_),
    .DE(_00085_),
    .Q(\w[29][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][6]$_SDFFCE_PN0P_  (.D(_01229_),
    .DE(_00085_),
    .Q(\w[29][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][7]$_SDFFCE_PN0P_  (.D(_01230_),
    .DE(_00085_),
    .Q(\w[29][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][8]$_SDFFCE_PN0P_  (.D(_01231_),
    .DE(_00085_),
    .Q(\w[29][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][9]$_SDFFCE_PN0P_  (.D(_01232_),
    .DE(_00085_),
    .Q(\w[29][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][0]$_DFFE_PP_  (.D(_00385_),
    .DE(_00116_),
    .Q(\w[2][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][10]$_DFFE_PP_  (.D(_00386_),
    .DE(_00116_),
    .Q(\w[2][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][11]$_DFFE_PP_  (.D(_00387_),
    .DE(_00116_),
    .Q(\w[2][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][12]$_DFFE_PP_  (.D(_00388_),
    .DE(_00116_),
    .Q(\w[2][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][13]$_DFFE_PP_  (.D(_00389_),
    .DE(_00116_),
    .Q(\w[2][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][14]$_DFFE_PP_  (.D(_00390_),
    .DE(_00116_),
    .Q(\w[2][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][15]$_DFFE_PP_  (.D(_00391_),
    .DE(_00116_),
    .Q(\w[2][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][16]$_DFFE_PP_  (.D(_00392_),
    .DE(_00116_),
    .Q(\w[2][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][17]$_DFFE_PP_  (.D(_00393_),
    .DE(_00116_),
    .Q(\w[2][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][18]$_DFFE_PP_  (.D(_00394_),
    .DE(_00116_),
    .Q(\w[2][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][19]$_DFFE_PP_  (.D(_00395_),
    .DE(_00116_),
    .Q(\w[2][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][1]$_DFFE_PP_  (.D(_00396_),
    .DE(_00116_),
    .Q(\w[2][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][20]$_DFFE_PP_  (.D(_00397_),
    .DE(_00116_),
    .Q(\w[2][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][21]$_DFFE_PP_  (.D(_00398_),
    .DE(_00116_),
    .Q(\w[2][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][22]$_DFFE_PP_  (.D(_00399_),
    .DE(_00116_),
    .Q(\w[2][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][23]$_DFFE_PP_  (.D(_00400_),
    .DE(_00116_),
    .Q(\w[2][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][24]$_DFFE_PP_  (.D(_00401_),
    .DE(_00116_),
    .Q(\w[2][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][25]$_DFFE_PP_  (.D(_00402_),
    .DE(_00116_),
    .Q(\w[2][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][26]$_DFFE_PP_  (.D(_00403_),
    .DE(_00116_),
    .Q(\w[2][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][27]$_DFFE_PP_  (.D(_00404_),
    .DE(_00116_),
    .Q(\w[2][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][28]$_DFFE_PP_  (.D(_00405_),
    .DE(_00116_),
    .Q(\w[2][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][29]$_DFFE_PP_  (.D(_00406_),
    .DE(_00116_),
    .Q(\w[2][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][2]$_DFFE_PP_  (.D(_00407_),
    .DE(_00116_),
    .Q(\w[2][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][30]$_DFFE_PP_  (.D(_00408_),
    .DE(_00116_),
    .Q(\w[2][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][31]$_DFFE_PP_  (.D(_00409_),
    .DE(_00116_),
    .Q(\w[2][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][3]$_DFFE_PP_  (.D(_00410_),
    .DE(_00116_),
    .Q(\w[2][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][4]$_DFFE_PP_  (.D(_00411_),
    .DE(_00116_),
    .Q(\w[2][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][5]$_DFFE_PP_  (.D(_00412_),
    .DE(_00116_),
    .Q(\w[2][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][6]$_DFFE_PP_  (.D(_00413_),
    .DE(_00116_),
    .Q(\w[2][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][7]$_DFFE_PP_  (.D(_00414_),
    .DE(_00116_),
    .Q(\w[2][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][8]$_DFFE_PP_  (.D(_00415_),
    .DE(_00116_),
    .Q(\w[2][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][9]$_DFFE_PP_  (.D(_00416_),
    .DE(_00116_),
    .Q(\w[2][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][0]$_SDFFCE_PN0P_  (.D(_01233_),
    .DE(_00115_),
    .Q(\w[30][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][10]$_SDFFCE_PN0P_  (.D(_01234_),
    .DE(_00115_),
    .Q(\w[30][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][11]$_SDFFCE_PN0P_  (.D(_01235_),
    .DE(_00115_),
    .Q(\w[30][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][12]$_SDFFCE_PN0P_  (.D(_01236_),
    .DE(_00115_),
    .Q(\w[30][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][13]$_SDFFCE_PN0P_  (.D(_01237_),
    .DE(_00115_),
    .Q(\w[30][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][14]$_SDFFCE_PN0P_  (.D(_01238_),
    .DE(_00115_),
    .Q(\w[30][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][15]$_SDFFCE_PN0P_  (.D(_01239_),
    .DE(_00115_),
    .Q(\w[30][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][16]$_SDFFCE_PN0P_  (.D(_01240_),
    .DE(_00115_),
    .Q(\w[30][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][17]$_SDFFCE_PN0P_  (.D(_01241_),
    .DE(_00115_),
    .Q(\w[30][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][18]$_SDFFCE_PN0P_  (.D(_01242_),
    .DE(_00115_),
    .Q(\w[30][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][19]$_SDFFCE_PN0P_  (.D(_01243_),
    .DE(_00115_),
    .Q(\w[30][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][1]$_SDFFCE_PN0P_  (.D(_01244_),
    .DE(_00115_),
    .Q(\w[30][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][20]$_SDFFCE_PN0P_  (.D(_01245_),
    .DE(_00115_),
    .Q(\w[30][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][21]$_SDFFCE_PN0P_  (.D(_01246_),
    .DE(_00115_),
    .Q(\w[30][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][22]$_SDFFCE_PN0P_  (.D(_01247_),
    .DE(_00115_),
    .Q(\w[30][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][23]$_SDFFCE_PN0P_  (.D(_01248_),
    .DE(_00115_),
    .Q(\w[30][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][24]$_SDFFCE_PN0P_  (.D(_01249_),
    .DE(_00115_),
    .Q(\w[30][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][25]$_SDFFCE_PN0P_  (.D(_01250_),
    .DE(_00115_),
    .Q(\w[30][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][26]$_SDFFCE_PN0P_  (.D(_01251_),
    .DE(_00115_),
    .Q(\w[30][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][27]$_SDFFCE_PN0P_  (.D(_01252_),
    .DE(_00115_),
    .Q(\w[30][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][28]$_SDFFCE_PN0P_  (.D(_01253_),
    .DE(_00115_),
    .Q(\w[30][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][29]$_SDFFCE_PN0P_  (.D(_01254_),
    .DE(_00115_),
    .Q(\w[30][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][2]$_SDFFCE_PN0P_  (.D(_01255_),
    .DE(_00115_),
    .Q(\w[30][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][30]$_SDFFCE_PN0P_  (.D(_01256_),
    .DE(_00115_),
    .Q(\w[30][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][31]$_SDFFCE_PN0P_  (.D(_01257_),
    .DE(_00115_),
    .Q(\w[30][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][3]$_SDFFCE_PN0P_  (.D(_01258_),
    .DE(_00115_),
    .Q(\w[30][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][4]$_SDFFCE_PN0P_  (.D(_01259_),
    .DE(_00115_),
    .Q(\w[30][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][5]$_SDFFCE_PN0P_  (.D(_01260_),
    .DE(_00115_),
    .Q(\w[30][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][6]$_SDFFCE_PN0P_  (.D(_01261_),
    .DE(_00115_),
    .Q(\w[30][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][7]$_SDFFCE_PN0P_  (.D(_01262_),
    .DE(_00115_),
    .Q(\w[30][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][8]$_SDFFCE_PN0P_  (.D(_01263_),
    .DE(_00115_),
    .Q(\w[30][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][9]$_SDFFCE_PN0P_  (.D(_01264_),
    .DE(_00115_),
    .Q(\w[30][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][0]$_SDFFCE_PN0P_  (.D(_01265_),
    .DE(_00084_),
    .Q(\w[31][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][10]$_SDFFCE_PN0P_  (.D(_01266_),
    .DE(_00084_),
    .Q(\w[31][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][11]$_SDFFCE_PN0P_  (.D(_01267_),
    .DE(_00084_),
    .Q(\w[31][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][12]$_SDFFCE_PN0P_  (.D(_01268_),
    .DE(_00084_),
    .Q(\w[31][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][13]$_SDFFCE_PN0P_  (.D(_01269_),
    .DE(_00084_),
    .Q(\w[31][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][14]$_SDFFCE_PN0P_  (.D(_01270_),
    .DE(_00084_),
    .Q(\w[31][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][15]$_SDFFCE_PN0P_  (.D(_01271_),
    .DE(_00084_),
    .Q(\w[31][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][16]$_SDFFCE_PN0P_  (.D(_01272_),
    .DE(_00084_),
    .Q(\w[31][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][17]$_SDFFCE_PN0P_  (.D(_01273_),
    .DE(_00084_),
    .Q(\w[31][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][18]$_SDFFCE_PN0P_  (.D(_01274_),
    .DE(_00084_),
    .Q(\w[31][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][19]$_SDFFCE_PN0P_  (.D(_01275_),
    .DE(_00084_),
    .Q(\w[31][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][1]$_SDFFCE_PN0P_  (.D(_01276_),
    .DE(_00084_),
    .Q(\w[31][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][20]$_SDFFCE_PN0P_  (.D(_01277_),
    .DE(_00084_),
    .Q(\w[31][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][21]$_SDFFCE_PN0P_  (.D(_01278_),
    .DE(_00084_),
    .Q(\w[31][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][22]$_SDFFCE_PN0P_  (.D(_01279_),
    .DE(_00084_),
    .Q(\w[31][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][23]$_SDFFCE_PN0P_  (.D(_01280_),
    .DE(_00084_),
    .Q(\w[31][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][24]$_SDFFCE_PN0P_  (.D(_01281_),
    .DE(_00084_),
    .Q(\w[31][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][25]$_SDFFCE_PN0P_  (.D(_01282_),
    .DE(_00084_),
    .Q(\w[31][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][26]$_SDFFCE_PN0P_  (.D(_01283_),
    .DE(_00084_),
    .Q(\w[31][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][27]$_SDFFCE_PN0P_  (.D(_01284_),
    .DE(_00084_),
    .Q(\w[31][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][28]$_SDFFCE_PN0P_  (.D(_01285_),
    .DE(_00084_),
    .Q(\w[31][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][29]$_SDFFCE_PN0P_  (.D(_01286_),
    .DE(_00084_),
    .Q(\w[31][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][2]$_SDFFCE_PN0P_  (.D(_01287_),
    .DE(_00084_),
    .Q(\w[31][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][30]$_SDFFCE_PN0P_  (.D(_01288_),
    .DE(_00084_),
    .Q(\w[31][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][31]$_SDFFCE_PN0P_  (.D(_01289_),
    .DE(_00084_),
    .Q(\w[31][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][3]$_SDFFCE_PN0P_  (.D(_01290_),
    .DE(_00084_),
    .Q(\w[31][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][4]$_SDFFCE_PN0P_  (.D(_01291_),
    .DE(_00084_),
    .Q(\w[31][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][5]$_SDFFCE_PN0P_  (.D(_01292_),
    .DE(_00084_),
    .Q(\w[31][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][6]$_SDFFCE_PN0P_  (.D(_01293_),
    .DE(_00084_),
    .Q(\w[31][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][7]$_SDFFCE_PN0P_  (.D(_01294_),
    .DE(_00084_),
    .Q(\w[31][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][8]$_SDFFCE_PN0P_  (.D(_01295_),
    .DE(_00084_),
    .Q(\w[31][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][9]$_SDFFCE_PN0P_  (.D(_01296_),
    .DE(_00084_),
    .Q(\w[31][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][0]$_SDFFCE_PN0P_  (.D(_01297_),
    .DE(_00114_),
    .Q(\w[32][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][10]$_SDFFCE_PN0P_  (.D(_01298_),
    .DE(_00114_),
    .Q(\w[32][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][11]$_SDFFCE_PN0P_  (.D(_01299_),
    .DE(_00114_),
    .Q(\w[32][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][12]$_SDFFCE_PN0P_  (.D(_01300_),
    .DE(_00114_),
    .Q(\w[32][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][13]$_SDFFCE_PN0P_  (.D(_01301_),
    .DE(_00114_),
    .Q(\w[32][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][14]$_SDFFCE_PN0P_  (.D(_01302_),
    .DE(_00114_),
    .Q(\w[32][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][15]$_SDFFCE_PN0P_  (.D(_01303_),
    .DE(_00114_),
    .Q(\w[32][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][16]$_SDFFCE_PN0P_  (.D(_01304_),
    .DE(_00114_),
    .Q(\w[32][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][17]$_SDFFCE_PN0P_  (.D(_01305_),
    .DE(_00114_),
    .Q(\w[32][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][18]$_SDFFCE_PN0P_  (.D(_01306_),
    .DE(_00114_),
    .Q(\w[32][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][19]$_SDFFCE_PN0P_  (.D(_01307_),
    .DE(_00114_),
    .Q(\w[32][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][1]$_SDFFCE_PN0P_  (.D(_01308_),
    .DE(_00114_),
    .Q(\w[32][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][20]$_SDFFCE_PN0P_  (.D(_01309_),
    .DE(_00114_),
    .Q(\w[32][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][21]$_SDFFCE_PN0P_  (.D(_01310_),
    .DE(_00114_),
    .Q(\w[32][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][22]$_SDFFCE_PN0P_  (.D(_01311_),
    .DE(_00114_),
    .Q(\w[32][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][23]$_SDFFCE_PN0P_  (.D(_01312_),
    .DE(_00114_),
    .Q(\w[32][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][24]$_SDFFCE_PN0P_  (.D(_01313_),
    .DE(_00114_),
    .Q(\w[32][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][25]$_SDFFCE_PN0P_  (.D(_01314_),
    .DE(_00114_),
    .Q(\w[32][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][26]$_SDFFCE_PN0P_  (.D(_01315_),
    .DE(_00114_),
    .Q(\w[32][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][27]$_SDFFCE_PN0P_  (.D(_01316_),
    .DE(_00114_),
    .Q(\w[32][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][28]$_SDFFCE_PN0P_  (.D(_01317_),
    .DE(_00114_),
    .Q(\w[32][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][29]$_SDFFCE_PN0P_  (.D(_01318_),
    .DE(_00114_),
    .Q(\w[32][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][2]$_SDFFCE_PN0P_  (.D(_01319_),
    .DE(_00114_),
    .Q(\w[32][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][30]$_SDFFCE_PN0P_  (.D(_01320_),
    .DE(_00114_),
    .Q(\w[32][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][31]$_SDFFCE_PN0P_  (.D(_01321_),
    .DE(_00114_),
    .Q(\w[32][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][3]$_SDFFCE_PN0P_  (.D(_01322_),
    .DE(_00114_),
    .Q(\w[32][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][4]$_SDFFCE_PN0P_  (.D(_01323_),
    .DE(_00114_),
    .Q(\w[32][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][5]$_SDFFCE_PN0P_  (.D(_01324_),
    .DE(_00114_),
    .Q(\w[32][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][6]$_SDFFCE_PN0P_  (.D(_01325_),
    .DE(_00114_),
    .Q(\w[32][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][7]$_SDFFCE_PN0P_  (.D(_01326_),
    .DE(_00114_),
    .Q(\w[32][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][8]$_SDFFCE_PN0P_  (.D(_01327_),
    .DE(_00114_),
    .Q(\w[32][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][9]$_SDFFCE_PN0P_  (.D(_01328_),
    .DE(_00114_),
    .Q(\w[32][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][0]$_SDFFCE_PN0P_  (.D(_01329_),
    .DE(_00083_),
    .Q(\w[33][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][10]$_SDFFCE_PN0P_  (.D(_01330_),
    .DE(_00083_),
    .Q(\w[33][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][11]$_SDFFCE_PN0P_  (.D(_01331_),
    .DE(_00083_),
    .Q(\w[33][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][12]$_SDFFCE_PN0P_  (.D(_01332_),
    .DE(_00083_),
    .Q(\w[33][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][13]$_SDFFCE_PN0P_  (.D(_01333_),
    .DE(_00083_),
    .Q(\w[33][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][14]$_SDFFCE_PN0P_  (.D(_01334_),
    .DE(_00083_),
    .Q(\w[33][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][15]$_SDFFCE_PN0P_  (.D(_01335_),
    .DE(_00083_),
    .Q(\w[33][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][16]$_SDFFCE_PN0P_  (.D(_01336_),
    .DE(_00083_),
    .Q(\w[33][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][17]$_SDFFCE_PN0P_  (.D(_01337_),
    .DE(_00083_),
    .Q(\w[33][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][18]$_SDFFCE_PN0P_  (.D(_01338_),
    .DE(_00083_),
    .Q(\w[33][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][19]$_SDFFCE_PN0P_  (.D(_01339_),
    .DE(_00083_),
    .Q(\w[33][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][1]$_SDFFCE_PN0P_  (.D(_01340_),
    .DE(_00083_),
    .Q(\w[33][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][20]$_SDFFCE_PN0P_  (.D(_01341_),
    .DE(_00083_),
    .Q(\w[33][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][21]$_SDFFCE_PN0P_  (.D(_01342_),
    .DE(_00083_),
    .Q(\w[33][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][22]$_SDFFCE_PN0P_  (.D(_01343_),
    .DE(_00083_),
    .Q(\w[33][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][23]$_SDFFCE_PN0P_  (.D(_01344_),
    .DE(_00083_),
    .Q(\w[33][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][24]$_SDFFCE_PN0P_  (.D(_01345_),
    .DE(_00083_),
    .Q(\w[33][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][25]$_SDFFCE_PN0P_  (.D(_01346_),
    .DE(_00083_),
    .Q(\w[33][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][26]$_SDFFCE_PN0P_  (.D(_01347_),
    .DE(_00083_),
    .Q(\w[33][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][27]$_SDFFCE_PN0P_  (.D(_01348_),
    .DE(_00083_),
    .Q(\w[33][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][28]$_SDFFCE_PN0P_  (.D(_01349_),
    .DE(_00083_),
    .Q(\w[33][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][29]$_SDFFCE_PN0P_  (.D(_01350_),
    .DE(_00083_),
    .Q(\w[33][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][2]$_SDFFCE_PN0P_  (.D(_01351_),
    .DE(_00083_),
    .Q(\w[33][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][30]$_SDFFCE_PN0P_  (.D(_01352_),
    .DE(_00083_),
    .Q(\w[33][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][31]$_SDFFCE_PN0P_  (.D(_01353_),
    .DE(_00083_),
    .Q(\w[33][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][3]$_SDFFCE_PN0P_  (.D(_01354_),
    .DE(_00083_),
    .Q(\w[33][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][4]$_SDFFCE_PN0P_  (.D(_01355_),
    .DE(_00083_),
    .Q(\w[33][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][5]$_SDFFCE_PN0P_  (.D(_01356_),
    .DE(_00083_),
    .Q(\w[33][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][6]$_SDFFCE_PN0P_  (.D(_01357_),
    .DE(_00083_),
    .Q(\w[33][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][7]$_SDFFCE_PN0P_  (.D(_01358_),
    .DE(_00083_),
    .Q(\w[33][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][8]$_SDFFCE_PN0P_  (.D(_01359_),
    .DE(_00083_),
    .Q(\w[33][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][9]$_SDFFCE_PN0P_  (.D(_01360_),
    .DE(_00083_),
    .Q(\w[33][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][0]$_SDFFCE_PN0P_  (.D(_01361_),
    .DE(_00113_),
    .Q(\w[34][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][10]$_SDFFCE_PN0P_  (.D(_01362_),
    .DE(_00113_),
    .Q(\w[34][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][11]$_SDFFCE_PN0P_  (.D(_01363_),
    .DE(_00113_),
    .Q(\w[34][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][12]$_SDFFCE_PN0P_  (.D(_01364_),
    .DE(_00113_),
    .Q(\w[34][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][13]$_SDFFCE_PN0P_  (.D(_01365_),
    .DE(_00113_),
    .Q(\w[34][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][14]$_SDFFCE_PN0P_  (.D(_01366_),
    .DE(_00113_),
    .Q(\w[34][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][15]$_SDFFCE_PN0P_  (.D(_01367_),
    .DE(_00113_),
    .Q(\w[34][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][16]$_SDFFCE_PN0P_  (.D(_01368_),
    .DE(_00113_),
    .Q(\w[34][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][17]$_SDFFCE_PN0P_  (.D(_01369_),
    .DE(_00113_),
    .Q(\w[34][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][18]$_SDFFCE_PN0P_  (.D(_01370_),
    .DE(_00113_),
    .Q(\w[34][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][19]$_SDFFCE_PN0P_  (.D(_01371_),
    .DE(_00113_),
    .Q(\w[34][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][1]$_SDFFCE_PN0P_  (.D(_01372_),
    .DE(_00113_),
    .Q(\w[34][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][20]$_SDFFCE_PN0P_  (.D(_01373_),
    .DE(_00113_),
    .Q(\w[34][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][21]$_SDFFCE_PN0P_  (.D(_01374_),
    .DE(_00113_),
    .Q(\w[34][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][22]$_SDFFCE_PN0P_  (.D(_01375_),
    .DE(_00113_),
    .Q(\w[34][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][23]$_SDFFCE_PN0P_  (.D(_01376_),
    .DE(_00113_),
    .Q(\w[34][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][24]$_SDFFCE_PN0P_  (.D(_01377_),
    .DE(_00113_),
    .Q(\w[34][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][25]$_SDFFCE_PN0P_  (.D(_01378_),
    .DE(_00113_),
    .Q(\w[34][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][26]$_SDFFCE_PN0P_  (.D(_01379_),
    .DE(_00113_),
    .Q(\w[34][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][27]$_SDFFCE_PN0P_  (.D(_01380_),
    .DE(_00113_),
    .Q(\w[34][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][28]$_SDFFCE_PN0P_  (.D(_01381_),
    .DE(_00113_),
    .Q(\w[34][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][29]$_SDFFCE_PN0P_  (.D(_01382_),
    .DE(_00113_),
    .Q(\w[34][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][2]$_SDFFCE_PN0P_  (.D(_01383_),
    .DE(_00113_),
    .Q(\w[34][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][30]$_SDFFCE_PN0P_  (.D(_01384_),
    .DE(_00113_),
    .Q(\w[34][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][31]$_SDFFCE_PN0P_  (.D(_01385_),
    .DE(_00113_),
    .Q(\w[34][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][3]$_SDFFCE_PN0P_  (.D(_01386_),
    .DE(_00113_),
    .Q(\w[34][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][4]$_SDFFCE_PN0P_  (.D(_01387_),
    .DE(_00113_),
    .Q(\w[34][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][5]$_SDFFCE_PN0P_  (.D(_01388_),
    .DE(_00113_),
    .Q(\w[34][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][6]$_SDFFCE_PN0P_  (.D(_01389_),
    .DE(_00113_),
    .Q(\w[34][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][7]$_SDFFCE_PN0P_  (.D(_01390_),
    .DE(_00113_),
    .Q(\w[34][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][8]$_SDFFCE_PN0P_  (.D(_01391_),
    .DE(_00113_),
    .Q(\w[34][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][9]$_SDFFCE_PN0P_  (.D(_01392_),
    .DE(_00113_),
    .Q(\w[34][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][0]$_SDFFCE_PN0P_  (.D(_01393_),
    .DE(_00082_),
    .Q(\w[35][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][10]$_SDFFCE_PN0P_  (.D(_01394_),
    .DE(_00082_),
    .Q(\w[35][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][11]$_SDFFCE_PN0P_  (.D(_01395_),
    .DE(_00082_),
    .Q(\w[35][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][12]$_SDFFCE_PN0P_  (.D(_01396_),
    .DE(_00082_),
    .Q(\w[35][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][13]$_SDFFCE_PN0P_  (.D(_01397_),
    .DE(_00082_),
    .Q(\w[35][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][14]$_SDFFCE_PN0P_  (.D(_01398_),
    .DE(_00082_),
    .Q(\w[35][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][15]$_SDFFCE_PN0P_  (.D(_01399_),
    .DE(_00082_),
    .Q(\w[35][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][16]$_SDFFCE_PN0P_  (.D(_01400_),
    .DE(_00082_),
    .Q(\w[35][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][17]$_SDFFCE_PN0P_  (.D(_01401_),
    .DE(_00082_),
    .Q(\w[35][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][18]$_SDFFCE_PN0P_  (.D(_01402_),
    .DE(_00082_),
    .Q(\w[35][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][19]$_SDFFCE_PN0P_  (.D(_01403_),
    .DE(_00082_),
    .Q(\w[35][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][1]$_SDFFCE_PN0P_  (.D(_01404_),
    .DE(_00082_),
    .Q(\w[35][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][20]$_SDFFCE_PN0P_  (.D(_01405_),
    .DE(_00082_),
    .Q(\w[35][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][21]$_SDFFCE_PN0P_  (.D(_01406_),
    .DE(_00082_),
    .Q(\w[35][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][22]$_SDFFCE_PN0P_  (.D(_01407_),
    .DE(_00082_),
    .Q(\w[35][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][23]$_SDFFCE_PN0P_  (.D(_01408_),
    .DE(_00082_),
    .Q(\w[35][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][24]$_SDFFCE_PN0P_  (.D(_01409_),
    .DE(_00082_),
    .Q(\w[35][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][25]$_SDFFCE_PN0P_  (.D(_01410_),
    .DE(_00082_),
    .Q(\w[35][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][26]$_SDFFCE_PN0P_  (.D(_01411_),
    .DE(_00082_),
    .Q(\w[35][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][27]$_SDFFCE_PN0P_  (.D(_01412_),
    .DE(_00082_),
    .Q(\w[35][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][28]$_SDFFCE_PN0P_  (.D(_01413_),
    .DE(_00082_),
    .Q(\w[35][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][29]$_SDFFCE_PN0P_  (.D(_01414_),
    .DE(_00082_),
    .Q(\w[35][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][2]$_SDFFCE_PN0P_  (.D(_01415_),
    .DE(_00082_),
    .Q(\w[35][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][30]$_SDFFCE_PN0P_  (.D(_01416_),
    .DE(_00082_),
    .Q(\w[35][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][31]$_SDFFCE_PN0P_  (.D(_01417_),
    .DE(_00082_),
    .Q(\w[35][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][3]$_SDFFCE_PN0P_  (.D(_01418_),
    .DE(_00082_),
    .Q(\w[35][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][4]$_SDFFCE_PN0P_  (.D(_01419_),
    .DE(_00082_),
    .Q(\w[35][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][5]$_SDFFCE_PN0P_  (.D(_01420_),
    .DE(_00082_),
    .Q(\w[35][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][6]$_SDFFCE_PN0P_  (.D(_01421_),
    .DE(_00082_),
    .Q(\w[35][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][7]$_SDFFCE_PN0P_  (.D(_01422_),
    .DE(_00082_),
    .Q(\w[35][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][8]$_SDFFCE_PN0P_  (.D(_01423_),
    .DE(_00082_),
    .Q(\w[35][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][9]$_SDFFCE_PN0P_  (.D(_01424_),
    .DE(_00082_),
    .Q(\w[35][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][0]$_SDFFCE_PN0P_  (.D(_01425_),
    .DE(_00112_),
    .Q(\w[36][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][10]$_SDFFCE_PN0P_  (.D(_01426_),
    .DE(_00112_),
    .Q(\w[36][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][11]$_SDFFCE_PN0P_  (.D(_01427_),
    .DE(_00112_),
    .Q(\w[36][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][12]$_SDFFCE_PN0P_  (.D(_01428_),
    .DE(_00112_),
    .Q(\w[36][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][13]$_SDFFCE_PN0P_  (.D(_01429_),
    .DE(_00112_),
    .Q(\w[36][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][14]$_SDFFCE_PN0P_  (.D(_01430_),
    .DE(_00112_),
    .Q(\w[36][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][15]$_SDFFCE_PN0P_  (.D(_01431_),
    .DE(_00112_),
    .Q(\w[36][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][16]$_SDFFCE_PN0P_  (.D(_01432_),
    .DE(_00112_),
    .Q(\w[36][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][17]$_SDFFCE_PN0P_  (.D(_01433_),
    .DE(_00112_),
    .Q(\w[36][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][18]$_SDFFCE_PN0P_  (.D(_01434_),
    .DE(_00112_),
    .Q(\w[36][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][19]$_SDFFCE_PN0P_  (.D(_01435_),
    .DE(_00112_),
    .Q(\w[36][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][1]$_SDFFCE_PN0P_  (.D(_01436_),
    .DE(_00112_),
    .Q(\w[36][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][20]$_SDFFCE_PN0P_  (.D(_01437_),
    .DE(_00112_),
    .Q(\w[36][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][21]$_SDFFCE_PN0P_  (.D(_01438_),
    .DE(_00112_),
    .Q(\w[36][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][22]$_SDFFCE_PN0P_  (.D(_01439_),
    .DE(_00112_),
    .Q(\w[36][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][23]$_SDFFCE_PN0P_  (.D(_01440_),
    .DE(_00112_),
    .Q(\w[36][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][24]$_SDFFCE_PN0P_  (.D(_01441_),
    .DE(_00112_),
    .Q(\w[36][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][25]$_SDFFCE_PN0P_  (.D(_01442_),
    .DE(_00112_),
    .Q(\w[36][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][26]$_SDFFCE_PN0P_  (.D(_01443_),
    .DE(_00112_),
    .Q(\w[36][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][27]$_SDFFCE_PN0P_  (.D(_01444_),
    .DE(_00112_),
    .Q(\w[36][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][28]$_SDFFCE_PN0P_  (.D(_01445_),
    .DE(_00112_),
    .Q(\w[36][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][29]$_SDFFCE_PN0P_  (.D(_01446_),
    .DE(_00112_),
    .Q(\w[36][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][2]$_SDFFCE_PN0P_  (.D(_01447_),
    .DE(_00112_),
    .Q(\w[36][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][30]$_SDFFCE_PN0P_  (.D(_01448_),
    .DE(_00112_),
    .Q(\w[36][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][31]$_SDFFCE_PN0P_  (.D(_01449_),
    .DE(_00112_),
    .Q(\w[36][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][3]$_SDFFCE_PN0P_  (.D(_01450_),
    .DE(_00112_),
    .Q(\w[36][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][4]$_SDFFCE_PN0P_  (.D(_01451_),
    .DE(_00112_),
    .Q(\w[36][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][5]$_SDFFCE_PN0P_  (.D(_01452_),
    .DE(_00112_),
    .Q(\w[36][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][6]$_SDFFCE_PN0P_  (.D(_01453_),
    .DE(_00112_),
    .Q(\w[36][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][7]$_SDFFCE_PN0P_  (.D(_01454_),
    .DE(_00112_),
    .Q(\w[36][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][8]$_SDFFCE_PN0P_  (.D(_01455_),
    .DE(_00112_),
    .Q(\w[36][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][9]$_SDFFCE_PN0P_  (.D(_01456_),
    .DE(_00112_),
    .Q(\w[36][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][0]$_SDFFCE_PN0P_  (.D(_01457_),
    .DE(_00081_),
    .Q(\w[37][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][10]$_SDFFCE_PN0P_  (.D(_01458_),
    .DE(_00081_),
    .Q(\w[37][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][11]$_SDFFCE_PN0P_  (.D(_01459_),
    .DE(_00081_),
    .Q(\w[37][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][12]$_SDFFCE_PN0P_  (.D(_01460_),
    .DE(_00081_),
    .Q(\w[37][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][13]$_SDFFCE_PN0P_  (.D(_01461_),
    .DE(_00081_),
    .Q(\w[37][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][14]$_SDFFCE_PN0P_  (.D(_01462_),
    .DE(_00081_),
    .Q(\w[37][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][15]$_SDFFCE_PN0P_  (.D(_01463_),
    .DE(_00081_),
    .Q(\w[37][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][16]$_SDFFCE_PN0P_  (.D(_01464_),
    .DE(_00081_),
    .Q(\w[37][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][17]$_SDFFCE_PN0P_  (.D(_01465_),
    .DE(_00081_),
    .Q(\w[37][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][18]$_SDFFCE_PN0P_  (.D(_01466_),
    .DE(_00081_),
    .Q(\w[37][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][19]$_SDFFCE_PN0P_  (.D(_01467_),
    .DE(_00081_),
    .Q(\w[37][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][1]$_SDFFCE_PN0P_  (.D(_01468_),
    .DE(_00081_),
    .Q(\w[37][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][20]$_SDFFCE_PN0P_  (.D(_01469_),
    .DE(_00081_),
    .Q(\w[37][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][21]$_SDFFCE_PN0P_  (.D(_01470_),
    .DE(_00081_),
    .Q(\w[37][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][22]$_SDFFCE_PN0P_  (.D(_01471_),
    .DE(_00081_),
    .Q(\w[37][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][23]$_SDFFCE_PN0P_  (.D(_01472_),
    .DE(_00081_),
    .Q(\w[37][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][24]$_SDFFCE_PN0P_  (.D(_01473_),
    .DE(_00081_),
    .Q(\w[37][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][25]$_SDFFCE_PN0P_  (.D(_01474_),
    .DE(_00081_),
    .Q(\w[37][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][26]$_SDFFCE_PN0P_  (.D(_01475_),
    .DE(_00081_),
    .Q(\w[37][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][27]$_SDFFCE_PN0P_  (.D(_01476_),
    .DE(_00081_),
    .Q(\w[37][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][28]$_SDFFCE_PN0P_  (.D(_01477_),
    .DE(_00081_),
    .Q(\w[37][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][29]$_SDFFCE_PN0P_  (.D(_01478_),
    .DE(_00081_),
    .Q(\w[37][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][2]$_SDFFCE_PN0P_  (.D(_01479_),
    .DE(_00081_),
    .Q(\w[37][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][30]$_SDFFCE_PN0P_  (.D(_01480_),
    .DE(_00081_),
    .Q(\w[37][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][31]$_SDFFCE_PN0P_  (.D(_01481_),
    .DE(_00081_),
    .Q(\w[37][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][3]$_SDFFCE_PN0P_  (.D(_01482_),
    .DE(_00081_),
    .Q(\w[37][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][4]$_SDFFCE_PN0P_  (.D(_01483_),
    .DE(_00081_),
    .Q(\w[37][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][5]$_SDFFCE_PN0P_  (.D(_01484_),
    .DE(_00081_),
    .Q(\w[37][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][6]$_SDFFCE_PN0P_  (.D(_01485_),
    .DE(_00081_),
    .Q(\w[37][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][7]$_SDFFCE_PN0P_  (.D(_01486_),
    .DE(_00081_),
    .Q(\w[37][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][8]$_SDFFCE_PN0P_  (.D(_01487_),
    .DE(_00081_),
    .Q(\w[37][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][9]$_SDFFCE_PN0P_  (.D(_01488_),
    .DE(_00081_),
    .Q(\w[37][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][0]$_SDFFCE_PN0P_  (.D(_01489_),
    .DE(_00111_),
    .Q(\w[38][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][10]$_SDFFCE_PN0P_  (.D(_01490_),
    .DE(_00111_),
    .Q(\w[38][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][11]$_SDFFCE_PN0P_  (.D(_01491_),
    .DE(_00111_),
    .Q(\w[38][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][12]$_SDFFCE_PN0P_  (.D(_01492_),
    .DE(_00111_),
    .Q(\w[38][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][13]$_SDFFCE_PN0P_  (.D(_01493_),
    .DE(_00111_),
    .Q(\w[38][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][14]$_SDFFCE_PN0P_  (.D(_01494_),
    .DE(_00111_),
    .Q(\w[38][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][15]$_SDFFCE_PN0P_  (.D(_01495_),
    .DE(_00111_),
    .Q(\w[38][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][16]$_SDFFCE_PN0P_  (.D(_01496_),
    .DE(_00111_),
    .Q(\w[38][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][17]$_SDFFCE_PN0P_  (.D(_01497_),
    .DE(_00111_),
    .Q(\w[38][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][18]$_SDFFCE_PN0P_  (.D(_01498_),
    .DE(_00111_),
    .Q(\w[38][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][19]$_SDFFCE_PN0P_  (.D(_01499_),
    .DE(_00111_),
    .Q(\w[38][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][1]$_SDFFCE_PN0P_  (.D(_01500_),
    .DE(_00111_),
    .Q(\w[38][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][20]$_SDFFCE_PN0P_  (.D(_01501_),
    .DE(_00111_),
    .Q(\w[38][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][21]$_SDFFCE_PN0P_  (.D(_01502_),
    .DE(_00111_),
    .Q(\w[38][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][22]$_SDFFCE_PN0P_  (.D(_01503_),
    .DE(_00111_),
    .Q(\w[38][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][23]$_SDFFCE_PN0P_  (.D(_01504_),
    .DE(_00111_),
    .Q(\w[38][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][24]$_SDFFCE_PN0P_  (.D(_01505_),
    .DE(_00111_),
    .Q(\w[38][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][25]$_SDFFCE_PN0P_  (.D(_01506_),
    .DE(_00111_),
    .Q(\w[38][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][26]$_SDFFCE_PN0P_  (.D(_01507_),
    .DE(_00111_),
    .Q(\w[38][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][27]$_SDFFCE_PN0P_  (.D(_01508_),
    .DE(_00111_),
    .Q(\w[38][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][28]$_SDFFCE_PN0P_  (.D(_01509_),
    .DE(_00111_),
    .Q(\w[38][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][29]$_SDFFCE_PN0P_  (.D(_01510_),
    .DE(_00111_),
    .Q(\w[38][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][2]$_SDFFCE_PN0P_  (.D(_01511_),
    .DE(_00111_),
    .Q(\w[38][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][30]$_SDFFCE_PN0P_  (.D(_01512_),
    .DE(_00111_),
    .Q(\w[38][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][31]$_SDFFCE_PN0P_  (.D(_01513_),
    .DE(_00111_),
    .Q(\w[38][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][3]$_SDFFCE_PN0P_  (.D(_01514_),
    .DE(_00111_),
    .Q(\w[38][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][4]$_SDFFCE_PN0P_  (.D(_01515_),
    .DE(_00111_),
    .Q(\w[38][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][5]$_SDFFCE_PN0P_  (.D(_01516_),
    .DE(_00111_),
    .Q(\w[38][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][6]$_SDFFCE_PN0P_  (.D(_01517_),
    .DE(_00111_),
    .Q(\w[38][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][7]$_SDFFCE_PN0P_  (.D(_01518_),
    .DE(_00111_),
    .Q(\w[38][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][8]$_SDFFCE_PN0P_  (.D(_01519_),
    .DE(_00111_),
    .Q(\w[38][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][9]$_SDFFCE_PN0P_  (.D(_01520_),
    .DE(_00111_),
    .Q(\w[38][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][0]$_SDFFCE_PN0P_  (.D(_01521_),
    .DE(_00080_),
    .Q(\w[39][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][10]$_SDFFCE_PN0P_  (.D(_01522_),
    .DE(_00080_),
    .Q(\w[39][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][11]$_SDFFCE_PN0P_  (.D(_01523_),
    .DE(_00080_),
    .Q(\w[39][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][12]$_SDFFCE_PN0P_  (.D(_01524_),
    .DE(_00080_),
    .Q(\w[39][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][13]$_SDFFCE_PN0P_  (.D(_01525_),
    .DE(_00080_),
    .Q(\w[39][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][14]$_SDFFCE_PN0P_  (.D(_01526_),
    .DE(_00080_),
    .Q(\w[39][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][15]$_SDFFCE_PN0P_  (.D(_01527_),
    .DE(_00080_),
    .Q(\w[39][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][16]$_SDFFCE_PN0P_  (.D(_01528_),
    .DE(_00080_),
    .Q(\w[39][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][17]$_SDFFCE_PN0P_  (.D(_01529_),
    .DE(_00080_),
    .Q(\w[39][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][18]$_SDFFCE_PN0P_  (.D(_01530_),
    .DE(_00080_),
    .Q(\w[39][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][19]$_SDFFCE_PN0P_  (.D(_01531_),
    .DE(_00080_),
    .Q(\w[39][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][1]$_SDFFCE_PN0P_  (.D(_01532_),
    .DE(_00080_),
    .Q(\w[39][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][20]$_SDFFCE_PN0P_  (.D(_01533_),
    .DE(_00080_),
    .Q(\w[39][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][21]$_SDFFCE_PN0P_  (.D(_01534_),
    .DE(_00080_),
    .Q(\w[39][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][22]$_SDFFCE_PN0P_  (.D(_01535_),
    .DE(_00080_),
    .Q(\w[39][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][23]$_SDFFCE_PN0P_  (.D(_01536_),
    .DE(_00080_),
    .Q(\w[39][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][24]$_SDFFCE_PN0P_  (.D(_01537_),
    .DE(_00080_),
    .Q(\w[39][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][25]$_SDFFCE_PN0P_  (.D(_01538_),
    .DE(_00080_),
    .Q(\w[39][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][26]$_SDFFCE_PN0P_  (.D(_01539_),
    .DE(_00080_),
    .Q(\w[39][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][27]$_SDFFCE_PN0P_  (.D(_01540_),
    .DE(_00080_),
    .Q(\w[39][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][28]$_SDFFCE_PN0P_  (.D(_01541_),
    .DE(_00080_),
    .Q(\w[39][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][29]$_SDFFCE_PN0P_  (.D(_01542_),
    .DE(_00080_),
    .Q(\w[39][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][2]$_SDFFCE_PN0P_  (.D(_01543_),
    .DE(_00080_),
    .Q(\w[39][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][30]$_SDFFCE_PN0P_  (.D(_01544_),
    .DE(_00080_),
    .Q(\w[39][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][31]$_SDFFCE_PN0P_  (.D(_01545_),
    .DE(_00080_),
    .Q(\w[39][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][3]$_SDFFCE_PN0P_  (.D(_01546_),
    .DE(_00080_),
    .Q(\w[39][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][4]$_SDFFCE_PN0P_  (.D(_01547_),
    .DE(_00080_),
    .Q(\w[39][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][5]$_SDFFCE_PN0P_  (.D(_01548_),
    .DE(_00080_),
    .Q(\w[39][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][6]$_SDFFCE_PN0P_  (.D(_01549_),
    .DE(_00080_),
    .Q(\w[39][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][7]$_SDFFCE_PN0P_  (.D(_01550_),
    .DE(_00080_),
    .Q(\w[39][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][8]$_SDFFCE_PN0P_  (.D(_01551_),
    .DE(_00080_),
    .Q(\w[39][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][9]$_SDFFCE_PN0P_  (.D(_01552_),
    .DE(_00080_),
    .Q(\w[39][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][0]$_DFFE_PP_  (.D(_00417_),
    .DE(_00079_),
    .Q(\w[3][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][10]$_DFFE_PP_  (.D(_00418_),
    .DE(_00079_),
    .Q(\w[3][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][11]$_DFFE_PP_  (.D(_00419_),
    .DE(_00079_),
    .Q(\w[3][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][12]$_DFFE_PP_  (.D(_00420_),
    .DE(_00079_),
    .Q(\w[3][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][13]$_DFFE_PP_  (.D(_00421_),
    .DE(_00079_),
    .Q(\w[3][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][14]$_DFFE_PP_  (.D(_00422_),
    .DE(_00079_),
    .Q(\w[3][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][15]$_DFFE_PP_  (.D(_00423_),
    .DE(_00079_),
    .Q(\w[3][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][16]$_DFFE_PP_  (.D(_00424_),
    .DE(_00079_),
    .Q(\w[3][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][17]$_DFFE_PP_  (.D(_00425_),
    .DE(_00079_),
    .Q(\w[3][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][18]$_DFFE_PP_  (.D(_00426_),
    .DE(_00079_),
    .Q(\w[3][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][19]$_DFFE_PP_  (.D(_00427_),
    .DE(_00079_),
    .Q(\w[3][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][1]$_DFFE_PP_  (.D(_00428_),
    .DE(_00079_),
    .Q(\w[3][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][20]$_DFFE_PP_  (.D(_00429_),
    .DE(_00079_),
    .Q(\w[3][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][21]$_DFFE_PP_  (.D(_00430_),
    .DE(_00079_),
    .Q(\w[3][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][22]$_DFFE_PP_  (.D(_00431_),
    .DE(_00079_),
    .Q(\w[3][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][23]$_DFFE_PP_  (.D(_00432_),
    .DE(_00079_),
    .Q(\w[3][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][24]$_DFFE_PP_  (.D(_00433_),
    .DE(_00079_),
    .Q(\w[3][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][25]$_DFFE_PP_  (.D(_00434_),
    .DE(_00079_),
    .Q(\w[3][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][26]$_DFFE_PP_  (.D(_00435_),
    .DE(_00079_),
    .Q(\w[3][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][27]$_DFFE_PP_  (.D(_00436_),
    .DE(_00079_),
    .Q(\w[3][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][28]$_DFFE_PP_  (.D(_00437_),
    .DE(_00079_),
    .Q(\w[3][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][29]$_DFFE_PP_  (.D(_00438_),
    .DE(_00079_),
    .Q(\w[3][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][2]$_DFFE_PP_  (.D(_00439_),
    .DE(_00079_),
    .Q(\w[3][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][30]$_DFFE_PP_  (.D(_00440_),
    .DE(_00079_),
    .Q(\w[3][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][31]$_DFFE_PP_  (.D(_00441_),
    .DE(_00079_),
    .Q(\w[3][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][3]$_DFFE_PP_  (.D(_00442_),
    .DE(_00079_),
    .Q(\w[3][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][4]$_DFFE_PP_  (.D(_00443_),
    .DE(_00079_),
    .Q(\w[3][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][5]$_DFFE_PP_  (.D(_00444_),
    .DE(_00079_),
    .Q(\w[3][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][6]$_DFFE_PP_  (.D(_00445_),
    .DE(_00079_),
    .Q(\w[3][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][7]$_DFFE_PP_  (.D(_00446_),
    .DE(_00079_),
    .Q(\w[3][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][8]$_DFFE_PP_  (.D(_00447_),
    .DE(_00079_),
    .Q(\w[3][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][9]$_DFFE_PP_  (.D(_00448_),
    .DE(_00079_),
    .Q(\w[3][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][0]$_SDFFCE_PN0P_  (.D(_01553_),
    .DE(_00110_),
    .Q(\w[40][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][10]$_SDFFCE_PN0P_  (.D(_01554_),
    .DE(_00110_),
    .Q(\w[40][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][11]$_SDFFCE_PN0P_  (.D(_01555_),
    .DE(_00110_),
    .Q(\w[40][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][12]$_SDFFCE_PN0P_  (.D(_01556_),
    .DE(_00110_),
    .Q(\w[40][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][13]$_SDFFCE_PN0P_  (.D(_01557_),
    .DE(_00110_),
    .Q(\w[40][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][14]$_SDFFCE_PN0P_  (.D(_01558_),
    .DE(_00110_),
    .Q(\w[40][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][15]$_SDFFCE_PN0P_  (.D(_01559_),
    .DE(_00110_),
    .Q(\w[40][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][16]$_SDFFCE_PN0P_  (.D(_01560_),
    .DE(_00110_),
    .Q(\w[40][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][17]$_SDFFCE_PN0P_  (.D(_01561_),
    .DE(_00110_),
    .Q(\w[40][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][18]$_SDFFCE_PN0P_  (.D(_01562_),
    .DE(_00110_),
    .Q(\w[40][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][19]$_SDFFCE_PN0P_  (.D(_01563_),
    .DE(_00110_),
    .Q(\w[40][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][1]$_SDFFCE_PN0P_  (.D(_01564_),
    .DE(_00110_),
    .Q(\w[40][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][20]$_SDFFCE_PN0P_  (.D(_01565_),
    .DE(_00110_),
    .Q(\w[40][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][21]$_SDFFCE_PN0P_  (.D(_01566_),
    .DE(_00110_),
    .Q(\w[40][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][22]$_SDFFCE_PN0P_  (.D(_01567_),
    .DE(_00110_),
    .Q(\w[40][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][23]$_SDFFCE_PN0P_  (.D(_01568_),
    .DE(_00110_),
    .Q(\w[40][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][24]$_SDFFCE_PN0P_  (.D(_01569_),
    .DE(_00110_),
    .Q(\w[40][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][25]$_SDFFCE_PN0P_  (.D(_01570_),
    .DE(_00110_),
    .Q(\w[40][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][26]$_SDFFCE_PN0P_  (.D(_01571_),
    .DE(_00110_),
    .Q(\w[40][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][27]$_SDFFCE_PN0P_  (.D(_01572_),
    .DE(_00110_),
    .Q(\w[40][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][28]$_SDFFCE_PN0P_  (.D(_01573_),
    .DE(_00110_),
    .Q(\w[40][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][29]$_SDFFCE_PN0P_  (.D(_01574_),
    .DE(_00110_),
    .Q(\w[40][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][2]$_SDFFCE_PN0P_  (.D(_01575_),
    .DE(_00110_),
    .Q(\w[40][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][30]$_SDFFCE_PN0P_  (.D(_01576_),
    .DE(_00110_),
    .Q(\w[40][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][31]$_SDFFCE_PN0P_  (.D(_01577_),
    .DE(_00110_),
    .Q(\w[40][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][3]$_SDFFCE_PN0P_  (.D(_01578_),
    .DE(_00110_),
    .Q(\w[40][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][4]$_SDFFCE_PN0P_  (.D(_01579_),
    .DE(_00110_),
    .Q(\w[40][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][5]$_SDFFCE_PN0P_  (.D(_01580_),
    .DE(_00110_),
    .Q(\w[40][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][6]$_SDFFCE_PN0P_  (.D(_01581_),
    .DE(_00110_),
    .Q(\w[40][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][7]$_SDFFCE_PN0P_  (.D(_01582_),
    .DE(_00110_),
    .Q(\w[40][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][8]$_SDFFCE_PN0P_  (.D(_01583_),
    .DE(_00110_),
    .Q(\w[40][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][9]$_SDFFCE_PN0P_  (.D(_01584_),
    .DE(_00110_),
    .Q(\w[40][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][0]$_SDFFCE_PN0P_  (.D(_01585_),
    .DE(_00078_),
    .Q(\w[41][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][10]$_SDFFCE_PN0P_  (.D(_01586_),
    .DE(_00078_),
    .Q(\w[41][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][11]$_SDFFCE_PN0P_  (.D(_01587_),
    .DE(_00078_),
    .Q(\w[41][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][12]$_SDFFCE_PN0P_  (.D(_01588_),
    .DE(_00078_),
    .Q(\w[41][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][13]$_SDFFCE_PN0P_  (.D(_01589_),
    .DE(_00078_),
    .Q(\w[41][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][14]$_SDFFCE_PN0P_  (.D(_01590_),
    .DE(_00078_),
    .Q(\w[41][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][15]$_SDFFCE_PN0P_  (.D(_01591_),
    .DE(_00078_),
    .Q(\w[41][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][16]$_SDFFCE_PN0P_  (.D(_01592_),
    .DE(_00078_),
    .Q(\w[41][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][17]$_SDFFCE_PN0P_  (.D(_01593_),
    .DE(_00078_),
    .Q(\w[41][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][18]$_SDFFCE_PN0P_  (.D(_01594_),
    .DE(_00078_),
    .Q(\w[41][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][19]$_SDFFCE_PN0P_  (.D(_01595_),
    .DE(_00078_),
    .Q(\w[41][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][1]$_SDFFCE_PN0P_  (.D(_01596_),
    .DE(_00078_),
    .Q(\w[41][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][20]$_SDFFCE_PN0P_  (.D(_01597_),
    .DE(_00078_),
    .Q(\w[41][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][21]$_SDFFCE_PN0P_  (.D(_01598_),
    .DE(_00078_),
    .Q(\w[41][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][22]$_SDFFCE_PN0P_  (.D(_01599_),
    .DE(_00078_),
    .Q(\w[41][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][23]$_SDFFCE_PN0P_  (.D(_01600_),
    .DE(_00078_),
    .Q(\w[41][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][24]$_SDFFCE_PN0P_  (.D(_01601_),
    .DE(_00078_),
    .Q(\w[41][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][25]$_SDFFCE_PN0P_  (.D(_01602_),
    .DE(_00078_),
    .Q(\w[41][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][26]$_SDFFCE_PN0P_  (.D(_01603_),
    .DE(_00078_),
    .Q(\w[41][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][27]$_SDFFCE_PN0P_  (.D(_01604_),
    .DE(_00078_),
    .Q(\w[41][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][28]$_SDFFCE_PN0P_  (.D(_01605_),
    .DE(_00078_),
    .Q(\w[41][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][29]$_SDFFCE_PN0P_  (.D(_01606_),
    .DE(_00078_),
    .Q(\w[41][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][2]$_SDFFCE_PN0P_  (.D(_01607_),
    .DE(_00078_),
    .Q(\w[41][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][30]$_SDFFCE_PN0P_  (.D(_01608_),
    .DE(_00078_),
    .Q(\w[41][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][31]$_SDFFCE_PN0P_  (.D(_01609_),
    .DE(_00078_),
    .Q(\w[41][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][3]$_SDFFCE_PN0P_  (.D(_01610_),
    .DE(_00078_),
    .Q(\w[41][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][4]$_SDFFCE_PN0P_  (.D(_01611_),
    .DE(_00078_),
    .Q(\w[41][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][5]$_SDFFCE_PN0P_  (.D(_01612_),
    .DE(_00078_),
    .Q(\w[41][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][6]$_SDFFCE_PN0P_  (.D(_01613_),
    .DE(_00078_),
    .Q(\w[41][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][7]$_SDFFCE_PN0P_  (.D(_01614_),
    .DE(_00078_),
    .Q(\w[41][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][8]$_SDFFCE_PN0P_  (.D(_01615_),
    .DE(_00078_),
    .Q(\w[41][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][9]$_SDFFCE_PN0P_  (.D(_01616_),
    .DE(_00078_),
    .Q(\w[41][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][0]$_SDFFCE_PN0P_  (.D(_01617_),
    .DE(_00109_),
    .Q(\w[42][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][10]$_SDFFCE_PN0P_  (.D(_01618_),
    .DE(_00109_),
    .Q(\w[42][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][11]$_SDFFCE_PN0P_  (.D(_01619_),
    .DE(_00109_),
    .Q(\w[42][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][12]$_SDFFCE_PN0P_  (.D(_01620_),
    .DE(_00109_),
    .Q(\w[42][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][13]$_SDFFCE_PN0P_  (.D(_01621_),
    .DE(_00109_),
    .Q(\w[42][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][14]$_SDFFCE_PN0P_  (.D(_01622_),
    .DE(_00109_),
    .Q(\w[42][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][15]$_SDFFCE_PN0P_  (.D(_01623_),
    .DE(_00109_),
    .Q(\w[42][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][16]$_SDFFCE_PN0P_  (.D(_01624_),
    .DE(_00109_),
    .Q(\w[42][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][17]$_SDFFCE_PN0P_  (.D(_01625_),
    .DE(_00109_),
    .Q(\w[42][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][18]$_SDFFCE_PN0P_  (.D(_01626_),
    .DE(_00109_),
    .Q(\w[42][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][19]$_SDFFCE_PN0P_  (.D(_01627_),
    .DE(_00109_),
    .Q(\w[42][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][1]$_SDFFCE_PN0P_  (.D(_01628_),
    .DE(_00109_),
    .Q(\w[42][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][20]$_SDFFCE_PN0P_  (.D(_01629_),
    .DE(_00109_),
    .Q(\w[42][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][21]$_SDFFCE_PN0P_  (.D(_01630_),
    .DE(_00109_),
    .Q(\w[42][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][22]$_SDFFCE_PN0P_  (.D(_01631_),
    .DE(_00109_),
    .Q(\w[42][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][23]$_SDFFCE_PN0P_  (.D(_01632_),
    .DE(_00109_),
    .Q(\w[42][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][24]$_SDFFCE_PN0P_  (.D(_01633_),
    .DE(_00109_),
    .Q(\w[42][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][25]$_SDFFCE_PN0P_  (.D(_01634_),
    .DE(_00109_),
    .Q(\w[42][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][26]$_SDFFCE_PN0P_  (.D(_01635_),
    .DE(_00109_),
    .Q(\w[42][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][27]$_SDFFCE_PN0P_  (.D(_01636_),
    .DE(_00109_),
    .Q(\w[42][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][28]$_SDFFCE_PN0P_  (.D(_01637_),
    .DE(_00109_),
    .Q(\w[42][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][29]$_SDFFCE_PN0P_  (.D(_01638_),
    .DE(_00109_),
    .Q(\w[42][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][2]$_SDFFCE_PN0P_  (.D(_01639_),
    .DE(_00109_),
    .Q(\w[42][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][30]$_SDFFCE_PN0P_  (.D(_01640_),
    .DE(_00109_),
    .Q(\w[42][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][31]$_SDFFCE_PN0P_  (.D(_01641_),
    .DE(_00109_),
    .Q(\w[42][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][3]$_SDFFCE_PN0P_  (.D(_01642_),
    .DE(_00109_),
    .Q(\w[42][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][4]$_SDFFCE_PN0P_  (.D(_01643_),
    .DE(_00109_),
    .Q(\w[42][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][5]$_SDFFCE_PN0P_  (.D(_01644_),
    .DE(_00109_),
    .Q(\w[42][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][6]$_SDFFCE_PN0P_  (.D(_01645_),
    .DE(_00109_),
    .Q(\w[42][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][7]$_SDFFCE_PN0P_  (.D(_01646_),
    .DE(_00109_),
    .Q(\w[42][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][8]$_SDFFCE_PN0P_  (.D(_01647_),
    .DE(_00109_),
    .Q(\w[42][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][9]$_SDFFCE_PN0P_  (.D(_01648_),
    .DE(_00109_),
    .Q(\w[42][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][0]$_SDFFCE_PN0P_  (.D(_01649_),
    .DE(_00077_),
    .Q(\w[43][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][10]$_SDFFCE_PN0P_  (.D(_01650_),
    .DE(_00077_),
    .Q(\w[43][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][11]$_SDFFCE_PN0P_  (.D(_01651_),
    .DE(_00077_),
    .Q(\w[43][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][12]$_SDFFCE_PN0P_  (.D(_01652_),
    .DE(_00077_),
    .Q(\w[43][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][13]$_SDFFCE_PN0P_  (.D(_01653_),
    .DE(_00077_),
    .Q(\w[43][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][14]$_SDFFCE_PN0P_  (.D(_01654_),
    .DE(_00077_),
    .Q(\w[43][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][15]$_SDFFCE_PN0P_  (.D(_01655_),
    .DE(_00077_),
    .Q(\w[43][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][16]$_SDFFCE_PN0P_  (.D(_01656_),
    .DE(_00077_),
    .Q(\w[43][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][17]$_SDFFCE_PN0P_  (.D(_01657_),
    .DE(_00077_),
    .Q(\w[43][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][18]$_SDFFCE_PN0P_  (.D(_01658_),
    .DE(_00077_),
    .Q(\w[43][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][19]$_SDFFCE_PN0P_  (.D(_01659_),
    .DE(_00077_),
    .Q(\w[43][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][1]$_SDFFCE_PN0P_  (.D(_01660_),
    .DE(_00077_),
    .Q(\w[43][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][20]$_SDFFCE_PN0P_  (.D(_01661_),
    .DE(_00077_),
    .Q(\w[43][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][21]$_SDFFCE_PN0P_  (.D(_01662_),
    .DE(_00077_),
    .Q(\w[43][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][22]$_SDFFCE_PN0P_  (.D(_01663_),
    .DE(_00077_),
    .Q(\w[43][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][23]$_SDFFCE_PN0P_  (.D(_01664_),
    .DE(_00077_),
    .Q(\w[43][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][24]$_SDFFCE_PN0P_  (.D(_01665_),
    .DE(_00077_),
    .Q(\w[43][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][25]$_SDFFCE_PN0P_  (.D(_01666_),
    .DE(_00077_),
    .Q(\w[43][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][26]$_SDFFCE_PN0P_  (.D(_01667_),
    .DE(_00077_),
    .Q(\w[43][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][27]$_SDFFCE_PN0P_  (.D(_01668_),
    .DE(_00077_),
    .Q(\w[43][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][28]$_SDFFCE_PN0P_  (.D(_01669_),
    .DE(_00077_),
    .Q(\w[43][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][29]$_SDFFCE_PN0P_  (.D(_01670_),
    .DE(_00077_),
    .Q(\w[43][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][2]$_SDFFCE_PN0P_  (.D(_01671_),
    .DE(_00077_),
    .Q(\w[43][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][30]$_SDFFCE_PN0P_  (.D(_01672_),
    .DE(_00077_),
    .Q(\w[43][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][31]$_SDFFCE_PN0P_  (.D(_01673_),
    .DE(_00077_),
    .Q(\w[43][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][3]$_SDFFCE_PN0P_  (.D(_01674_),
    .DE(_00077_),
    .Q(\w[43][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][4]$_SDFFCE_PN0P_  (.D(_01675_),
    .DE(_00077_),
    .Q(\w[43][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][5]$_SDFFCE_PN0P_  (.D(_01676_),
    .DE(_00077_),
    .Q(\w[43][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][6]$_SDFFCE_PN0P_  (.D(_01677_),
    .DE(_00077_),
    .Q(\w[43][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][7]$_SDFFCE_PN0P_  (.D(_01678_),
    .DE(_00077_),
    .Q(\w[43][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][8]$_SDFFCE_PN0P_  (.D(_01679_),
    .DE(_00077_),
    .Q(\w[43][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][9]$_SDFFCE_PN0P_  (.D(_01680_),
    .DE(_00077_),
    .Q(\w[43][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][0]$_SDFFCE_PN0P_  (.D(_01681_),
    .DE(_00108_),
    .Q(\w[44][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][10]$_SDFFCE_PN0P_  (.D(_01682_),
    .DE(_00108_),
    .Q(\w[44][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][11]$_SDFFCE_PN0P_  (.D(_01683_),
    .DE(_00108_),
    .Q(\w[44][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][12]$_SDFFCE_PN0P_  (.D(_01684_),
    .DE(_00108_),
    .Q(\w[44][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][13]$_SDFFCE_PN0P_  (.D(_01685_),
    .DE(_00108_),
    .Q(\w[44][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][14]$_SDFFCE_PN0P_  (.D(_01686_),
    .DE(_00108_),
    .Q(\w[44][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][15]$_SDFFCE_PN0P_  (.D(_01687_),
    .DE(_00108_),
    .Q(\w[44][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][16]$_SDFFCE_PN0P_  (.D(_01688_),
    .DE(_00108_),
    .Q(\w[44][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][17]$_SDFFCE_PN0P_  (.D(_01689_),
    .DE(_00108_),
    .Q(\w[44][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][18]$_SDFFCE_PN0P_  (.D(_01690_),
    .DE(_00108_),
    .Q(\w[44][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][19]$_SDFFCE_PN0P_  (.D(_01691_),
    .DE(_00108_),
    .Q(\w[44][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][1]$_SDFFCE_PN0P_  (.D(_01692_),
    .DE(_00108_),
    .Q(\w[44][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][20]$_SDFFCE_PN0P_  (.D(_01693_),
    .DE(_00108_),
    .Q(\w[44][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][21]$_SDFFCE_PN0P_  (.D(_01694_),
    .DE(_00108_),
    .Q(\w[44][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][22]$_SDFFCE_PN0P_  (.D(_01695_),
    .DE(_00108_),
    .Q(\w[44][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][23]$_SDFFCE_PN0P_  (.D(_01696_),
    .DE(_00108_),
    .Q(\w[44][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][24]$_SDFFCE_PN0P_  (.D(_01697_),
    .DE(_00108_),
    .Q(\w[44][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][25]$_SDFFCE_PN0P_  (.D(_01698_),
    .DE(_00108_),
    .Q(\w[44][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][26]$_SDFFCE_PN0P_  (.D(_01699_),
    .DE(_00108_),
    .Q(\w[44][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][27]$_SDFFCE_PN0P_  (.D(_01700_),
    .DE(_00108_),
    .Q(\w[44][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][28]$_SDFFCE_PN0P_  (.D(_01701_),
    .DE(_00108_),
    .Q(\w[44][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][29]$_SDFFCE_PN0P_  (.D(_01702_),
    .DE(_00108_),
    .Q(\w[44][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][2]$_SDFFCE_PN0P_  (.D(_01703_),
    .DE(_00108_),
    .Q(\w[44][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][30]$_SDFFCE_PN0P_  (.D(_01704_),
    .DE(_00108_),
    .Q(\w[44][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][31]$_SDFFCE_PN0P_  (.D(_01705_),
    .DE(_00108_),
    .Q(\w[44][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][3]$_SDFFCE_PN0P_  (.D(_01706_),
    .DE(_00108_),
    .Q(\w[44][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][4]$_SDFFCE_PN0P_  (.D(_01707_),
    .DE(_00108_),
    .Q(\w[44][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][5]$_SDFFCE_PN0P_  (.D(_01708_),
    .DE(_00108_),
    .Q(\w[44][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][6]$_SDFFCE_PN0P_  (.D(_01709_),
    .DE(_00108_),
    .Q(\w[44][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][7]$_SDFFCE_PN0P_  (.D(_01710_),
    .DE(_00108_),
    .Q(\w[44][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][8]$_SDFFCE_PN0P_  (.D(_01711_),
    .DE(_00108_),
    .Q(\w[44][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][9]$_SDFFCE_PN0P_  (.D(_01712_),
    .DE(_00108_),
    .Q(\w[44][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][0]$_SDFFCE_PN0P_  (.D(_01713_),
    .DE(_00076_),
    .Q(\w[45][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][10]$_SDFFCE_PN0P_  (.D(_01714_),
    .DE(_00076_),
    .Q(\w[45][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][11]$_SDFFCE_PN0P_  (.D(_01715_),
    .DE(_00076_),
    .Q(\w[45][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][12]$_SDFFCE_PN0P_  (.D(_01716_),
    .DE(_00076_),
    .Q(\w[45][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][13]$_SDFFCE_PN0P_  (.D(_01717_),
    .DE(_00076_),
    .Q(\w[45][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][14]$_SDFFCE_PN0P_  (.D(_01718_),
    .DE(_00076_),
    .Q(\w[45][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][15]$_SDFFCE_PN0P_  (.D(_01719_),
    .DE(_00076_),
    .Q(\w[45][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][16]$_SDFFCE_PN0P_  (.D(_01720_),
    .DE(_00076_),
    .Q(\w[45][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][17]$_SDFFCE_PN0P_  (.D(_01721_),
    .DE(_00076_),
    .Q(\w[45][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][18]$_SDFFCE_PN0P_  (.D(_01722_),
    .DE(_00076_),
    .Q(\w[45][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][19]$_SDFFCE_PN0P_  (.D(_01723_),
    .DE(_00076_),
    .Q(\w[45][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][1]$_SDFFCE_PN0P_  (.D(_01724_),
    .DE(_00076_),
    .Q(\w[45][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][20]$_SDFFCE_PN0P_  (.D(_01725_),
    .DE(_00076_),
    .Q(\w[45][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][21]$_SDFFCE_PN0P_  (.D(_01726_),
    .DE(_00076_),
    .Q(\w[45][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][22]$_SDFFCE_PN0P_  (.D(_01727_),
    .DE(_00076_),
    .Q(\w[45][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][23]$_SDFFCE_PN0P_  (.D(_01728_),
    .DE(_00076_),
    .Q(\w[45][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][24]$_SDFFCE_PN0P_  (.D(_01729_),
    .DE(_00076_),
    .Q(\w[45][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][25]$_SDFFCE_PN0P_  (.D(_01730_),
    .DE(_00076_),
    .Q(\w[45][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][26]$_SDFFCE_PN0P_  (.D(_01731_),
    .DE(_00076_),
    .Q(\w[45][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][27]$_SDFFCE_PN0P_  (.D(_01732_),
    .DE(_00076_),
    .Q(\w[45][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][28]$_SDFFCE_PN0P_  (.D(_01733_),
    .DE(_00076_),
    .Q(\w[45][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][29]$_SDFFCE_PN0P_  (.D(_01734_),
    .DE(_00076_),
    .Q(\w[45][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][2]$_SDFFCE_PN0P_  (.D(_01735_),
    .DE(_00076_),
    .Q(\w[45][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][30]$_SDFFCE_PN0P_  (.D(_01736_),
    .DE(_00076_),
    .Q(\w[45][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][31]$_SDFFCE_PN0P_  (.D(_01737_),
    .DE(_00076_),
    .Q(\w[45][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][3]$_SDFFCE_PN0P_  (.D(_01738_),
    .DE(_00076_),
    .Q(\w[45][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][4]$_SDFFCE_PN0P_  (.D(_01739_),
    .DE(_00076_),
    .Q(\w[45][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][5]$_SDFFCE_PN0P_  (.D(_01740_),
    .DE(_00076_),
    .Q(\w[45][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][6]$_SDFFCE_PN0P_  (.D(_01741_),
    .DE(_00076_),
    .Q(\w[45][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][7]$_SDFFCE_PN0P_  (.D(_01742_),
    .DE(_00076_),
    .Q(\w[45][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][8]$_SDFFCE_PN0P_  (.D(_01743_),
    .DE(_00076_),
    .Q(\w[45][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][9]$_SDFFCE_PN0P_  (.D(_01744_),
    .DE(_00076_),
    .Q(\w[45][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][0]$_SDFFCE_PN0P_  (.D(_01745_),
    .DE(_00107_),
    .Q(\w[46][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][10]$_SDFFCE_PN0P_  (.D(_01746_),
    .DE(_00107_),
    .Q(\w[46][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][11]$_SDFFCE_PN0P_  (.D(_01747_),
    .DE(_00107_),
    .Q(\w[46][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][12]$_SDFFCE_PN0P_  (.D(_01748_),
    .DE(_00107_),
    .Q(\w[46][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][13]$_SDFFCE_PN0P_  (.D(_01749_),
    .DE(_00107_),
    .Q(\w[46][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][14]$_SDFFCE_PN0P_  (.D(_01750_),
    .DE(_00107_),
    .Q(\w[46][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][15]$_SDFFCE_PN0P_  (.D(_01751_),
    .DE(_00107_),
    .Q(\w[46][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][16]$_SDFFCE_PN0P_  (.D(_01752_),
    .DE(_00107_),
    .Q(\w[46][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][17]$_SDFFCE_PN0P_  (.D(_01753_),
    .DE(_00107_),
    .Q(\w[46][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][18]$_SDFFCE_PN0P_  (.D(_01754_),
    .DE(_00107_),
    .Q(\w[46][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][19]$_SDFFCE_PN0P_  (.D(_01755_),
    .DE(_00107_),
    .Q(\w[46][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][1]$_SDFFCE_PN0P_  (.D(_01756_),
    .DE(_00107_),
    .Q(\w[46][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][20]$_SDFFCE_PN0P_  (.D(_01757_),
    .DE(_00107_),
    .Q(\w[46][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][21]$_SDFFCE_PN0P_  (.D(_01758_),
    .DE(_00107_),
    .Q(\w[46][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][22]$_SDFFCE_PN0P_  (.D(_01759_),
    .DE(_00107_),
    .Q(\w[46][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][23]$_SDFFCE_PN0P_  (.D(_01760_),
    .DE(_00107_),
    .Q(\w[46][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][24]$_SDFFCE_PN0P_  (.D(_01761_),
    .DE(_00107_),
    .Q(\w[46][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][25]$_SDFFCE_PN0P_  (.D(_01762_),
    .DE(_00107_),
    .Q(\w[46][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][26]$_SDFFCE_PN0P_  (.D(_01763_),
    .DE(_00107_),
    .Q(\w[46][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][27]$_SDFFCE_PN0P_  (.D(_01764_),
    .DE(_00107_),
    .Q(\w[46][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][28]$_SDFFCE_PN0P_  (.D(_01765_),
    .DE(_00107_),
    .Q(\w[46][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][29]$_SDFFCE_PN0P_  (.D(_01766_),
    .DE(_00107_),
    .Q(\w[46][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][2]$_SDFFCE_PN0P_  (.D(_01767_),
    .DE(_00107_),
    .Q(\w[46][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][30]$_SDFFCE_PN0P_  (.D(_01768_),
    .DE(_00107_),
    .Q(\w[46][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][31]$_SDFFCE_PN0P_  (.D(_01769_),
    .DE(_00107_),
    .Q(\w[46][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][3]$_SDFFCE_PN0P_  (.D(_01770_),
    .DE(_00107_),
    .Q(\w[46][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][4]$_SDFFCE_PN0P_  (.D(_01771_),
    .DE(_00107_),
    .Q(\w[46][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][5]$_SDFFCE_PN0P_  (.D(_01772_),
    .DE(_00107_),
    .Q(\w[46][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][6]$_SDFFCE_PN0P_  (.D(_01773_),
    .DE(_00107_),
    .Q(\w[46][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][7]$_SDFFCE_PN0P_  (.D(_01774_),
    .DE(_00107_),
    .Q(\w[46][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][8]$_SDFFCE_PN0P_  (.D(_01775_),
    .DE(_00107_),
    .Q(\w[46][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][9]$_SDFFCE_PN0P_  (.D(_01776_),
    .DE(_00107_),
    .Q(\w[46][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][0]$_SDFFCE_PN0P_  (.D(_01777_),
    .DE(_00075_),
    .Q(\w[47][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][10]$_SDFFCE_PN0P_  (.D(_01778_),
    .DE(_00075_),
    .Q(\w[47][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][11]$_SDFFCE_PN0P_  (.D(_01779_),
    .DE(_00075_),
    .Q(\w[47][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][12]$_SDFFCE_PN0P_  (.D(_01780_),
    .DE(_00075_),
    .Q(\w[47][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][13]$_SDFFCE_PN0P_  (.D(_01781_),
    .DE(_00075_),
    .Q(\w[47][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][14]$_SDFFCE_PN0P_  (.D(_01782_),
    .DE(_00075_),
    .Q(\w[47][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][15]$_SDFFCE_PN0P_  (.D(_01783_),
    .DE(_00075_),
    .Q(\w[47][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][16]$_SDFFCE_PN0P_  (.D(_01784_),
    .DE(_00075_),
    .Q(\w[47][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][17]$_SDFFCE_PN0P_  (.D(_01785_),
    .DE(_00075_),
    .Q(\w[47][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][18]$_SDFFCE_PN0P_  (.D(_01786_),
    .DE(_00075_),
    .Q(\w[47][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][19]$_SDFFCE_PN0P_  (.D(_01787_),
    .DE(_00075_),
    .Q(\w[47][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][1]$_SDFFCE_PN0P_  (.D(_01788_),
    .DE(_00075_),
    .Q(\w[47][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][20]$_SDFFCE_PN0P_  (.D(_01789_),
    .DE(_00075_),
    .Q(\w[47][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][21]$_SDFFCE_PN0P_  (.D(_01790_),
    .DE(_00075_),
    .Q(\w[47][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][22]$_SDFFCE_PN0P_  (.D(_01791_),
    .DE(_00075_),
    .Q(\w[47][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][23]$_SDFFCE_PN0P_  (.D(_01792_),
    .DE(_00075_),
    .Q(\w[47][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][24]$_SDFFCE_PN0P_  (.D(_01793_),
    .DE(_00075_),
    .Q(\w[47][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][25]$_SDFFCE_PN0P_  (.D(_01794_),
    .DE(_00075_),
    .Q(\w[47][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][26]$_SDFFCE_PN0P_  (.D(_01795_),
    .DE(_00075_),
    .Q(\w[47][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][27]$_SDFFCE_PN0P_  (.D(_01796_),
    .DE(_00075_),
    .Q(\w[47][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][28]$_SDFFCE_PN0P_  (.D(_01797_),
    .DE(_00075_),
    .Q(\w[47][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][29]$_SDFFCE_PN0P_  (.D(_01798_),
    .DE(_00075_),
    .Q(\w[47][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][2]$_SDFFCE_PN0P_  (.D(_01799_),
    .DE(_00075_),
    .Q(\w[47][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][30]$_SDFFCE_PN0P_  (.D(_01800_),
    .DE(_00075_),
    .Q(\w[47][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][31]$_SDFFCE_PN0P_  (.D(_01801_),
    .DE(_00075_),
    .Q(\w[47][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][3]$_SDFFCE_PN0P_  (.D(_01802_),
    .DE(_00075_),
    .Q(\w[47][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][4]$_SDFFCE_PN0P_  (.D(_01803_),
    .DE(_00075_),
    .Q(\w[47][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][5]$_SDFFCE_PN0P_  (.D(_01804_),
    .DE(_00075_),
    .Q(\w[47][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][6]$_SDFFCE_PN0P_  (.D(_01805_),
    .DE(_00075_),
    .Q(\w[47][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][7]$_SDFFCE_PN0P_  (.D(_01806_),
    .DE(_00075_),
    .Q(\w[47][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][8]$_SDFFCE_PN0P_  (.D(_01807_),
    .DE(_00075_),
    .Q(\w[47][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][9]$_SDFFCE_PN0P_  (.D(_01808_),
    .DE(_00075_),
    .Q(\w[47][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][0]$_SDFFCE_PN0P_  (.D(_01809_),
    .DE(_00106_),
    .Q(\w[48][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][10]$_SDFFCE_PN0P_  (.D(_01810_),
    .DE(_00106_),
    .Q(\w[48][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][11]$_SDFFCE_PN0P_  (.D(_01811_),
    .DE(_00106_),
    .Q(\w[48][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][12]$_SDFFCE_PN0P_  (.D(_01812_),
    .DE(_00106_),
    .Q(\w[48][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][13]$_SDFFCE_PN0P_  (.D(_01813_),
    .DE(_00106_),
    .Q(\w[48][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][14]$_SDFFCE_PN0P_  (.D(_01814_),
    .DE(_00106_),
    .Q(\w[48][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][15]$_SDFFCE_PN0P_  (.D(_01815_),
    .DE(_00106_),
    .Q(\w[48][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][16]$_SDFFCE_PN0P_  (.D(_01816_),
    .DE(_00106_),
    .Q(\w[48][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][17]$_SDFFCE_PN0P_  (.D(_01817_),
    .DE(_00106_),
    .Q(\w[48][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][18]$_SDFFCE_PN0P_  (.D(_01818_),
    .DE(_00106_),
    .Q(\w[48][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][19]$_SDFFCE_PN0P_  (.D(_01819_),
    .DE(_00106_),
    .Q(\w[48][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][1]$_SDFFCE_PN0P_  (.D(_01820_),
    .DE(_00106_),
    .Q(\w[48][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][20]$_SDFFCE_PN0P_  (.D(_01821_),
    .DE(_00106_),
    .Q(\w[48][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][21]$_SDFFCE_PN0P_  (.D(_01822_),
    .DE(_00106_),
    .Q(\w[48][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][22]$_SDFFCE_PN0P_  (.D(_01823_),
    .DE(_00106_),
    .Q(\w[48][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][23]$_SDFFCE_PN0P_  (.D(_01824_),
    .DE(_00106_),
    .Q(\w[48][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][24]$_SDFFCE_PN0P_  (.D(_01825_),
    .DE(_00106_),
    .Q(\w[48][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][25]$_SDFFCE_PN0P_  (.D(_01826_),
    .DE(_00106_),
    .Q(\w[48][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][26]$_SDFFCE_PN0P_  (.D(_01827_),
    .DE(_00106_),
    .Q(\w[48][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][27]$_SDFFCE_PN0P_  (.D(_01828_),
    .DE(_00106_),
    .Q(\w[48][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][28]$_SDFFCE_PN0P_  (.D(_01829_),
    .DE(_00106_),
    .Q(\w[48][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][29]$_SDFFCE_PN0P_  (.D(_01830_),
    .DE(_00106_),
    .Q(\w[48][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][2]$_SDFFCE_PN0P_  (.D(_01831_),
    .DE(_00106_),
    .Q(\w[48][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][30]$_SDFFCE_PN0P_  (.D(_01832_),
    .DE(_00106_),
    .Q(\w[48][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][31]$_SDFFCE_PN0P_  (.D(_01833_),
    .DE(_00106_),
    .Q(\w[48][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][3]$_SDFFCE_PN0P_  (.D(_01834_),
    .DE(_00106_),
    .Q(\w[48][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][4]$_SDFFCE_PN0P_  (.D(_01835_),
    .DE(_00106_),
    .Q(\w[48][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][5]$_SDFFCE_PN0P_  (.D(_01836_),
    .DE(_00106_),
    .Q(\w[48][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][6]$_SDFFCE_PN0P_  (.D(_01837_),
    .DE(_00106_),
    .Q(\w[48][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][7]$_SDFFCE_PN0P_  (.D(_01838_),
    .DE(_00106_),
    .Q(\w[48][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][8]$_SDFFCE_PN0P_  (.D(_01839_),
    .DE(_00106_),
    .Q(\w[48][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][9]$_SDFFCE_PN0P_  (.D(_01840_),
    .DE(_00106_),
    .Q(\w[48][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][0]$_SDFFCE_PN0P_  (.D(_01841_),
    .DE(_00074_),
    .Q(\w[49][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][10]$_SDFFCE_PN0P_  (.D(_01842_),
    .DE(_00074_),
    .Q(\w[49][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][11]$_SDFFCE_PN0P_  (.D(_01843_),
    .DE(_00074_),
    .Q(\w[49][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][12]$_SDFFCE_PN0P_  (.D(_01844_),
    .DE(_00074_),
    .Q(\w[49][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][13]$_SDFFCE_PN0P_  (.D(_01845_),
    .DE(_00074_),
    .Q(\w[49][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][14]$_SDFFCE_PN0P_  (.D(_01846_),
    .DE(_00074_),
    .Q(\w[49][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][15]$_SDFFCE_PN0P_  (.D(_01847_),
    .DE(_00074_),
    .Q(\w[49][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][16]$_SDFFCE_PN0P_  (.D(_01848_),
    .DE(_00074_),
    .Q(\w[49][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][17]$_SDFFCE_PN0P_  (.D(_01849_),
    .DE(_00074_),
    .Q(\w[49][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][18]$_SDFFCE_PN0P_  (.D(_01850_),
    .DE(_00074_),
    .Q(\w[49][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][19]$_SDFFCE_PN0P_  (.D(_01851_),
    .DE(_00074_),
    .Q(\w[49][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][1]$_SDFFCE_PN0P_  (.D(_01852_),
    .DE(_00074_),
    .Q(\w[49][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][20]$_SDFFCE_PN0P_  (.D(_01853_),
    .DE(_00074_),
    .Q(\w[49][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][21]$_SDFFCE_PN0P_  (.D(_01854_),
    .DE(_00074_),
    .Q(\w[49][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][22]$_SDFFCE_PN0P_  (.D(_01855_),
    .DE(_00074_),
    .Q(\w[49][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][23]$_SDFFCE_PN0P_  (.D(_01856_),
    .DE(_00074_),
    .Q(\w[49][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][24]$_SDFFCE_PN0P_  (.D(_01857_),
    .DE(_00074_),
    .Q(\w[49][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][25]$_SDFFCE_PN0P_  (.D(_01858_),
    .DE(_00074_),
    .Q(\w[49][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][26]$_SDFFCE_PN0P_  (.D(_01859_),
    .DE(_00074_),
    .Q(\w[49][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][27]$_SDFFCE_PN0P_  (.D(_01860_),
    .DE(_00074_),
    .Q(\w[49][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][28]$_SDFFCE_PN0P_  (.D(_01861_),
    .DE(_00074_),
    .Q(\w[49][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][29]$_SDFFCE_PN0P_  (.D(_01862_),
    .DE(_00074_),
    .Q(\w[49][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][2]$_SDFFCE_PN0P_  (.D(_01863_),
    .DE(_00074_),
    .Q(\w[49][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][30]$_SDFFCE_PN0P_  (.D(_01864_),
    .DE(_00074_),
    .Q(\w[49][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][31]$_SDFFCE_PN0P_  (.D(_01865_),
    .DE(_00074_),
    .Q(\w[49][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][3]$_SDFFCE_PN0P_  (.D(_01866_),
    .DE(_00074_),
    .Q(\w[49][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][4]$_SDFFCE_PN0P_  (.D(_01867_),
    .DE(_00074_),
    .Q(\w[49][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][5]$_SDFFCE_PN0P_  (.D(_01868_),
    .DE(_00074_),
    .Q(\w[49][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][6]$_SDFFCE_PN0P_  (.D(_01869_),
    .DE(_00074_),
    .Q(\w[49][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][7]$_SDFFCE_PN0P_  (.D(_01870_),
    .DE(_00074_),
    .Q(\w[49][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][8]$_SDFFCE_PN0P_  (.D(_01871_),
    .DE(_00074_),
    .Q(\w[49][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][9]$_SDFFCE_PN0P_  (.D(_01872_),
    .DE(_00074_),
    .Q(\w[49][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][0]$_DFFE_PP_  (.D(_00449_),
    .DE(_00105_),
    .Q(\w[4][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][10]$_DFFE_PP_  (.D(_00450_),
    .DE(_00105_),
    .Q(\w[4][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][11]$_DFFE_PP_  (.D(_00451_),
    .DE(_00105_),
    .Q(\w[4][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][12]$_DFFE_PP_  (.D(_00452_),
    .DE(_00105_),
    .Q(\w[4][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][13]$_DFFE_PP_  (.D(_00453_),
    .DE(_00105_),
    .Q(\w[4][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][14]$_DFFE_PP_  (.D(_00454_),
    .DE(_00105_),
    .Q(\w[4][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][15]$_DFFE_PP_  (.D(_00455_),
    .DE(_00105_),
    .Q(\w[4][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][16]$_DFFE_PP_  (.D(_00456_),
    .DE(_00105_),
    .Q(\w[4][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][17]$_DFFE_PP_  (.D(_00457_),
    .DE(_00105_),
    .Q(\w[4][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][18]$_DFFE_PP_  (.D(_00458_),
    .DE(_00105_),
    .Q(\w[4][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][19]$_DFFE_PP_  (.D(_00459_),
    .DE(_00105_),
    .Q(\w[4][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][1]$_DFFE_PP_  (.D(_00460_),
    .DE(_00105_),
    .Q(\w[4][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][20]$_DFFE_PP_  (.D(_00461_),
    .DE(_00105_),
    .Q(\w[4][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][21]$_DFFE_PP_  (.D(_00462_),
    .DE(_00105_),
    .Q(\w[4][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][22]$_DFFE_PP_  (.D(_00463_),
    .DE(_00105_),
    .Q(\w[4][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][23]$_DFFE_PP_  (.D(_00464_),
    .DE(_00105_),
    .Q(\w[4][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][24]$_DFFE_PP_  (.D(_00465_),
    .DE(_00105_),
    .Q(\w[4][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][25]$_DFFE_PP_  (.D(_00466_),
    .DE(_00105_),
    .Q(\w[4][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][26]$_DFFE_PP_  (.D(_00467_),
    .DE(_00105_),
    .Q(\w[4][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][27]$_DFFE_PP_  (.D(_00468_),
    .DE(_00105_),
    .Q(\w[4][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][28]$_DFFE_PP_  (.D(_00469_),
    .DE(_00105_),
    .Q(\w[4][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][29]$_DFFE_PP_  (.D(_00470_),
    .DE(_00105_),
    .Q(\w[4][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][2]$_DFFE_PP_  (.D(_00471_),
    .DE(_00105_),
    .Q(\w[4][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][30]$_DFFE_PP_  (.D(_00472_),
    .DE(_00105_),
    .Q(\w[4][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][31]$_DFFE_PP_  (.D(_00473_),
    .DE(_00105_),
    .Q(\w[4][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][3]$_DFFE_PP_  (.D(_00474_),
    .DE(_00105_),
    .Q(\w[4][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][4]$_DFFE_PP_  (.D(_00475_),
    .DE(_00105_),
    .Q(\w[4][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][5]$_DFFE_PP_  (.D(_00476_),
    .DE(_00105_),
    .Q(\w[4][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][6]$_DFFE_PP_  (.D(_00477_),
    .DE(_00105_),
    .Q(\w[4][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][7]$_DFFE_PP_  (.D(_00478_),
    .DE(_00105_),
    .Q(\w[4][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][8]$_DFFE_PP_  (.D(_00479_),
    .DE(_00105_),
    .Q(\w[4][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][9]$_DFFE_PP_  (.D(_00480_),
    .DE(_00105_),
    .Q(\w[4][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][0]$_SDFFCE_PN0P_  (.D(_01873_),
    .DE(_00104_),
    .Q(\w[50][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][10]$_SDFFCE_PN0P_  (.D(_01874_),
    .DE(_00104_),
    .Q(\w[50][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][11]$_SDFFCE_PN0P_  (.D(_01875_),
    .DE(_00104_),
    .Q(\w[50][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][12]$_SDFFCE_PN0P_  (.D(_01876_),
    .DE(_00104_),
    .Q(\w[50][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][13]$_SDFFCE_PN0P_  (.D(_01877_),
    .DE(_00104_),
    .Q(\w[50][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][14]$_SDFFCE_PN0P_  (.D(_01878_),
    .DE(_00104_),
    .Q(\w[50][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][15]$_SDFFCE_PN0P_  (.D(_01879_),
    .DE(_00104_),
    .Q(\w[50][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][16]$_SDFFCE_PN0P_  (.D(_01880_),
    .DE(_00104_),
    .Q(\w[50][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][17]$_SDFFCE_PN0P_  (.D(_01881_),
    .DE(_00104_),
    .Q(\w[50][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][18]$_SDFFCE_PN0P_  (.D(_01882_),
    .DE(_00104_),
    .Q(\w[50][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][19]$_SDFFCE_PN0P_  (.D(_01883_),
    .DE(_00104_),
    .Q(\w[50][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][1]$_SDFFCE_PN0P_  (.D(_01884_),
    .DE(_00104_),
    .Q(\w[50][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][20]$_SDFFCE_PN0P_  (.D(_01885_),
    .DE(_00104_),
    .Q(\w[50][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][21]$_SDFFCE_PN0P_  (.D(_01886_),
    .DE(_00104_),
    .Q(\w[50][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][22]$_SDFFCE_PN0P_  (.D(_01887_),
    .DE(_00104_),
    .Q(\w[50][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][23]$_SDFFCE_PN0P_  (.D(_01888_),
    .DE(_00104_),
    .Q(\w[50][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][24]$_SDFFCE_PN0P_  (.D(_01889_),
    .DE(_00104_),
    .Q(\w[50][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][25]$_SDFFCE_PN0P_  (.D(_01890_),
    .DE(_00104_),
    .Q(\w[50][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][26]$_SDFFCE_PN0P_  (.D(_01891_),
    .DE(_00104_),
    .Q(\w[50][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][27]$_SDFFCE_PN0P_  (.D(_01892_),
    .DE(_00104_),
    .Q(\w[50][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][28]$_SDFFCE_PN0P_  (.D(_01893_),
    .DE(_00104_),
    .Q(\w[50][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][29]$_SDFFCE_PN0P_  (.D(_01894_),
    .DE(_00104_),
    .Q(\w[50][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][2]$_SDFFCE_PN0P_  (.D(_01895_),
    .DE(_00104_),
    .Q(\w[50][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][30]$_SDFFCE_PN0P_  (.D(_01896_),
    .DE(_00104_),
    .Q(\w[50][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][31]$_SDFFCE_PN0P_  (.D(_01897_),
    .DE(_00104_),
    .Q(\w[50][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][3]$_SDFFCE_PN0P_  (.D(_01898_),
    .DE(_00104_),
    .Q(\w[50][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][4]$_SDFFCE_PN0P_  (.D(_01899_),
    .DE(_00104_),
    .Q(\w[50][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][5]$_SDFFCE_PN0P_  (.D(_01900_),
    .DE(_00104_),
    .Q(\w[50][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][6]$_SDFFCE_PN0P_  (.D(_01901_),
    .DE(_00104_),
    .Q(\w[50][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][7]$_SDFFCE_PN0P_  (.D(_01902_),
    .DE(_00104_),
    .Q(\w[50][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][8]$_SDFFCE_PN0P_  (.D(_01903_),
    .DE(_00104_),
    .Q(\w[50][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][9]$_SDFFCE_PN0P_  (.D(_01904_),
    .DE(_00104_),
    .Q(\w[50][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][0]$_SDFFCE_PN0P_  (.D(_01905_),
    .DE(_00073_),
    .Q(\w[51][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][10]$_SDFFCE_PN0P_  (.D(_01906_),
    .DE(_00073_),
    .Q(\w[51][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][11]$_SDFFCE_PN0P_  (.D(_01907_),
    .DE(_00073_),
    .Q(\w[51][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][12]$_SDFFCE_PN0P_  (.D(_01908_),
    .DE(_00073_),
    .Q(\w[51][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][13]$_SDFFCE_PN0P_  (.D(_01909_),
    .DE(_00073_),
    .Q(\w[51][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][14]$_SDFFCE_PN0P_  (.D(_01910_),
    .DE(_00073_),
    .Q(\w[51][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][15]$_SDFFCE_PN0P_  (.D(_01911_),
    .DE(_00073_),
    .Q(\w[51][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][16]$_SDFFCE_PN0P_  (.D(_01912_),
    .DE(_00073_),
    .Q(\w[51][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][17]$_SDFFCE_PN0P_  (.D(_01913_),
    .DE(_00073_),
    .Q(\w[51][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][18]$_SDFFCE_PN0P_  (.D(_01914_),
    .DE(_00073_),
    .Q(\w[51][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][19]$_SDFFCE_PN0P_  (.D(_01915_),
    .DE(_00073_),
    .Q(\w[51][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][1]$_SDFFCE_PN0P_  (.D(_01916_),
    .DE(_00073_),
    .Q(\w[51][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][20]$_SDFFCE_PN0P_  (.D(_01917_),
    .DE(_00073_),
    .Q(\w[51][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][21]$_SDFFCE_PN0P_  (.D(_01918_),
    .DE(_00073_),
    .Q(\w[51][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][22]$_SDFFCE_PN0P_  (.D(_01919_),
    .DE(_00073_),
    .Q(\w[51][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][23]$_SDFFCE_PN0P_  (.D(_01920_),
    .DE(_00073_),
    .Q(\w[51][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][24]$_SDFFCE_PN0P_  (.D(_01921_),
    .DE(_00073_),
    .Q(\w[51][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][25]$_SDFFCE_PN0P_  (.D(_01922_),
    .DE(_00073_),
    .Q(\w[51][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][26]$_SDFFCE_PN0P_  (.D(_01923_),
    .DE(_00073_),
    .Q(\w[51][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][27]$_SDFFCE_PN0P_  (.D(_01924_),
    .DE(_00073_),
    .Q(\w[51][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][28]$_SDFFCE_PN0P_  (.D(_01925_),
    .DE(_00073_),
    .Q(\w[51][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][29]$_SDFFCE_PN0P_  (.D(_01926_),
    .DE(_00073_),
    .Q(\w[51][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][2]$_SDFFCE_PN0P_  (.D(_01927_),
    .DE(_00073_),
    .Q(\w[51][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][30]$_SDFFCE_PN0P_  (.D(_01928_),
    .DE(_00073_),
    .Q(\w[51][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][31]$_SDFFCE_PN0P_  (.D(_01929_),
    .DE(_00073_),
    .Q(\w[51][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][3]$_SDFFCE_PN0P_  (.D(_01930_),
    .DE(_00073_),
    .Q(\w[51][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][4]$_SDFFCE_PN0P_  (.D(_01931_),
    .DE(_00073_),
    .Q(\w[51][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][5]$_SDFFCE_PN0P_  (.D(_01932_),
    .DE(_00073_),
    .Q(\w[51][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][6]$_SDFFCE_PN0P_  (.D(_01933_),
    .DE(_00073_),
    .Q(\w[51][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][7]$_SDFFCE_PN0P_  (.D(_01934_),
    .DE(_00073_),
    .Q(\w[51][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][8]$_SDFFCE_PN0P_  (.D(_01935_),
    .DE(_00073_),
    .Q(\w[51][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][9]$_SDFFCE_PN0P_  (.D(_01936_),
    .DE(_00073_),
    .Q(\w[51][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][0]$_SDFFCE_PN0P_  (.D(_01937_),
    .DE(_00103_),
    .Q(\w[52][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][10]$_SDFFCE_PN0P_  (.D(_01938_),
    .DE(_00103_),
    .Q(\w[52][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][11]$_SDFFCE_PN0P_  (.D(_01939_),
    .DE(_00103_),
    .Q(\w[52][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][12]$_SDFFCE_PN0P_  (.D(_01940_),
    .DE(_00103_),
    .Q(\w[52][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][13]$_SDFFCE_PN0P_  (.D(_01941_),
    .DE(_00103_),
    .Q(\w[52][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][14]$_SDFFCE_PN0P_  (.D(_01942_),
    .DE(_00103_),
    .Q(\w[52][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][15]$_SDFFCE_PN0P_  (.D(_01943_),
    .DE(_00103_),
    .Q(\w[52][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][16]$_SDFFCE_PN0P_  (.D(_01944_),
    .DE(_00103_),
    .Q(\w[52][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][17]$_SDFFCE_PN0P_  (.D(_01945_),
    .DE(_00103_),
    .Q(\w[52][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][18]$_SDFFCE_PN0P_  (.D(_01946_),
    .DE(_00103_),
    .Q(\w[52][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][19]$_SDFFCE_PN0P_  (.D(_01947_),
    .DE(_00103_),
    .Q(\w[52][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][1]$_SDFFCE_PN0P_  (.D(_01948_),
    .DE(_00103_),
    .Q(\w[52][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][20]$_SDFFCE_PN0P_  (.D(_01949_),
    .DE(_00103_),
    .Q(\w[52][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][21]$_SDFFCE_PN0P_  (.D(_01950_),
    .DE(_00103_),
    .Q(\w[52][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][22]$_SDFFCE_PN0P_  (.D(_01951_),
    .DE(_00103_),
    .Q(\w[52][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][23]$_SDFFCE_PN0P_  (.D(_01952_),
    .DE(_00103_),
    .Q(\w[52][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][24]$_SDFFCE_PN0P_  (.D(_01953_),
    .DE(_00103_),
    .Q(\w[52][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][25]$_SDFFCE_PN0P_  (.D(_01954_),
    .DE(_00103_),
    .Q(\w[52][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][26]$_SDFFCE_PN0P_  (.D(_01955_),
    .DE(_00103_),
    .Q(\w[52][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][27]$_SDFFCE_PN0P_  (.D(_01956_),
    .DE(_00103_),
    .Q(\w[52][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][28]$_SDFFCE_PN0P_  (.D(_01957_),
    .DE(_00103_),
    .Q(\w[52][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][29]$_SDFFCE_PN0P_  (.D(_01958_),
    .DE(_00103_),
    .Q(\w[52][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][2]$_SDFFCE_PN0P_  (.D(_01959_),
    .DE(_00103_),
    .Q(\w[52][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][30]$_SDFFCE_PN0P_  (.D(_01960_),
    .DE(_00103_),
    .Q(\w[52][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][31]$_SDFFCE_PN0P_  (.D(_01961_),
    .DE(_00103_),
    .Q(\w[52][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][3]$_SDFFCE_PN0P_  (.D(_01962_),
    .DE(_00103_),
    .Q(\w[52][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][4]$_SDFFCE_PN0P_  (.D(_01963_),
    .DE(_00103_),
    .Q(\w[52][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][5]$_SDFFCE_PN0P_  (.D(_01964_),
    .DE(_00103_),
    .Q(\w[52][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][6]$_SDFFCE_PN0P_  (.D(_01965_),
    .DE(_00103_),
    .Q(\w[52][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][7]$_SDFFCE_PN0P_  (.D(_01966_),
    .DE(_00103_),
    .Q(\w[52][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][8]$_SDFFCE_PN0P_  (.D(_01967_),
    .DE(_00103_),
    .Q(\w[52][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][9]$_SDFFCE_PN0P_  (.D(_01968_),
    .DE(_00103_),
    .Q(\w[52][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][0]$_SDFFCE_PN0P_  (.D(_01969_),
    .DE(_00072_),
    .Q(\w[53][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][10]$_SDFFCE_PN0P_  (.D(_01970_),
    .DE(_00072_),
    .Q(\w[53][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][11]$_SDFFCE_PN0P_  (.D(_01971_),
    .DE(_00072_),
    .Q(\w[53][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][12]$_SDFFCE_PN0P_  (.D(_01972_),
    .DE(_00072_),
    .Q(\w[53][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][13]$_SDFFCE_PN0P_  (.D(_01973_),
    .DE(_00072_),
    .Q(\w[53][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][14]$_SDFFCE_PN0P_  (.D(_01974_),
    .DE(_00072_),
    .Q(\w[53][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][15]$_SDFFCE_PN0P_  (.D(_01975_),
    .DE(_00072_),
    .Q(\w[53][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][16]$_SDFFCE_PN0P_  (.D(_01976_),
    .DE(_00072_),
    .Q(\w[53][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][17]$_SDFFCE_PN0P_  (.D(_01977_),
    .DE(_00072_),
    .Q(\w[53][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][18]$_SDFFCE_PN0P_  (.D(_01978_),
    .DE(_00072_),
    .Q(\w[53][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][19]$_SDFFCE_PN0P_  (.D(_01979_),
    .DE(_00072_),
    .Q(\w[53][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][1]$_SDFFCE_PN0P_  (.D(_01980_),
    .DE(_00072_),
    .Q(\w[53][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][20]$_SDFFCE_PN0P_  (.D(_01981_),
    .DE(_00072_),
    .Q(\w[53][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][21]$_SDFFCE_PN0P_  (.D(_01982_),
    .DE(_00072_),
    .Q(\w[53][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][22]$_SDFFCE_PN0P_  (.D(_01983_),
    .DE(_00072_),
    .Q(\w[53][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][23]$_SDFFCE_PN0P_  (.D(_01984_),
    .DE(_00072_),
    .Q(\w[53][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][24]$_SDFFCE_PN0P_  (.D(_01985_),
    .DE(_00072_),
    .Q(\w[53][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][25]$_SDFFCE_PN0P_  (.D(_01986_),
    .DE(_00072_),
    .Q(\w[53][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][26]$_SDFFCE_PN0P_  (.D(_01987_),
    .DE(_00072_),
    .Q(\w[53][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][27]$_SDFFCE_PN0P_  (.D(_01988_),
    .DE(_00072_),
    .Q(\w[53][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][28]$_SDFFCE_PN0P_  (.D(_01989_),
    .DE(_00072_),
    .Q(\w[53][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][29]$_SDFFCE_PN0P_  (.D(_01990_),
    .DE(_00072_),
    .Q(\w[53][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][2]$_SDFFCE_PN0P_  (.D(_01991_),
    .DE(_00072_),
    .Q(\w[53][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][30]$_SDFFCE_PN0P_  (.D(_01992_),
    .DE(_00072_),
    .Q(\w[53][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][31]$_SDFFCE_PN0P_  (.D(_01993_),
    .DE(_00072_),
    .Q(\w[53][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][3]$_SDFFCE_PN0P_  (.D(_01994_),
    .DE(_00072_),
    .Q(\w[53][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][4]$_SDFFCE_PN0P_  (.D(_01995_),
    .DE(_00072_),
    .Q(\w[53][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][5]$_SDFFCE_PN0P_  (.D(_01996_),
    .DE(_00072_),
    .Q(\w[53][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][6]$_SDFFCE_PN0P_  (.D(_01997_),
    .DE(_00072_),
    .Q(\w[53][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][7]$_SDFFCE_PN0P_  (.D(_01998_),
    .DE(_00072_),
    .Q(\w[53][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][8]$_SDFFCE_PN0P_  (.D(_01999_),
    .DE(_00072_),
    .Q(\w[53][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][9]$_SDFFCE_PN0P_  (.D(_02000_),
    .DE(_00072_),
    .Q(\w[53][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][0]$_SDFFCE_PN0P_  (.D(_02001_),
    .DE(_00102_),
    .Q(\w[54][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][10]$_SDFFCE_PN0P_  (.D(_02002_),
    .DE(_00102_),
    .Q(\w[54][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][11]$_SDFFCE_PN0P_  (.D(_02003_),
    .DE(_00102_),
    .Q(\w[54][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][12]$_SDFFCE_PN0P_  (.D(_02004_),
    .DE(_00102_),
    .Q(\w[54][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][13]$_SDFFCE_PN0P_  (.D(_02005_),
    .DE(_00102_),
    .Q(\w[54][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][14]$_SDFFCE_PN0P_  (.D(_02006_),
    .DE(_00102_),
    .Q(\w[54][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][15]$_SDFFCE_PN0P_  (.D(_02007_),
    .DE(_00102_),
    .Q(\w[54][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][16]$_SDFFCE_PN0P_  (.D(_02008_),
    .DE(_00102_),
    .Q(\w[54][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][17]$_SDFFCE_PN0P_  (.D(_02009_),
    .DE(_00102_),
    .Q(\w[54][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][18]$_SDFFCE_PN0P_  (.D(_02010_),
    .DE(_00102_),
    .Q(\w[54][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][19]$_SDFFCE_PN0P_  (.D(_02011_),
    .DE(_00102_),
    .Q(\w[54][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][1]$_SDFFCE_PN0P_  (.D(_02012_),
    .DE(_00102_),
    .Q(\w[54][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][20]$_SDFFCE_PN0P_  (.D(_02013_),
    .DE(_00102_),
    .Q(\w[54][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][21]$_SDFFCE_PN0P_  (.D(_02014_),
    .DE(_00102_),
    .Q(\w[54][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][22]$_SDFFCE_PN0P_  (.D(_02015_),
    .DE(_00102_),
    .Q(\w[54][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][23]$_SDFFCE_PN0P_  (.D(_02016_),
    .DE(_00102_),
    .Q(\w[54][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][24]$_SDFFCE_PN0P_  (.D(_02017_),
    .DE(_00102_),
    .Q(\w[54][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][25]$_SDFFCE_PN0P_  (.D(_02018_),
    .DE(_00102_),
    .Q(\w[54][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][26]$_SDFFCE_PN0P_  (.D(_02019_),
    .DE(_00102_),
    .Q(\w[54][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][27]$_SDFFCE_PN0P_  (.D(_02020_),
    .DE(_00102_),
    .Q(\w[54][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][28]$_SDFFCE_PN0P_  (.D(_02021_),
    .DE(_00102_),
    .Q(\w[54][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][29]$_SDFFCE_PN0P_  (.D(_02022_),
    .DE(_00102_),
    .Q(\w[54][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][2]$_SDFFCE_PN0P_  (.D(_02023_),
    .DE(_00102_),
    .Q(\w[54][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][30]$_SDFFCE_PN0P_  (.D(_02024_),
    .DE(_00102_),
    .Q(\w[54][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][31]$_SDFFCE_PN0P_  (.D(_02025_),
    .DE(_00102_),
    .Q(\w[54][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][3]$_SDFFCE_PN0P_  (.D(_02026_),
    .DE(_00102_),
    .Q(\w[54][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][4]$_SDFFCE_PN0P_  (.D(_02027_),
    .DE(_00102_),
    .Q(\w[54][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][5]$_SDFFCE_PN0P_  (.D(_02028_),
    .DE(_00102_),
    .Q(\w[54][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][6]$_SDFFCE_PN0P_  (.D(_02029_),
    .DE(_00102_),
    .Q(\w[54][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][7]$_SDFFCE_PN0P_  (.D(_02030_),
    .DE(_00102_),
    .Q(\w[54][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][8]$_SDFFCE_PN0P_  (.D(_02031_),
    .DE(_00102_),
    .Q(\w[54][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][9]$_SDFFCE_PN0P_  (.D(_02032_),
    .DE(_00102_),
    .Q(\w[54][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][0]$_SDFFCE_PN0P_  (.D(_02033_),
    .DE(_00071_),
    .Q(\w[55][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][10]$_SDFFCE_PN0P_  (.D(_02034_),
    .DE(_00071_),
    .Q(\w[55][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][11]$_SDFFCE_PN0P_  (.D(_02035_),
    .DE(_00071_),
    .Q(\w[55][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][12]$_SDFFCE_PN0P_  (.D(_02036_),
    .DE(_00071_),
    .Q(\w[55][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][13]$_SDFFCE_PN0P_  (.D(_02037_),
    .DE(_00071_),
    .Q(\w[55][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][14]$_SDFFCE_PN0P_  (.D(_02038_),
    .DE(_00071_),
    .Q(\w[55][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][15]$_SDFFCE_PN0P_  (.D(_02039_),
    .DE(_00071_),
    .Q(\w[55][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][16]$_SDFFCE_PN0P_  (.D(_02040_),
    .DE(_00071_),
    .Q(\w[55][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][17]$_SDFFCE_PN0P_  (.D(_02041_),
    .DE(_00071_),
    .Q(\w[55][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][18]$_SDFFCE_PN0P_  (.D(_02042_),
    .DE(_00071_),
    .Q(\w[55][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][19]$_SDFFCE_PN0P_  (.D(_02043_),
    .DE(_00071_),
    .Q(\w[55][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][1]$_SDFFCE_PN0P_  (.D(_02044_),
    .DE(_00071_),
    .Q(\w[55][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][20]$_SDFFCE_PN0P_  (.D(_02045_),
    .DE(_00071_),
    .Q(\w[55][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][21]$_SDFFCE_PN0P_  (.D(_02046_),
    .DE(_00071_),
    .Q(\w[55][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][22]$_SDFFCE_PN0P_  (.D(_02047_),
    .DE(_00071_),
    .Q(\w[55][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][23]$_SDFFCE_PN0P_  (.D(_02048_),
    .DE(_00071_),
    .Q(\w[55][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][24]$_SDFFCE_PN0P_  (.D(_02049_),
    .DE(_00071_),
    .Q(\w[55][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][25]$_SDFFCE_PN0P_  (.D(_02050_),
    .DE(_00071_),
    .Q(\w[55][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][26]$_SDFFCE_PN0P_  (.D(_02051_),
    .DE(_00071_),
    .Q(\w[55][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][27]$_SDFFCE_PN0P_  (.D(_02052_),
    .DE(_00071_),
    .Q(\w[55][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][28]$_SDFFCE_PN0P_  (.D(_02053_),
    .DE(_00071_),
    .Q(\w[55][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][29]$_SDFFCE_PN0P_  (.D(_02054_),
    .DE(_00071_),
    .Q(\w[55][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][2]$_SDFFCE_PN0P_  (.D(_02055_),
    .DE(_00071_),
    .Q(\w[55][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][30]$_SDFFCE_PN0P_  (.D(_02056_),
    .DE(_00071_),
    .Q(\w[55][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][31]$_SDFFCE_PN0P_  (.D(_02057_),
    .DE(_00071_),
    .Q(\w[55][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][3]$_SDFFCE_PN0P_  (.D(_02058_),
    .DE(_00071_),
    .Q(\w[55][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][4]$_SDFFCE_PN0P_  (.D(_02059_),
    .DE(_00071_),
    .Q(\w[55][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][5]$_SDFFCE_PN0P_  (.D(_02060_),
    .DE(_00071_),
    .Q(\w[55][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][6]$_SDFFCE_PN0P_  (.D(_02061_),
    .DE(_00071_),
    .Q(\w[55][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][7]$_SDFFCE_PN0P_  (.D(_02062_),
    .DE(_00071_),
    .Q(\w[55][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][8]$_SDFFCE_PN0P_  (.D(_02063_),
    .DE(_00071_),
    .Q(\w[55][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][9]$_SDFFCE_PN0P_  (.D(_02064_),
    .DE(_00071_),
    .Q(\w[55][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][0]$_SDFFCE_PN0P_  (.D(_02065_),
    .DE(_00101_),
    .Q(\w[56][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][10]$_SDFFCE_PN0P_  (.D(_02066_),
    .DE(_00101_),
    .Q(\w[56][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][11]$_SDFFCE_PN0P_  (.D(_02067_),
    .DE(_00101_),
    .Q(\w[56][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][12]$_SDFFCE_PN0P_  (.D(_02068_),
    .DE(_00101_),
    .Q(\w[56][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][13]$_SDFFCE_PN0P_  (.D(_02069_),
    .DE(_00101_),
    .Q(\w[56][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][14]$_SDFFCE_PN0P_  (.D(_02070_),
    .DE(_00101_),
    .Q(\w[56][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][15]$_SDFFCE_PN0P_  (.D(_02071_),
    .DE(_00101_),
    .Q(\w[56][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][16]$_SDFFCE_PN0P_  (.D(_02072_),
    .DE(_00101_),
    .Q(\w[56][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][17]$_SDFFCE_PN0P_  (.D(_02073_),
    .DE(_00101_),
    .Q(\w[56][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][18]$_SDFFCE_PN0P_  (.D(_02074_),
    .DE(_00101_),
    .Q(\w[56][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][19]$_SDFFCE_PN0P_  (.D(_02075_),
    .DE(_00101_),
    .Q(\w[56][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][1]$_SDFFCE_PN0P_  (.D(_02076_),
    .DE(_00101_),
    .Q(\w[56][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][20]$_SDFFCE_PN0P_  (.D(_02077_),
    .DE(_00101_),
    .Q(\w[56][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][21]$_SDFFCE_PN0P_  (.D(_02078_),
    .DE(_00101_),
    .Q(\w[56][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][22]$_SDFFCE_PN0P_  (.D(_02079_),
    .DE(_00101_),
    .Q(\w[56][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][23]$_SDFFCE_PN0P_  (.D(_02080_),
    .DE(_00101_),
    .Q(\w[56][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][24]$_SDFFCE_PN0P_  (.D(_02081_),
    .DE(_00101_),
    .Q(\w[56][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][25]$_SDFFCE_PN0P_  (.D(_02082_),
    .DE(_00101_),
    .Q(\w[56][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][26]$_SDFFCE_PN0P_  (.D(_02083_),
    .DE(_00101_),
    .Q(\w[56][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][27]$_SDFFCE_PN0P_  (.D(_02084_),
    .DE(_00101_),
    .Q(\w[56][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][28]$_SDFFCE_PN0P_  (.D(_02085_),
    .DE(_00101_),
    .Q(\w[56][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][29]$_SDFFCE_PN0P_  (.D(_02086_),
    .DE(_00101_),
    .Q(\w[56][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][2]$_SDFFCE_PN0P_  (.D(_02087_),
    .DE(_00101_),
    .Q(\w[56][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][30]$_SDFFCE_PN0P_  (.D(_02088_),
    .DE(_00101_),
    .Q(\w[56][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][31]$_SDFFCE_PN0P_  (.D(_02089_),
    .DE(_00101_),
    .Q(\w[56][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][3]$_SDFFCE_PN0P_  (.D(_02090_),
    .DE(_00101_),
    .Q(\w[56][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][4]$_SDFFCE_PN0P_  (.D(_02091_),
    .DE(_00101_),
    .Q(\w[56][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][5]$_SDFFCE_PN0P_  (.D(_02092_),
    .DE(_00101_),
    .Q(\w[56][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][6]$_SDFFCE_PN0P_  (.D(_02093_),
    .DE(_00101_),
    .Q(\w[56][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][7]$_SDFFCE_PN0P_  (.D(_02094_),
    .DE(_00101_),
    .Q(\w[56][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][8]$_SDFFCE_PN0P_  (.D(_02095_),
    .DE(_00101_),
    .Q(\w[56][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][9]$_SDFFCE_PN0P_  (.D(_02096_),
    .DE(_00101_),
    .Q(\w[56][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][0]$_SDFFCE_PN0P_  (.D(_02097_),
    .DE(_00070_),
    .Q(\w[57][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][10]$_SDFFCE_PN0P_  (.D(_02098_),
    .DE(_00070_),
    .Q(\w[57][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][11]$_SDFFCE_PN0P_  (.D(_02099_),
    .DE(_00070_),
    .Q(\w[57][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][12]$_SDFFCE_PN0P_  (.D(_02100_),
    .DE(_00070_),
    .Q(\w[57][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][13]$_SDFFCE_PN0P_  (.D(_02101_),
    .DE(_00070_),
    .Q(\w[57][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][14]$_SDFFCE_PN0P_  (.D(_02102_),
    .DE(_00070_),
    .Q(\w[57][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][15]$_SDFFCE_PN0P_  (.D(_02103_),
    .DE(_00070_),
    .Q(\w[57][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][16]$_SDFFCE_PN0P_  (.D(_02104_),
    .DE(_00070_),
    .Q(\w[57][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][17]$_SDFFCE_PN0P_  (.D(_02105_),
    .DE(_00070_),
    .Q(\w[57][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][18]$_SDFFCE_PN0P_  (.D(_02106_),
    .DE(_00070_),
    .Q(\w[57][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][19]$_SDFFCE_PN0P_  (.D(_02107_),
    .DE(_00070_),
    .Q(\w[57][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][1]$_SDFFCE_PN0P_  (.D(_02108_),
    .DE(_00070_),
    .Q(\w[57][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][20]$_SDFFCE_PN0P_  (.D(_02109_),
    .DE(_00070_),
    .Q(\w[57][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][21]$_SDFFCE_PN0P_  (.D(_02110_),
    .DE(_00070_),
    .Q(\w[57][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][22]$_SDFFCE_PN0P_  (.D(_02111_),
    .DE(_00070_),
    .Q(\w[57][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][23]$_SDFFCE_PN0P_  (.D(_02112_),
    .DE(_00070_),
    .Q(\w[57][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][24]$_SDFFCE_PN0P_  (.D(_02113_),
    .DE(_00070_),
    .Q(\w[57][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][25]$_SDFFCE_PN0P_  (.D(_02114_),
    .DE(_00070_),
    .Q(\w[57][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][26]$_SDFFCE_PN0P_  (.D(_02115_),
    .DE(_00070_),
    .Q(\w[57][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][27]$_SDFFCE_PN0P_  (.D(_02116_),
    .DE(_00070_),
    .Q(\w[57][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][28]$_SDFFCE_PN0P_  (.D(_02117_),
    .DE(_00070_),
    .Q(\w[57][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][29]$_SDFFCE_PN0P_  (.D(_02118_),
    .DE(_00070_),
    .Q(\w[57][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][2]$_SDFFCE_PN0P_  (.D(_02119_),
    .DE(_00070_),
    .Q(\w[57][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][30]$_SDFFCE_PN0P_  (.D(_02120_),
    .DE(_00070_),
    .Q(\w[57][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][31]$_SDFFCE_PN0P_  (.D(_02121_),
    .DE(_00070_),
    .Q(\w[57][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][3]$_SDFFCE_PN0P_  (.D(_02122_),
    .DE(_00070_),
    .Q(\w[57][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][4]$_SDFFCE_PN0P_  (.D(_02123_),
    .DE(_00070_),
    .Q(\w[57][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][5]$_SDFFCE_PN0P_  (.D(_02124_),
    .DE(_00070_),
    .Q(\w[57][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][6]$_SDFFCE_PN0P_  (.D(_02125_),
    .DE(_00070_),
    .Q(\w[57][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][7]$_SDFFCE_PN0P_  (.D(_02126_),
    .DE(_00070_),
    .Q(\w[57][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][8]$_SDFFCE_PN0P_  (.D(_02127_),
    .DE(_00070_),
    .Q(\w[57][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][9]$_SDFFCE_PN0P_  (.D(_02128_),
    .DE(_00070_),
    .Q(\w[57][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][0]$_SDFFCE_PN0P_  (.D(_02129_),
    .DE(_00100_),
    .Q(\w[58][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][10]$_SDFFCE_PN0P_  (.D(_02130_),
    .DE(_00100_),
    .Q(\w[58][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][11]$_SDFFCE_PN0P_  (.D(_02131_),
    .DE(_00100_),
    .Q(\w[58][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][12]$_SDFFCE_PN0P_  (.D(_02132_),
    .DE(_00100_),
    .Q(\w[58][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][13]$_SDFFCE_PN0P_  (.D(_02133_),
    .DE(_00100_),
    .Q(\w[58][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][14]$_SDFFCE_PN0P_  (.D(_02134_),
    .DE(_00100_),
    .Q(\w[58][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][15]$_SDFFCE_PN0P_  (.D(_02135_),
    .DE(_00100_),
    .Q(\w[58][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][16]$_SDFFCE_PN0P_  (.D(_02136_),
    .DE(_00100_),
    .Q(\w[58][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][17]$_SDFFCE_PN0P_  (.D(_02137_),
    .DE(_00100_),
    .Q(\w[58][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][18]$_SDFFCE_PN0P_  (.D(_02138_),
    .DE(_00100_),
    .Q(\w[58][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][19]$_SDFFCE_PN0P_  (.D(_02139_),
    .DE(_00100_),
    .Q(\w[58][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][1]$_SDFFCE_PN0P_  (.D(_02140_),
    .DE(_00100_),
    .Q(\w[58][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][20]$_SDFFCE_PN0P_  (.D(_02141_),
    .DE(_00100_),
    .Q(\w[58][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][21]$_SDFFCE_PN0P_  (.D(_02142_),
    .DE(_00100_),
    .Q(\w[58][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][22]$_SDFFCE_PN0P_  (.D(_02143_),
    .DE(_00100_),
    .Q(\w[58][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][23]$_SDFFCE_PN0P_  (.D(_02144_),
    .DE(_00100_),
    .Q(\w[58][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][24]$_SDFFCE_PN0P_  (.D(_02145_),
    .DE(_00100_),
    .Q(\w[58][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][25]$_SDFFCE_PN0P_  (.D(_02146_),
    .DE(_00100_),
    .Q(\w[58][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][26]$_SDFFCE_PN0P_  (.D(_02147_),
    .DE(_00100_),
    .Q(\w[58][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][27]$_SDFFCE_PN0P_  (.D(_02148_),
    .DE(_00100_),
    .Q(\w[58][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][28]$_SDFFCE_PN0P_  (.D(_02149_),
    .DE(_00100_),
    .Q(\w[58][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][29]$_SDFFCE_PN0P_  (.D(_02150_),
    .DE(_00100_),
    .Q(\w[58][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][2]$_SDFFCE_PN0P_  (.D(_02151_),
    .DE(_00100_),
    .Q(\w[58][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][30]$_SDFFCE_PN0P_  (.D(_02152_),
    .DE(_00100_),
    .Q(\w[58][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][31]$_SDFFCE_PN0P_  (.D(_02153_),
    .DE(_00100_),
    .Q(\w[58][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][3]$_SDFFCE_PN0P_  (.D(_02154_),
    .DE(_00100_),
    .Q(\w[58][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][4]$_SDFFCE_PN0P_  (.D(_02155_),
    .DE(_00100_),
    .Q(\w[58][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][5]$_SDFFCE_PN0P_  (.D(_02156_),
    .DE(_00100_),
    .Q(\w[58][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][6]$_SDFFCE_PN0P_  (.D(_02157_),
    .DE(_00100_),
    .Q(\w[58][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][7]$_SDFFCE_PN0P_  (.D(_02158_),
    .DE(_00100_),
    .Q(\w[58][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][8]$_SDFFCE_PN0P_  (.D(_02159_),
    .DE(_00100_),
    .Q(\w[58][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][9]$_SDFFCE_PN0P_  (.D(_02160_),
    .DE(_00100_),
    .Q(\w[58][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][0]$_SDFFCE_PN0P_  (.D(_02161_),
    .DE(_00069_),
    .Q(\w[59][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][10]$_SDFFCE_PN0P_  (.D(_02162_),
    .DE(_00069_),
    .Q(\w[59][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][11]$_SDFFCE_PN0P_  (.D(_02163_),
    .DE(_00069_),
    .Q(\w[59][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][12]$_SDFFCE_PN0P_  (.D(_02164_),
    .DE(_00069_),
    .Q(\w[59][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][13]$_SDFFCE_PN0P_  (.D(_02165_),
    .DE(_00069_),
    .Q(\w[59][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][14]$_SDFFCE_PN0P_  (.D(_02166_),
    .DE(_00069_),
    .Q(\w[59][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][15]$_SDFFCE_PN0P_  (.D(_02167_),
    .DE(_00069_),
    .Q(\w[59][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][16]$_SDFFCE_PN0P_  (.D(_02168_),
    .DE(_00069_),
    .Q(\w[59][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][17]$_SDFFCE_PN0P_  (.D(_02169_),
    .DE(_00069_),
    .Q(\w[59][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][18]$_SDFFCE_PN0P_  (.D(_02170_),
    .DE(_00069_),
    .Q(\w[59][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][19]$_SDFFCE_PN0P_  (.D(_02171_),
    .DE(_00069_),
    .Q(\w[59][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][1]$_SDFFCE_PN0P_  (.D(_02172_),
    .DE(_00069_),
    .Q(\w[59][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][20]$_SDFFCE_PN0P_  (.D(_02173_),
    .DE(_00069_),
    .Q(\w[59][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][21]$_SDFFCE_PN0P_  (.D(_02174_),
    .DE(_00069_),
    .Q(\w[59][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][22]$_SDFFCE_PN0P_  (.D(_02175_),
    .DE(_00069_),
    .Q(\w[59][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][23]$_SDFFCE_PN0P_  (.D(_02176_),
    .DE(_00069_),
    .Q(\w[59][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][24]$_SDFFCE_PN0P_  (.D(_02177_),
    .DE(_00069_),
    .Q(\w[59][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][25]$_SDFFCE_PN0P_  (.D(_02178_),
    .DE(_00069_),
    .Q(\w[59][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][26]$_SDFFCE_PN0P_  (.D(_02179_),
    .DE(_00069_),
    .Q(\w[59][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][27]$_SDFFCE_PN0P_  (.D(_02180_),
    .DE(_00069_),
    .Q(\w[59][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][28]$_SDFFCE_PN0P_  (.D(_02181_),
    .DE(_00069_),
    .Q(\w[59][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][29]$_SDFFCE_PN0P_  (.D(_02182_),
    .DE(_00069_),
    .Q(\w[59][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][2]$_SDFFCE_PN0P_  (.D(_02183_),
    .DE(_00069_),
    .Q(\w[59][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][30]$_SDFFCE_PN0P_  (.D(_02184_),
    .DE(_00069_),
    .Q(\w[59][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][31]$_SDFFCE_PN0P_  (.D(_02185_),
    .DE(_00069_),
    .Q(\w[59][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][3]$_SDFFCE_PN0P_  (.D(_02186_),
    .DE(_00069_),
    .Q(\w[59][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][4]$_SDFFCE_PN0P_  (.D(_02187_),
    .DE(_00069_),
    .Q(\w[59][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][5]$_SDFFCE_PN0P_  (.D(_02188_),
    .DE(_00069_),
    .Q(\w[59][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][6]$_SDFFCE_PN0P_  (.D(_02189_),
    .DE(_00069_),
    .Q(\w[59][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][7]$_SDFFCE_PN0P_  (.D(_02190_),
    .DE(_00069_),
    .Q(\w[59][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][8]$_SDFFCE_PN0P_  (.D(_02191_),
    .DE(_00069_),
    .Q(\w[59][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][9]$_SDFFCE_PN0P_  (.D(_02192_),
    .DE(_00069_),
    .Q(\w[59][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][0]$_DFFE_PP_  (.D(_00481_),
    .DE(_00068_),
    .Q(\w[5][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][10]$_DFFE_PP_  (.D(_00482_),
    .DE(_00068_),
    .Q(\w[5][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][11]$_DFFE_PP_  (.D(_00483_),
    .DE(_00068_),
    .Q(\w[5][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][12]$_DFFE_PP_  (.D(_00484_),
    .DE(_00068_),
    .Q(\w[5][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][13]$_DFFE_PP_  (.D(_00485_),
    .DE(_00068_),
    .Q(\w[5][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][14]$_DFFE_PP_  (.D(_00486_),
    .DE(_00068_),
    .Q(\w[5][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][15]$_DFFE_PP_  (.D(_00487_),
    .DE(_00068_),
    .Q(\w[5][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][16]$_DFFE_PP_  (.D(_00488_),
    .DE(_00068_),
    .Q(\w[5][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][17]$_DFFE_PP_  (.D(_00489_),
    .DE(_00068_),
    .Q(\w[5][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][18]$_DFFE_PP_  (.D(_00490_),
    .DE(_00068_),
    .Q(\w[5][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][19]$_DFFE_PP_  (.D(_00491_),
    .DE(_00068_),
    .Q(\w[5][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][1]$_DFFE_PP_  (.D(_00492_),
    .DE(_00068_),
    .Q(\w[5][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][20]$_DFFE_PP_  (.D(_00493_),
    .DE(_00068_),
    .Q(\w[5][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][21]$_DFFE_PP_  (.D(_00494_),
    .DE(_00068_),
    .Q(\w[5][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][22]$_DFFE_PP_  (.D(_00495_),
    .DE(_00068_),
    .Q(\w[5][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][23]$_DFFE_PP_  (.D(_00496_),
    .DE(_00068_),
    .Q(\w[5][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][24]$_DFFE_PP_  (.D(_00497_),
    .DE(_00068_),
    .Q(\w[5][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][25]$_DFFE_PP_  (.D(_00498_),
    .DE(_00068_),
    .Q(\w[5][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][26]$_DFFE_PP_  (.D(_00499_),
    .DE(_00068_),
    .Q(\w[5][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][27]$_DFFE_PP_  (.D(_00500_),
    .DE(_00068_),
    .Q(\w[5][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][28]$_DFFE_PP_  (.D(_00501_),
    .DE(_00068_),
    .Q(\w[5][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][29]$_DFFE_PP_  (.D(_00502_),
    .DE(_00068_),
    .Q(\w[5][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][2]$_DFFE_PP_  (.D(_00503_),
    .DE(_00068_),
    .Q(\w[5][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][30]$_DFFE_PP_  (.D(_00504_),
    .DE(_00068_),
    .Q(\w[5][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][31]$_DFFE_PP_  (.D(_00505_),
    .DE(_00068_),
    .Q(\w[5][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][3]$_DFFE_PP_  (.D(_00506_),
    .DE(_00068_),
    .Q(\w[5][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][4]$_DFFE_PP_  (.D(_00507_),
    .DE(_00068_),
    .Q(\w[5][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][5]$_DFFE_PP_  (.D(_00508_),
    .DE(_00068_),
    .Q(\w[5][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][6]$_DFFE_PP_  (.D(_00509_),
    .DE(_00068_),
    .Q(\w[5][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][7]$_DFFE_PP_  (.D(_00510_),
    .DE(_00068_),
    .Q(\w[5][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][8]$_DFFE_PP_  (.D(_00511_),
    .DE(_00068_),
    .Q(\w[5][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][9]$_DFFE_PP_  (.D(_00512_),
    .DE(_00068_),
    .Q(\w[5][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][0]$_SDFFCE_PN0P_  (.D(_02193_),
    .DE(_00099_),
    .Q(\w[60][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][10]$_SDFFCE_PN0P_  (.D(_02194_),
    .DE(_00099_),
    .Q(\w[60][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][11]$_SDFFCE_PN0P_  (.D(_02195_),
    .DE(_00099_),
    .Q(\w[60][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][12]$_SDFFCE_PN0P_  (.D(_02196_),
    .DE(_00099_),
    .Q(\w[60][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][13]$_SDFFCE_PN0P_  (.D(_02197_),
    .DE(_00099_),
    .Q(\w[60][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][14]$_SDFFCE_PN0P_  (.D(_02198_),
    .DE(_00099_),
    .Q(\w[60][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][15]$_SDFFCE_PN0P_  (.D(_02199_),
    .DE(_00099_),
    .Q(\w[60][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][16]$_SDFFCE_PN0P_  (.D(_02200_),
    .DE(_00099_),
    .Q(\w[60][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][17]$_SDFFCE_PN0P_  (.D(_02201_),
    .DE(_00099_),
    .Q(\w[60][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][18]$_SDFFCE_PN0P_  (.D(_02202_),
    .DE(_00099_),
    .Q(\w[60][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][19]$_SDFFCE_PN0P_  (.D(_02203_),
    .DE(_00099_),
    .Q(\w[60][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][1]$_SDFFCE_PN0P_  (.D(_02204_),
    .DE(_00099_),
    .Q(\w[60][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][20]$_SDFFCE_PN0P_  (.D(_02205_),
    .DE(_00099_),
    .Q(\w[60][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][21]$_SDFFCE_PN0P_  (.D(_02206_),
    .DE(_00099_),
    .Q(\w[60][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][22]$_SDFFCE_PN0P_  (.D(_02207_),
    .DE(_00099_),
    .Q(\w[60][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][23]$_SDFFCE_PN0P_  (.D(_02208_),
    .DE(_00099_),
    .Q(\w[60][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][24]$_SDFFCE_PN0P_  (.D(_02209_),
    .DE(_00099_),
    .Q(\w[60][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][25]$_SDFFCE_PN0P_  (.D(_02210_),
    .DE(_00099_),
    .Q(\w[60][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][26]$_SDFFCE_PN0P_  (.D(_02211_),
    .DE(_00099_),
    .Q(\w[60][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][27]$_SDFFCE_PN0P_  (.D(_02212_),
    .DE(_00099_),
    .Q(\w[60][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][28]$_SDFFCE_PN0P_  (.D(_02213_),
    .DE(_00099_),
    .Q(\w[60][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][29]$_SDFFCE_PN0P_  (.D(_02214_),
    .DE(_00099_),
    .Q(\w[60][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][2]$_SDFFCE_PN0P_  (.D(_02215_),
    .DE(_00099_),
    .Q(\w[60][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][30]$_SDFFCE_PN0P_  (.D(_02216_),
    .DE(_00099_),
    .Q(\w[60][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][31]$_SDFFCE_PN0P_  (.D(_02217_),
    .DE(_00099_),
    .Q(\w[60][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][3]$_SDFFCE_PN0P_  (.D(_02218_),
    .DE(_00099_),
    .Q(\w[60][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][4]$_SDFFCE_PN0P_  (.D(_02219_),
    .DE(_00099_),
    .Q(\w[60][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][5]$_SDFFCE_PN0P_  (.D(_02220_),
    .DE(_00099_),
    .Q(\w[60][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][6]$_SDFFCE_PN0P_  (.D(_02221_),
    .DE(_00099_),
    .Q(\w[60][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][7]$_SDFFCE_PN0P_  (.D(_02222_),
    .DE(_00099_),
    .Q(\w[60][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][8]$_SDFFCE_PN0P_  (.D(_02223_),
    .DE(_00099_),
    .Q(\w[60][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][9]$_SDFFCE_PN0P_  (.D(_02224_),
    .DE(_00099_),
    .Q(\w[60][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][0]$_SDFFCE_PN0P_  (.D(_02225_),
    .DE(_00067_),
    .Q(\w[61][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][10]$_SDFFCE_PN0P_  (.D(_02226_),
    .DE(_00067_),
    .Q(\w[61][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][11]$_SDFFCE_PN0P_  (.D(_02227_),
    .DE(_00067_),
    .Q(\w[61][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][12]$_SDFFCE_PN0P_  (.D(_02228_),
    .DE(_00067_),
    .Q(\w[61][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][13]$_SDFFCE_PN0P_  (.D(_02229_),
    .DE(_00067_),
    .Q(\w[61][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][14]$_SDFFCE_PN0P_  (.D(_02230_),
    .DE(_00067_),
    .Q(\w[61][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][15]$_SDFFCE_PN0P_  (.D(_02231_),
    .DE(_00067_),
    .Q(\w[61][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][16]$_SDFFCE_PN0P_  (.D(_02232_),
    .DE(_00067_),
    .Q(\w[61][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][17]$_SDFFCE_PN0P_  (.D(_02233_),
    .DE(_00067_),
    .Q(\w[61][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][18]$_SDFFCE_PN0P_  (.D(_02234_),
    .DE(_00067_),
    .Q(\w[61][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][19]$_SDFFCE_PN0P_  (.D(_02235_),
    .DE(_00067_),
    .Q(\w[61][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][1]$_SDFFCE_PN0P_  (.D(_02236_),
    .DE(_00067_),
    .Q(\w[61][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][20]$_SDFFCE_PN0P_  (.D(_02237_),
    .DE(_00067_),
    .Q(\w[61][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][21]$_SDFFCE_PN0P_  (.D(_02238_),
    .DE(_00067_),
    .Q(\w[61][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][22]$_SDFFCE_PN0P_  (.D(_02239_),
    .DE(_00067_),
    .Q(\w[61][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][23]$_SDFFCE_PN0P_  (.D(_02240_),
    .DE(_00067_),
    .Q(\w[61][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][24]$_SDFFCE_PN0P_  (.D(_02241_),
    .DE(_00067_),
    .Q(\w[61][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][25]$_SDFFCE_PN0P_  (.D(_02242_),
    .DE(_00067_),
    .Q(\w[61][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][26]$_SDFFCE_PN0P_  (.D(_02243_),
    .DE(_00067_),
    .Q(\w[61][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][27]$_SDFFCE_PN0P_  (.D(_02244_),
    .DE(_00067_),
    .Q(\w[61][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][28]$_SDFFCE_PN0P_  (.D(_02245_),
    .DE(_00067_),
    .Q(\w[61][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][29]$_SDFFCE_PN0P_  (.D(_02246_),
    .DE(_00067_),
    .Q(\w[61][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][2]$_SDFFCE_PN0P_  (.D(_02247_),
    .DE(_00067_),
    .Q(\w[61][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][30]$_SDFFCE_PN0P_  (.D(_02248_),
    .DE(_00067_),
    .Q(\w[61][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][31]$_SDFFCE_PN0P_  (.D(_02249_),
    .DE(_00067_),
    .Q(\w[61][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][3]$_SDFFCE_PN0P_  (.D(_02250_),
    .DE(_00067_),
    .Q(\w[61][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][4]$_SDFFCE_PN0P_  (.D(_02251_),
    .DE(_00067_),
    .Q(\w[61][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][5]$_SDFFCE_PN0P_  (.D(_02252_),
    .DE(_00067_),
    .Q(\w[61][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][6]$_SDFFCE_PN0P_  (.D(_02253_),
    .DE(_00067_),
    .Q(\w[61][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][7]$_SDFFCE_PN0P_  (.D(_02254_),
    .DE(_00067_),
    .Q(\w[61][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][8]$_SDFFCE_PN0P_  (.D(_02255_),
    .DE(_00067_),
    .Q(\w[61][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][9]$_SDFFCE_PN0P_  (.D(_02256_),
    .DE(_00067_),
    .Q(\w[61][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][0]$_SDFFCE_PN0P_  (.D(_02257_),
    .DE(_00098_),
    .Q(\w[62][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][10]$_SDFFCE_PN0P_  (.D(_02258_),
    .DE(_00098_),
    .Q(\w[62][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][11]$_SDFFCE_PN0P_  (.D(_02259_),
    .DE(_00098_),
    .Q(\w[62][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][12]$_SDFFCE_PN0P_  (.D(_02260_),
    .DE(_00098_),
    .Q(\w[62][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][13]$_SDFFCE_PN0P_  (.D(_02261_),
    .DE(_00098_),
    .Q(\w[62][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][14]$_SDFFCE_PN0P_  (.D(_02262_),
    .DE(_00098_),
    .Q(\w[62][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][15]$_SDFFCE_PN0P_  (.D(_02263_),
    .DE(_00098_),
    .Q(\w[62][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][16]$_SDFFCE_PN0P_  (.D(_02264_),
    .DE(_00098_),
    .Q(\w[62][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][17]$_SDFFCE_PN0P_  (.D(_02265_),
    .DE(_00098_),
    .Q(\w[62][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][18]$_SDFFCE_PN0P_  (.D(_02266_),
    .DE(_00098_),
    .Q(\w[62][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][19]$_SDFFCE_PN0P_  (.D(_02267_),
    .DE(_00098_),
    .Q(\w[62][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][1]$_SDFFCE_PN0P_  (.D(_02268_),
    .DE(_00098_),
    .Q(\w[62][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][20]$_SDFFCE_PN0P_  (.D(_02269_),
    .DE(_00098_),
    .Q(\w[62][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][21]$_SDFFCE_PN0P_  (.D(_02270_),
    .DE(_00098_),
    .Q(\w[62][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][22]$_SDFFCE_PN0P_  (.D(_02271_),
    .DE(_00098_),
    .Q(\w[62][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][23]$_SDFFCE_PN0P_  (.D(_02272_),
    .DE(_00098_),
    .Q(\w[62][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][24]$_SDFFCE_PN0P_  (.D(_02273_),
    .DE(_00098_),
    .Q(\w[62][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][25]$_SDFFCE_PN0P_  (.D(_02274_),
    .DE(_00098_),
    .Q(\w[62][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][26]$_SDFFCE_PN0P_  (.D(_02275_),
    .DE(_00098_),
    .Q(\w[62][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][27]$_SDFFCE_PN0P_  (.D(_02276_),
    .DE(_00098_),
    .Q(\w[62][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][28]$_SDFFCE_PN0P_  (.D(_02277_),
    .DE(_00098_),
    .Q(\w[62][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][29]$_SDFFCE_PN0P_  (.D(_02278_),
    .DE(_00098_),
    .Q(\w[62][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][2]$_SDFFCE_PN0P_  (.D(_02279_),
    .DE(_00098_),
    .Q(\w[62][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][30]$_SDFFCE_PN0P_  (.D(_02280_),
    .DE(_00098_),
    .Q(\w[62][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][31]$_SDFFCE_PN0P_  (.D(_02281_),
    .DE(_00098_),
    .Q(\w[62][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][3]$_SDFFCE_PN0P_  (.D(_02282_),
    .DE(_00098_),
    .Q(\w[62][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][4]$_SDFFCE_PN0P_  (.D(_02283_),
    .DE(_00098_),
    .Q(\w[62][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][5]$_SDFFCE_PN0P_  (.D(_02284_),
    .DE(_00098_),
    .Q(\w[62][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][6]$_SDFFCE_PN0P_  (.D(_02285_),
    .DE(_00098_),
    .Q(\w[62][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][7]$_SDFFCE_PN0P_  (.D(_02286_),
    .DE(_00098_),
    .Q(\w[62][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][8]$_SDFFCE_PN0P_  (.D(_02287_),
    .DE(_00098_),
    .Q(\w[62][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][9]$_SDFFCE_PN0P_  (.D(_02288_),
    .DE(_00098_),
    .Q(\w[62][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][0]$_SDFFCE_PN0P_  (.D(_02289_),
    .DE(_00066_),
    .Q(\w[63][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][10]$_SDFFCE_PN0P_  (.D(_02290_),
    .DE(_00066_),
    .Q(\w[63][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][11]$_SDFFCE_PN0P_  (.D(_02291_),
    .DE(_00066_),
    .Q(\w[63][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][12]$_SDFFCE_PN0P_  (.D(_02292_),
    .DE(_00066_),
    .Q(\w[63][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][13]$_SDFFCE_PN0P_  (.D(_02293_),
    .DE(_00066_),
    .Q(\w[63][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][14]$_SDFFCE_PN0P_  (.D(_02294_),
    .DE(_00066_),
    .Q(\w[63][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][15]$_SDFFCE_PN0P_  (.D(_02295_),
    .DE(_00066_),
    .Q(\w[63][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][16]$_SDFFCE_PN0P_  (.D(_02296_),
    .DE(_00066_),
    .Q(\w[63][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][17]$_SDFFCE_PN0P_  (.D(_02297_),
    .DE(_00066_),
    .Q(\w[63][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][18]$_SDFFCE_PN0P_  (.D(_02298_),
    .DE(_00066_),
    .Q(\w[63][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][19]$_SDFFCE_PN0P_  (.D(_02299_),
    .DE(_00066_),
    .Q(\w[63][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][1]$_SDFFCE_PN0P_  (.D(_02300_),
    .DE(_00066_),
    .Q(\w[63][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][20]$_SDFFCE_PN0P_  (.D(_02301_),
    .DE(_00066_),
    .Q(\w[63][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][21]$_SDFFCE_PN0P_  (.D(_02302_),
    .DE(_00066_),
    .Q(\w[63][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][22]$_SDFFCE_PN0P_  (.D(_02303_),
    .DE(_00066_),
    .Q(\w[63][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][23]$_SDFFCE_PN0P_  (.D(_02304_),
    .DE(_00066_),
    .Q(\w[63][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][24]$_SDFFCE_PN0P_  (.D(_02305_),
    .DE(_00066_),
    .Q(\w[63][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][25]$_SDFFCE_PN0P_  (.D(_02306_),
    .DE(_00066_),
    .Q(\w[63][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][26]$_SDFFCE_PN0P_  (.D(_02307_),
    .DE(_00066_),
    .Q(\w[63][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][27]$_SDFFCE_PN0P_  (.D(_02308_),
    .DE(_00066_),
    .Q(\w[63][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][28]$_SDFFCE_PN0P_  (.D(_02309_),
    .DE(_00066_),
    .Q(\w[63][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][29]$_SDFFCE_PN0P_  (.D(_02310_),
    .DE(_00066_),
    .Q(\w[63][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][2]$_SDFFCE_PN0P_  (.D(_02311_),
    .DE(_00066_),
    .Q(\w[63][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][30]$_SDFFCE_PN0P_  (.D(_02312_),
    .DE(_00066_),
    .Q(\w[63][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][31]$_SDFFCE_PN0P_  (.D(_02313_),
    .DE(_00066_),
    .Q(\w[63][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][3]$_SDFFCE_PN0P_  (.D(_02314_),
    .DE(_00066_),
    .Q(\w[63][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][4]$_SDFFCE_PN0P_  (.D(_02315_),
    .DE(_00066_),
    .Q(\w[63][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][5]$_SDFFCE_PN0P_  (.D(_02316_),
    .DE(_00066_),
    .Q(\w[63][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][6]$_SDFFCE_PN0P_  (.D(_02317_),
    .DE(_00066_),
    .Q(\w[63][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][7]$_SDFFCE_PN0P_  (.D(_02318_),
    .DE(_00066_),
    .Q(\w[63][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][8]$_SDFFCE_PN0P_  (.D(_02319_),
    .DE(_00066_),
    .Q(\w[63][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][9]$_SDFFCE_PN0P_  (.D(_02320_),
    .DE(_00066_),
    .Q(\w[63][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][0]$_DFFE_PP_  (.D(_00513_),
    .DE(_00097_),
    .Q(\w[6][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][10]$_DFFE_PP_  (.D(_00514_),
    .DE(_00097_),
    .Q(\w[6][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][11]$_DFFE_PP_  (.D(_00515_),
    .DE(_00097_),
    .Q(\w[6][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][12]$_DFFE_PP_  (.D(_00516_),
    .DE(_00097_),
    .Q(\w[6][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][13]$_DFFE_PP_  (.D(_00517_),
    .DE(_00097_),
    .Q(\w[6][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][14]$_DFFE_PP_  (.D(_00518_),
    .DE(_00097_),
    .Q(\w[6][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][15]$_DFFE_PP_  (.D(_00519_),
    .DE(_00097_),
    .Q(\w[6][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][16]$_DFFE_PP_  (.D(_00520_),
    .DE(_00097_),
    .Q(\w[6][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][17]$_DFFE_PP_  (.D(_00521_),
    .DE(_00097_),
    .Q(\w[6][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][18]$_DFFE_PP_  (.D(_00522_),
    .DE(_00097_),
    .Q(\w[6][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][19]$_DFFE_PP_  (.D(_00523_),
    .DE(_00097_),
    .Q(\w[6][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][1]$_DFFE_PP_  (.D(_00524_),
    .DE(_00097_),
    .Q(\w[6][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][20]$_DFFE_PP_  (.D(_00525_),
    .DE(_00097_),
    .Q(\w[6][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][21]$_DFFE_PP_  (.D(_00526_),
    .DE(_00097_),
    .Q(\w[6][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][22]$_DFFE_PP_  (.D(_00527_),
    .DE(_00097_),
    .Q(\w[6][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][23]$_DFFE_PP_  (.D(_00528_),
    .DE(_00097_),
    .Q(\w[6][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][24]$_DFFE_PP_  (.D(_00529_),
    .DE(_00097_),
    .Q(\w[6][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][25]$_DFFE_PP_  (.D(_00530_),
    .DE(_00097_),
    .Q(\w[6][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][26]$_DFFE_PP_  (.D(_00531_),
    .DE(_00097_),
    .Q(\w[6][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][27]$_DFFE_PP_  (.D(_00532_),
    .DE(_00097_),
    .Q(\w[6][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][28]$_DFFE_PP_  (.D(_00533_),
    .DE(_00097_),
    .Q(\w[6][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][29]$_DFFE_PP_  (.D(_00534_),
    .DE(_00097_),
    .Q(\w[6][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][2]$_DFFE_PP_  (.D(_00535_),
    .DE(_00097_),
    .Q(\w[6][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][30]$_DFFE_PP_  (.D(_00536_),
    .DE(_00097_),
    .Q(\w[6][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][31]$_DFFE_PP_  (.D(_00537_),
    .DE(_00097_),
    .Q(\w[6][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][3]$_DFFE_PP_  (.D(_00538_),
    .DE(_00097_),
    .Q(\w[6][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][4]$_DFFE_PP_  (.D(_00539_),
    .DE(_00097_),
    .Q(\w[6][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][5]$_DFFE_PP_  (.D(_00540_),
    .DE(_00097_),
    .Q(\w[6][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][6]$_DFFE_PP_  (.D(_00541_),
    .DE(_00097_),
    .Q(\w[6][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][7]$_DFFE_PP_  (.D(_00542_),
    .DE(_00097_),
    .Q(\w[6][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][8]$_DFFE_PP_  (.D(_00543_),
    .DE(_00097_),
    .Q(\w[6][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][9]$_DFFE_PP_  (.D(_00544_),
    .DE(_00097_),
    .Q(\w[6][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][0]$_DFFE_PP_  (.D(_00545_),
    .DE(_00065_),
    .Q(\w[7][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][10]$_DFFE_PP_  (.D(_00546_),
    .DE(_00065_),
    .Q(\w[7][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][11]$_DFFE_PP_  (.D(_00547_),
    .DE(_00065_),
    .Q(\w[7][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][12]$_DFFE_PP_  (.D(_00548_),
    .DE(_00065_),
    .Q(\w[7][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][13]$_DFFE_PP_  (.D(_00549_),
    .DE(_00065_),
    .Q(\w[7][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][14]$_DFFE_PP_  (.D(_00550_),
    .DE(_00065_),
    .Q(\w[7][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][15]$_DFFE_PP_  (.D(_00551_),
    .DE(_00065_),
    .Q(\w[7][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][16]$_DFFE_PP_  (.D(_00552_),
    .DE(_00065_),
    .Q(\w[7][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][17]$_DFFE_PP_  (.D(_00553_),
    .DE(_00065_),
    .Q(\w[7][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][18]$_DFFE_PP_  (.D(_00554_),
    .DE(_00065_),
    .Q(\w[7][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][19]$_DFFE_PP_  (.D(_00555_),
    .DE(_00065_),
    .Q(\w[7][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][1]$_DFFE_PP_  (.D(_00556_),
    .DE(_00065_),
    .Q(\w[7][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][20]$_DFFE_PP_  (.D(_00557_),
    .DE(_00065_),
    .Q(\w[7][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][21]$_DFFE_PP_  (.D(_00558_),
    .DE(_00065_),
    .Q(\w[7][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][22]$_DFFE_PP_  (.D(_00559_),
    .DE(_00065_),
    .Q(\w[7][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][23]$_DFFE_PP_  (.D(_00560_),
    .DE(_00065_),
    .Q(\w[7][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][24]$_DFFE_PP_  (.D(_00561_),
    .DE(_00065_),
    .Q(\w[7][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][25]$_DFFE_PP_  (.D(_00562_),
    .DE(_00065_),
    .Q(\w[7][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][26]$_DFFE_PP_  (.D(_00563_),
    .DE(_00065_),
    .Q(\w[7][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][27]$_DFFE_PP_  (.D(_00564_),
    .DE(_00065_),
    .Q(\w[7][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][28]$_DFFE_PP_  (.D(_00565_),
    .DE(_00065_),
    .Q(\w[7][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][29]$_DFFE_PP_  (.D(_00566_),
    .DE(_00065_),
    .Q(\w[7][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][2]$_DFFE_PP_  (.D(_00567_),
    .DE(_00065_),
    .Q(\w[7][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][30]$_DFFE_PP_  (.D(_00568_),
    .DE(_00065_),
    .Q(\w[7][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][31]$_DFFE_PP_  (.D(_00569_),
    .DE(_00065_),
    .Q(\w[7][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][3]$_DFFE_PP_  (.D(_00570_),
    .DE(_00065_),
    .Q(\w[7][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][4]$_DFFE_PP_  (.D(_00571_),
    .DE(_00065_),
    .Q(\w[7][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][5]$_DFFE_PP_  (.D(_00572_),
    .DE(_00065_),
    .Q(\w[7][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][6]$_DFFE_PP_  (.D(_00573_),
    .DE(_00065_),
    .Q(\w[7][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][7]$_DFFE_PP_  (.D(_00574_),
    .DE(_00065_),
    .Q(\w[7][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][8]$_DFFE_PP_  (.D(_00575_),
    .DE(_00065_),
    .Q(\w[7][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][9]$_DFFE_PP_  (.D(_00576_),
    .DE(_00065_),
    .Q(\w[7][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][0]$_DFFE_PP_  (.D(_00577_),
    .DE(_00096_),
    .Q(\w[8][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][10]$_DFFE_PP_  (.D(_00578_),
    .DE(_00096_),
    .Q(\w[8][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][11]$_DFFE_PP_  (.D(_00579_),
    .DE(_00096_),
    .Q(\w[8][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][12]$_DFFE_PP_  (.D(_00580_),
    .DE(_00096_),
    .Q(\w[8][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][13]$_DFFE_PP_  (.D(_00581_),
    .DE(_00096_),
    .Q(\w[8][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][14]$_DFFE_PP_  (.D(_00582_),
    .DE(_00096_),
    .Q(\w[8][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][15]$_DFFE_PP_  (.D(_00583_),
    .DE(_00096_),
    .Q(\w[8][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][16]$_DFFE_PP_  (.D(_00584_),
    .DE(_00096_),
    .Q(\w[8][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][17]$_DFFE_PP_  (.D(_00585_),
    .DE(_00096_),
    .Q(\w[8][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][18]$_DFFE_PP_  (.D(_00586_),
    .DE(_00096_),
    .Q(\w[8][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][19]$_DFFE_PP_  (.D(_00587_),
    .DE(_00096_),
    .Q(\w[8][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][1]$_DFFE_PP_  (.D(_00588_),
    .DE(_00096_),
    .Q(\w[8][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][20]$_DFFE_PP_  (.D(_00589_),
    .DE(_00096_),
    .Q(\w[8][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][21]$_DFFE_PP_  (.D(_00590_),
    .DE(_00096_),
    .Q(\w[8][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][22]$_DFFE_PP_  (.D(_00591_),
    .DE(_00096_),
    .Q(\w[8][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][23]$_DFFE_PP_  (.D(_00592_),
    .DE(_00096_),
    .Q(\w[8][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][24]$_DFFE_PP_  (.D(_00593_),
    .DE(_00096_),
    .Q(\w[8][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][25]$_DFFE_PP_  (.D(_00594_),
    .DE(_00096_),
    .Q(\w[8][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][26]$_DFFE_PP_  (.D(_00595_),
    .DE(_00096_),
    .Q(\w[8][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][27]$_DFFE_PP_  (.D(_00596_),
    .DE(_00096_),
    .Q(\w[8][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][28]$_DFFE_PP_  (.D(_00597_),
    .DE(_00096_),
    .Q(\w[8][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][29]$_DFFE_PP_  (.D(_00598_),
    .DE(_00096_),
    .Q(\w[8][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][2]$_DFFE_PP_  (.D(_00599_),
    .DE(_00096_),
    .Q(\w[8][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][30]$_DFFE_PP_  (.D(_00600_),
    .DE(_00096_),
    .Q(\w[8][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][31]$_DFFE_PP_  (.D(_00601_),
    .DE(_00096_),
    .Q(\w[8][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][3]$_DFFE_PP_  (.D(_00602_),
    .DE(_00096_),
    .Q(\w[8][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][4]$_DFFE_PP_  (.D(_00603_),
    .DE(_00096_),
    .Q(\w[8][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][5]$_DFFE_PP_  (.D(_00604_),
    .DE(_00096_),
    .Q(\w[8][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][6]$_DFFE_PP_  (.D(_00605_),
    .DE(_00096_),
    .Q(\w[8][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][7]$_DFFE_PP_  (.D(_00606_),
    .DE(_00096_),
    .Q(\w[8][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][8]$_DFFE_PP_  (.D(_00607_),
    .DE(_00096_),
    .Q(\w[8][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][9]$_DFFE_PP_  (.D(_00608_),
    .DE(_00096_),
    .Q(\w[8][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][0]$_DFFE_PP_  (.D(_00609_),
    .DE(_00064_),
    .Q(\w[9][0] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][10]$_DFFE_PP_  (.D(_00610_),
    .DE(_00064_),
    .Q(\w[9][10] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][11]$_DFFE_PP_  (.D(_00611_),
    .DE(_00064_),
    .Q(\w[9][11] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][12]$_DFFE_PP_  (.D(_00612_),
    .DE(_00064_),
    .Q(\w[9][12] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][13]$_DFFE_PP_  (.D(_00613_),
    .DE(_00064_),
    .Q(\w[9][13] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][14]$_DFFE_PP_  (.D(_00614_),
    .DE(_00064_),
    .Q(\w[9][14] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][15]$_DFFE_PP_  (.D(_00615_),
    .DE(_00064_),
    .Q(\w[9][15] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][16]$_DFFE_PP_  (.D(_00616_),
    .DE(_00064_),
    .Q(\w[9][16] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][17]$_DFFE_PP_  (.D(_00617_),
    .DE(_00064_),
    .Q(\w[9][17] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][18]$_DFFE_PP_  (.D(_00618_),
    .DE(_00064_),
    .Q(\w[9][18] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][19]$_DFFE_PP_  (.D(_00619_),
    .DE(_00064_),
    .Q(\w[9][19] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][1]$_DFFE_PP_  (.D(_00620_),
    .DE(_00064_),
    .Q(\w[9][1] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][20]$_DFFE_PP_  (.D(_00621_),
    .DE(_00064_),
    .Q(\w[9][20] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][21]$_DFFE_PP_  (.D(_00622_),
    .DE(_00064_),
    .Q(\w[9][21] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][22]$_DFFE_PP_  (.D(_00623_),
    .DE(_00064_),
    .Q(\w[9][22] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][23]$_DFFE_PP_  (.D(_00624_),
    .DE(_00064_),
    .Q(\w[9][23] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][24]$_DFFE_PP_  (.D(_00625_),
    .DE(_00064_),
    .Q(\w[9][24] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][25]$_DFFE_PP_  (.D(_00626_),
    .DE(_00064_),
    .Q(\w[9][25] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][26]$_DFFE_PP_  (.D(_00627_),
    .DE(_00064_),
    .Q(\w[9][26] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][27]$_DFFE_PP_  (.D(_00628_),
    .DE(_00064_),
    .Q(\w[9][27] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][28]$_DFFE_PP_  (.D(_00629_),
    .DE(_00064_),
    .Q(\w[9][28] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][29]$_DFFE_PP_  (.D(_00630_),
    .DE(_00064_),
    .Q(\w[9][29] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][2]$_DFFE_PP_  (.D(_00631_),
    .DE(_00064_),
    .Q(\w[9][2] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][30]$_DFFE_PP_  (.D(_00632_),
    .DE(_00064_),
    .Q(\w[9][30] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][31]$_DFFE_PP_  (.D(_00633_),
    .DE(_00064_),
    .Q(\w[9][31] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][3]$_DFFE_PP_  (.D(_00634_),
    .DE(_00064_),
    .Q(\w[9][3] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][4]$_DFFE_PP_  (.D(_00635_),
    .DE(_00064_),
    .Q(\w[9][4] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][5]$_DFFE_PP_  (.D(_00636_),
    .DE(_00064_),
    .Q(\w[9][5] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][6]$_DFFE_PP_  (.D(_00637_),
    .DE(_00064_),
    .Q(\w[9][6] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][7]$_DFFE_PP_  (.D(_00638_),
    .DE(_00064_),
    .Q(\w[9][7] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][8]$_DFFE_PP_  (.D(_00639_),
    .DE(_00064_),
    .Q(\w[9][8] ),
    .CLK(clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][9]$_DFFE_PP_  (.D(_00640_),
    .DE(_00064_),
    .Q(\w[9][9] ),
    .CLK(clk));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_00_  (.A(\w_new_calc1.w_15[18] ),
    .B(\w_new_calc1.w_15[7] ),
    .C(\w_new_calc1.w_15[3] ),
    .X(\w_new_calc1.temp1[0] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_01_  (.A(\w_new_calc1.w_15[13] ),
    .B(\w_new_calc1.w_15[28] ),
    .C(\w_new_calc1.w_15[17] ),
    .X(\w_new_calc1.temp1[10] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_02_  (.A(\w_new_calc1.w_15[18] ),
    .B(\w_new_calc1.w_15[14] ),
    .C(\w_new_calc1.w_15[29] ),
    .X(\w_new_calc1.temp1[11] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_03_  (.A(\w_new_calc1.w_15[19] ),
    .B(\w_new_calc1.w_15[15] ),
    .C(\w_new_calc1.w_15[30] ),
    .X(\w_new_calc1.temp1[12] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_04_  (.A(\w_new_calc1.w_15[20] ),
    .B(\w_new_calc1.w_15[16] ),
    .C(\w_new_calc1.w_15[31] ),
    .X(\w_new_calc1.temp1[13] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_05_  (.A(\w_new_calc1.w_15[21] ),
    .B(\w_new_calc1.w_15[17] ),
    .C(\w_new_calc1.w_15[0] ),
    .X(\w_new_calc1.temp1[14] ));
 sky130_fd_sc_hd__xor3_4 \w_new_calc1.s0/_06_  (.A(\w_new_calc1.w_15[18] ),
    .B(\w_new_calc1.w_15[22] ),
    .C(\w_new_calc1.w_15[1] ),
    .X(\w_new_calc1.temp1[15] ));
 sky130_fd_sc_hd__xor3_4 \w_new_calc1.s0/_07_  (.A(\w_new_calc1.w_15[19] ),
    .B(\w_new_calc1.w_15[23] ),
    .C(\w_new_calc1.w_15[2] ),
    .X(\w_new_calc1.temp1[16] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_08_  (.A(\w_new_calc1.w_15[20] ),
    .B(\w_new_calc1.w_15[24] ),
    .C(\w_new_calc1.w_15[3] ),
    .X(\w_new_calc1.temp1[17] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_09_  (.A(\w_new_calc1.w_15[21] ),
    .B(\w_new_calc1.w_15[25] ),
    .C(\w_new_calc1.w_15[4] ),
    .X(\w_new_calc1.temp1[18] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_10_  (.A(\w_new_calc1.w_15[22] ),
    .B(\w_new_calc1.w_15[26] ),
    .C(\w_new_calc1.w_15[5] ),
    .X(\w_new_calc1.temp1[19] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_11_  (.A(\w_new_calc1.w_15[19] ),
    .B(\w_new_calc1.w_15[8] ),
    .C(\w_new_calc1.w_15[4] ),
    .X(\w_new_calc1.temp1[1] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_12_  (.A(\w_new_calc1.w_15[23] ),
    .B(\w_new_calc1.w_15[27] ),
    .C(\w_new_calc1.w_15[6] ),
    .X(\w_new_calc1.temp1[20] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_13_  (.A(\w_new_calc1.w_15[7] ),
    .B(\w_new_calc1.w_15[24] ),
    .C(\w_new_calc1.w_15[28] ),
    .X(\w_new_calc1.temp1[21] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_14_  (.A(\w_new_calc1.w_15[8] ),
    .B(\w_new_calc1.w_15[25] ),
    .C(\w_new_calc1.w_15[29] ),
    .X(\w_new_calc1.temp1[22] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_15_  (.A(\w_new_calc1.w_15[9] ),
    .B(\w_new_calc1.w_15[26] ),
    .C(\w_new_calc1.w_15[30] ),
    .X(\w_new_calc1.temp1[23] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_16_  (.A(\w_new_calc1.w_15[10] ),
    .B(\w_new_calc1.w_15[27] ),
    .C(\w_new_calc1.w_15[31] ),
    .X(\w_new_calc1.temp1[24] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_17_  (.A(\w_new_calc1.w_15[11] ),
    .B(\w_new_calc1.w_15[28] ),
    .C(\w_new_calc1.w_15[0] ),
    .X(\w_new_calc1.temp1[25] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_18_  (.A(\w_new_calc1.w_15[12] ),
    .B(\w_new_calc1.w_15[29] ),
    .C(\w_new_calc1.w_15[1] ),
    .X(\w_new_calc1.temp1[26] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_19_  (.A(\w_new_calc1.w_15[13] ),
    .B(\w_new_calc1.w_15[30] ),
    .C(\w_new_calc1.w_15[2] ),
    .X(\w_new_calc1.temp1[27] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_20_  (.A(\w_new_calc1.w_15[14] ),
    .B(\w_new_calc1.w_15[31] ),
    .C(\w_new_calc1.w_15[3] ),
    .X(\w_new_calc1.temp1[28] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s0/_21_  (.A(\w_new_calc1.w_15[15] ),
    .B(\w_new_calc1.w_15[4] ),
    .X(\w_new_calc1.temp1[29] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_22_  (.A(\w_new_calc1.w_15[20] ),
    .B(\w_new_calc1.w_15[9] ),
    .C(\w_new_calc1.w_15[5] ),
    .X(\w_new_calc1.temp1[2] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s0/_23_  (.A(\w_new_calc1.w_15[16] ),
    .B(\w_new_calc1.w_15[5] ),
    .X(\w_new_calc1.temp1[30] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s0/_24_  (.A(\w_new_calc1.w_15[17] ),
    .B(\w_new_calc1.w_15[6] ),
    .X(\w_new_calc1.temp1[31] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_25_  (.A(\w_new_calc1.w_15[21] ),
    .B(\w_new_calc1.w_15[10] ),
    .C(\w_new_calc1.w_15[6] ),
    .X(\w_new_calc1.temp1[3] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_26_  (.A(\w_new_calc1.w_15[7] ),
    .B(\w_new_calc1.w_15[22] ),
    .C(\w_new_calc1.w_15[11] ),
    .X(\w_new_calc1.temp1[4] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_27_  (.A(\w_new_calc1.w_15[8] ),
    .B(\w_new_calc1.w_15[23] ),
    .C(\w_new_calc1.w_15[12] ),
    .X(\w_new_calc1.temp1[5] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_28_  (.A(\w_new_calc1.w_15[9] ),
    .B(\w_new_calc1.w_15[24] ),
    .C(\w_new_calc1.w_15[13] ),
    .X(\w_new_calc1.temp1[6] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_29_  (.A(\w_new_calc1.w_15[10] ),
    .B(\w_new_calc1.w_15[25] ),
    .C(\w_new_calc1.w_15[14] ),
    .X(\w_new_calc1.temp1[7] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_30_  (.A(\w_new_calc1.w_15[11] ),
    .B(\w_new_calc1.w_15[26] ),
    .C(\w_new_calc1.w_15[15] ),
    .X(\w_new_calc1.temp1[8] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s0/_31_  (.A(\w_new_calc1.w_15[12] ),
    .B(\w_new_calc1.w_15[27] ),
    .C(\w_new_calc1.w_15[16] ),
    .X(\w_new_calc1.temp1[9] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_00_  (.A(\w_new_calc1.w_2[19] ),
    .B(\w_new_calc1.w_2[17] ),
    .C(\w_new_calc1.w_2[10] ),
    .X(\w_new_calc1.temp2[0] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_01_  (.A(\w_new_calc1.w_2[20] ),
    .B(\w_new_calc1.w_2[27] ),
    .C(\w_new_calc1.w_2[29] ),
    .X(\w_new_calc1.temp2[10] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_02_  (.A(\w_new_calc1.w_2[21] ),
    .B(\w_new_calc1.w_2[28] ),
    .C(\w_new_calc1.w_2[30] ),
    .X(\w_new_calc1.temp2[11] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_03_  (.A(\w_new_calc1.w_2[22] ),
    .B(\w_new_calc1.w_2[29] ),
    .C(\w_new_calc1.w_2[31] ),
    .X(\w_new_calc1.temp2[12] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_04_  (.A(\w_new_calc1.w_2[23] ),
    .B(\w_new_calc1.w_2[30] ),
    .C(\w_new_calc1.w_2[0] ),
    .X(\w_new_calc1.temp2[13] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_05_  (.A(\w_new_calc1.w_2[24] ),
    .B(\w_new_calc1.w_2[31] ),
    .C(\w_new_calc1.w_2[1] ),
    .X(\w_new_calc1.temp2[14] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_06_  (.A(\w_new_calc1.w_2[25] ),
    .B(\w_new_calc1.w_2[0] ),
    .C(\w_new_calc1.w_2[2] ),
    .X(\w_new_calc1.temp2[15] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_07_  (.A(\w_new_calc1.w_2[26] ),
    .B(\w_new_calc1.w_2[1] ),
    .C(\w_new_calc1.w_2[3] ),
    .X(\w_new_calc1.temp2[16] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_08_  (.A(\w_new_calc1.w_2[27] ),
    .B(\w_new_calc1.w_2[2] ),
    .C(\w_new_calc1.w_2[4] ),
    .X(\w_new_calc1.temp2[17] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_09_  (.A(\w_new_calc1.w_2[28] ),
    .B(\w_new_calc1.w_2[3] ),
    .C(\w_new_calc1.w_2[5] ),
    .X(\w_new_calc1.temp2[18] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_10_  (.A(\w_new_calc1.w_2[29] ),
    .B(\w_new_calc1.w_2[4] ),
    .C(\w_new_calc1.w_2[6] ),
    .X(\w_new_calc1.temp2[19] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_11_  (.A(\w_new_calc1.w_2[20] ),
    .B(\w_new_calc1.w_2[18] ),
    .C(\w_new_calc1.w_2[11] ),
    .X(\w_new_calc1.temp2[1] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_12_  (.A(\w_new_calc1.w_2[30] ),
    .B(\w_new_calc1.w_2[5] ),
    .C(\w_new_calc1.w_2[7] ),
    .X(\w_new_calc1.temp2[20] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_13_  (.A(\w_new_calc1.w_2[31] ),
    .B(\w_new_calc1.w_2[6] ),
    .C(\w_new_calc1.w_2[8] ),
    .X(\w_new_calc1.temp2[21] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_14_  (.A(\w_new_calc1.w_2[7] ),
    .B(\w_new_calc1.w_2[9] ),
    .X(\w_new_calc1.temp2[22] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_15_  (.A(\w_new_calc1.w_2[8] ),
    .B(\w_new_calc1.w_2[10] ),
    .X(\w_new_calc1.temp2[23] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_16_  (.A(\w_new_calc1.w_2[11] ),
    .B(\w_new_calc1.w_2[9] ),
    .X(\w_new_calc1.temp2[24] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_17_  (.A(\w_new_calc1.w_2[10] ),
    .B(\w_new_calc1.w_2[12] ),
    .X(\w_new_calc1.temp2[25] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_18_  (.A(\w_new_calc1.w_2[11] ),
    .B(\w_new_calc1.w_2[13] ),
    .X(\w_new_calc1.temp2[26] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_19_  (.A(\w_new_calc1.w_2[12] ),
    .B(\w_new_calc1.w_2[14] ),
    .X(\w_new_calc1.temp2[27] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_20_  (.A(\w_new_calc1.w_2[13] ),
    .B(\w_new_calc1.w_2[15] ),
    .X(\w_new_calc1.temp2[28] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_21_  (.A(\w_new_calc1.w_2[14] ),
    .B(\w_new_calc1.w_2[16] ),
    .X(\w_new_calc1.temp2[29] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_22_  (.A(\w_new_calc1.w_2[19] ),
    .B(\w_new_calc1.w_2[21] ),
    .C(\w_new_calc1.w_2[12] ),
    .X(\w_new_calc1.temp2[2] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_23_  (.A(\w_new_calc1.w_2[17] ),
    .B(\w_new_calc1.w_2[15] ),
    .X(\w_new_calc1.temp2[30] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc1.s1/_24_  (.A(\w_new_calc1.w_2[18] ),
    .B(\w_new_calc1.w_2[16] ),
    .X(\w_new_calc1.temp2[31] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_25_  (.A(\w_new_calc1.w_2[20] ),
    .B(\w_new_calc1.w_2[22] ),
    .C(\w_new_calc1.w_2[13] ),
    .X(\w_new_calc1.temp2[3] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_26_  (.A(\w_new_calc1.w_2[21] ),
    .B(\w_new_calc1.w_2[23] ),
    .C(\w_new_calc1.w_2[14] ),
    .X(\w_new_calc1.temp2[4] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_27_  (.A(\w_new_calc1.w_2[22] ),
    .B(\w_new_calc1.w_2[24] ),
    .C(\w_new_calc1.w_2[15] ),
    .X(\w_new_calc1.temp2[5] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_28_  (.A(\w_new_calc1.w_2[23] ),
    .B(\w_new_calc1.w_2[25] ),
    .C(\w_new_calc1.w_2[16] ),
    .X(\w_new_calc1.temp2[6] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_29_  (.A(\w_new_calc1.w_2[17] ),
    .B(\w_new_calc1.w_2[24] ),
    .C(\w_new_calc1.w_2[26] ),
    .X(\w_new_calc1.temp2[7] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_30_  (.A(\w_new_calc1.w_2[18] ),
    .B(\w_new_calc1.w_2[25] ),
    .C(\w_new_calc1.w_2[27] ),
    .X(\w_new_calc1.temp2[8] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc1.s1/_31_  (.A(\w_new_calc1.w_2[19] ),
    .B(\w_new_calc1.w_2[26] ),
    .C(\w_new_calc1.w_2[28] ),
    .X(\w_new_calc1.temp2[9] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_00_  (.A(\w_new_calc2.w_15[18] ),
    .B(\w_new_calc2.w_15[7] ),
    .C(\w_new_calc2.w_15[3] ),
    .X(\w_new_calc2.temp1[0] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_01_  (.A(\w_new_calc2.w_15[13] ),
    .B(\w_new_calc2.w_15[28] ),
    .C(\w_new_calc2.w_15[17] ),
    .X(\w_new_calc2.temp1[10] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_02_  (.A(\w_new_calc2.w_15[18] ),
    .B(\w_new_calc2.w_15[14] ),
    .C(\w_new_calc2.w_15[29] ),
    .X(\w_new_calc2.temp1[11] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_03_  (.A(\w_new_calc2.w_15[19] ),
    .B(\w_new_calc2.w_15[15] ),
    .C(\w_new_calc2.w_15[30] ),
    .X(\w_new_calc2.temp1[12] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_04_  (.A(\w_new_calc2.w_15[20] ),
    .B(\w_new_calc2.w_15[16] ),
    .C(\w_new_calc2.w_15[31] ),
    .X(\w_new_calc2.temp1[13] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_05_  (.A(\w_new_calc2.w_15[21] ),
    .B(\w_new_calc2.w_15[17] ),
    .C(\w_new_calc2.w_15[0] ),
    .X(\w_new_calc2.temp1[14] ));
 sky130_fd_sc_hd__xor3_4 \w_new_calc2.s0/_06_  (.A(\w_new_calc2.w_15[18] ),
    .B(\w_new_calc2.w_15[22] ),
    .C(\w_new_calc2.w_15[1] ),
    .X(\w_new_calc2.temp1[15] ));
 sky130_fd_sc_hd__xor3_4 \w_new_calc2.s0/_07_  (.A(\w_new_calc2.w_15[19] ),
    .B(\w_new_calc2.w_15[23] ),
    .C(\w_new_calc2.w_15[2] ),
    .X(\w_new_calc2.temp1[16] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_08_  (.A(\w_new_calc2.w_15[20] ),
    .B(\w_new_calc2.w_15[24] ),
    .C(\w_new_calc2.w_15[3] ),
    .X(\w_new_calc2.temp1[17] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_09_  (.A(\w_new_calc2.w_15[21] ),
    .B(\w_new_calc2.w_15[25] ),
    .C(\w_new_calc2.w_15[4] ),
    .X(\w_new_calc2.temp1[18] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_10_  (.A(\w_new_calc2.w_15[22] ),
    .B(\w_new_calc2.w_15[26] ),
    .C(\w_new_calc2.w_15[5] ),
    .X(\w_new_calc2.temp1[19] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_11_  (.A(\w_new_calc2.w_15[19] ),
    .B(\w_new_calc2.w_15[8] ),
    .C(\w_new_calc2.w_15[4] ),
    .X(\w_new_calc2.temp1[1] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_12_  (.A(\w_new_calc2.w_15[23] ),
    .B(\w_new_calc2.w_15[27] ),
    .C(\w_new_calc2.w_15[6] ),
    .X(\w_new_calc2.temp1[20] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_13_  (.A(\w_new_calc2.w_15[7] ),
    .B(\w_new_calc2.w_15[24] ),
    .C(\w_new_calc2.w_15[28] ),
    .X(\w_new_calc2.temp1[21] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_14_  (.A(\w_new_calc2.w_15[8] ),
    .B(\w_new_calc2.w_15[25] ),
    .C(\w_new_calc2.w_15[29] ),
    .X(\w_new_calc2.temp1[22] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_15_  (.A(\w_new_calc2.w_15[9] ),
    .B(\w_new_calc2.w_15[26] ),
    .C(\w_new_calc2.w_15[30] ),
    .X(\w_new_calc2.temp1[23] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_16_  (.A(\w_new_calc2.w_15[10] ),
    .B(\w_new_calc2.w_15[27] ),
    .C(\w_new_calc2.w_15[31] ),
    .X(\w_new_calc2.temp1[24] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_17_  (.A(\w_new_calc2.w_15[11] ),
    .B(\w_new_calc2.w_15[28] ),
    .C(\w_new_calc2.w_15[0] ),
    .X(\w_new_calc2.temp1[25] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_18_  (.A(\w_new_calc2.w_15[12] ),
    .B(\w_new_calc2.w_15[29] ),
    .C(\w_new_calc2.w_15[1] ),
    .X(\w_new_calc2.temp1[26] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_19_  (.A(\w_new_calc2.w_15[13] ),
    .B(\w_new_calc2.w_15[30] ),
    .C(\w_new_calc2.w_15[2] ),
    .X(\w_new_calc2.temp1[27] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_20_  (.A(\w_new_calc2.w_15[14] ),
    .B(\w_new_calc2.w_15[31] ),
    .C(\w_new_calc2.w_15[3] ),
    .X(\w_new_calc2.temp1[28] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s0/_21_  (.A(\w_new_calc2.w_15[15] ),
    .B(\w_new_calc2.w_15[4] ),
    .X(\w_new_calc2.temp1[29] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_22_  (.A(\w_new_calc2.w_15[20] ),
    .B(\w_new_calc2.w_15[9] ),
    .C(\w_new_calc2.w_15[5] ),
    .X(\w_new_calc2.temp1[2] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s0/_23_  (.A(\w_new_calc2.w_15[16] ),
    .B(\w_new_calc2.w_15[5] ),
    .X(\w_new_calc2.temp1[30] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s0/_24_  (.A(\w_new_calc2.w_15[17] ),
    .B(\w_new_calc2.w_15[6] ),
    .X(\w_new_calc2.temp1[31] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_25_  (.A(\w_new_calc2.w_15[21] ),
    .B(\w_new_calc2.w_15[10] ),
    .C(\w_new_calc2.w_15[6] ),
    .X(\w_new_calc2.temp1[3] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_26_  (.A(\w_new_calc2.w_15[7] ),
    .B(\w_new_calc2.w_15[22] ),
    .C(\w_new_calc2.w_15[11] ),
    .X(\w_new_calc2.temp1[4] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_27_  (.A(\w_new_calc2.w_15[8] ),
    .B(\w_new_calc2.w_15[23] ),
    .C(\w_new_calc2.w_15[12] ),
    .X(\w_new_calc2.temp1[5] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_28_  (.A(\w_new_calc2.w_15[9] ),
    .B(\w_new_calc2.w_15[24] ),
    .C(\w_new_calc2.w_15[13] ),
    .X(\w_new_calc2.temp1[6] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_29_  (.A(\w_new_calc2.w_15[10] ),
    .B(\w_new_calc2.w_15[25] ),
    .C(\w_new_calc2.w_15[14] ),
    .X(\w_new_calc2.temp1[7] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_30_  (.A(\w_new_calc2.w_15[11] ),
    .B(\w_new_calc2.w_15[26] ),
    .C(\w_new_calc2.w_15[15] ),
    .X(\w_new_calc2.temp1[8] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s0/_31_  (.A(\w_new_calc2.w_15[12] ),
    .B(\w_new_calc2.w_15[27] ),
    .C(\w_new_calc2.w_15[16] ),
    .X(\w_new_calc2.temp1[9] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_00_  (.A(\w_new_calc2.w_2[19] ),
    .B(\w_new_calc2.w_2[17] ),
    .C(\w_new_calc2.w_2[10] ),
    .X(\w_new_calc2.temp2[0] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_01_  (.A(\w_new_calc2.w_2[20] ),
    .B(\w_new_calc2.w_2[27] ),
    .C(\w_new_calc2.w_2[29] ),
    .X(\w_new_calc2.temp2[10] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_02_  (.A(\w_new_calc2.w_2[21] ),
    .B(\w_new_calc2.w_2[28] ),
    .C(\w_new_calc2.w_2[30] ),
    .X(\w_new_calc2.temp2[11] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_03_  (.A(\w_new_calc2.w_2[22] ),
    .B(\w_new_calc2.w_2[29] ),
    .C(\w_new_calc2.w_2[31] ),
    .X(\w_new_calc2.temp2[12] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_04_  (.A(\w_new_calc2.w_2[23] ),
    .B(\w_new_calc2.w_2[30] ),
    .C(\w_new_calc2.w_2[0] ),
    .X(\w_new_calc2.temp2[13] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_05_  (.A(\w_new_calc2.w_2[24] ),
    .B(\w_new_calc2.w_2[31] ),
    .C(\w_new_calc2.w_2[1] ),
    .X(\w_new_calc2.temp2[14] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_06_  (.A(\w_new_calc2.w_2[25] ),
    .B(\w_new_calc2.w_2[0] ),
    .C(\w_new_calc2.w_2[2] ),
    .X(\w_new_calc2.temp2[15] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_07_  (.A(\w_new_calc2.w_2[26] ),
    .B(\w_new_calc2.w_2[1] ),
    .C(\w_new_calc2.w_2[3] ),
    .X(\w_new_calc2.temp2[16] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_08_  (.A(\w_new_calc2.w_2[27] ),
    .B(\w_new_calc2.w_2[2] ),
    .C(\w_new_calc2.w_2[4] ),
    .X(\w_new_calc2.temp2[17] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_09_  (.A(\w_new_calc2.w_2[28] ),
    .B(\w_new_calc2.w_2[3] ),
    .C(\w_new_calc2.w_2[5] ),
    .X(\w_new_calc2.temp2[18] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_10_  (.A(\w_new_calc2.w_2[29] ),
    .B(\w_new_calc2.w_2[4] ),
    .C(\w_new_calc2.w_2[6] ),
    .X(\w_new_calc2.temp2[19] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_11_  (.A(\w_new_calc2.w_2[20] ),
    .B(\w_new_calc2.w_2[18] ),
    .C(\w_new_calc2.w_2[11] ),
    .X(\w_new_calc2.temp2[1] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_12_  (.A(\w_new_calc2.w_2[30] ),
    .B(\w_new_calc2.w_2[5] ),
    .C(\w_new_calc2.w_2[7] ),
    .X(\w_new_calc2.temp2[20] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_13_  (.A(\w_new_calc2.w_2[31] ),
    .B(\w_new_calc2.w_2[6] ),
    .C(\w_new_calc2.w_2[8] ),
    .X(\w_new_calc2.temp2[21] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_14_  (.A(\w_new_calc2.w_2[7] ),
    .B(\w_new_calc2.w_2[9] ),
    .X(\w_new_calc2.temp2[22] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_15_  (.A(\w_new_calc2.w_2[8] ),
    .B(\w_new_calc2.w_2[10] ),
    .X(\w_new_calc2.temp2[23] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_16_  (.A(\w_new_calc2.w_2[11] ),
    .B(\w_new_calc2.w_2[9] ),
    .X(\w_new_calc2.temp2[24] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_17_  (.A(\w_new_calc2.w_2[10] ),
    .B(\w_new_calc2.w_2[12] ),
    .X(\w_new_calc2.temp2[25] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_18_  (.A(\w_new_calc2.w_2[11] ),
    .B(\w_new_calc2.w_2[13] ),
    .X(\w_new_calc2.temp2[26] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_19_  (.A(\w_new_calc2.w_2[12] ),
    .B(\w_new_calc2.w_2[14] ),
    .X(\w_new_calc2.temp2[27] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_20_  (.A(\w_new_calc2.w_2[13] ),
    .B(\w_new_calc2.w_2[15] ),
    .X(\w_new_calc2.temp2[28] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_21_  (.A(\w_new_calc2.w_2[14] ),
    .B(\w_new_calc2.w_2[16] ),
    .X(\w_new_calc2.temp2[29] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_22_  (.A(\w_new_calc2.w_2[19] ),
    .B(\w_new_calc2.w_2[21] ),
    .C(\w_new_calc2.w_2[12] ),
    .X(\w_new_calc2.temp2[2] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_23_  (.A(\w_new_calc2.w_2[17] ),
    .B(\w_new_calc2.w_2[15] ),
    .X(\w_new_calc2.temp2[30] ));
 sky130_fd_sc_hd__xor2_1 \w_new_calc2.s1/_24_  (.A(\w_new_calc2.w_2[18] ),
    .B(\w_new_calc2.w_2[16] ),
    .X(\w_new_calc2.temp2[31] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_25_  (.A(\w_new_calc2.w_2[20] ),
    .B(\w_new_calc2.w_2[22] ),
    .C(\w_new_calc2.w_2[13] ),
    .X(\w_new_calc2.temp2[3] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_26_  (.A(\w_new_calc2.w_2[21] ),
    .B(\w_new_calc2.w_2[23] ),
    .C(\w_new_calc2.w_2[14] ),
    .X(\w_new_calc2.temp2[4] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_27_  (.A(\w_new_calc2.w_2[22] ),
    .B(\w_new_calc2.w_2[24] ),
    .C(\w_new_calc2.w_2[15] ),
    .X(\w_new_calc2.temp2[5] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_28_  (.A(\w_new_calc2.w_2[23] ),
    .B(\w_new_calc2.w_2[25] ),
    .C(\w_new_calc2.w_2[16] ),
    .X(\w_new_calc2.temp2[6] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_29_  (.A(\w_new_calc2.w_2[17] ),
    .B(\w_new_calc2.w_2[24] ),
    .C(\w_new_calc2.w_2[26] ),
    .X(\w_new_calc2.temp2[7] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_30_  (.A(\w_new_calc2.w_2[18] ),
    .B(\w_new_calc2.w_2[25] ),
    .C(\w_new_calc2.w_2[27] ),
    .X(\w_new_calc2.temp2[8] ));
 sky130_fd_sc_hd__xor3_1 \w_new_calc2.s1/_31_  (.A(\w_new_calc2.w_2[19] ),
    .B(\w_new_calc2.w_2[26] ),
    .C(\w_new_calc2.w_2[28] ),
    .X(\w_new_calc2.temp2[9] ));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[0]$_DFF_P_  (.D(_00000_),
    .Q(\w_value1[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[10]$_DFF_P_  (.D(_00001_),
    .Q(\w_value1[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[11]$_DFF_P_  (.D(_00002_),
    .Q(\w_value1[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[12]$_DFF_P_  (.D(_00003_),
    .Q(\w_value1[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[13]$_DFF_P_  (.D(_00004_),
    .Q(\w_value1[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[14]$_DFF_P_  (.D(_00005_),
    .Q(\w_value1[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[15]$_DFF_P_  (.D(_00006_),
    .Q(\w_value1[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[16]$_DFF_P_  (.D(_00007_),
    .Q(\w_value1[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[17]$_DFF_P_  (.D(_00008_),
    .Q(\w_value1[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[18]$_DFF_P_  (.D(_00009_),
    .Q(\w_value1[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[19]$_DFF_P_  (.D(_00010_),
    .Q(\w_value1[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[1]$_DFF_P_  (.D(_00011_),
    .Q(\w_value1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[20]$_DFF_P_  (.D(_00012_),
    .Q(\w_value1[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[21]$_DFF_P_  (.D(_00013_),
    .Q(\w_value1[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[22]$_DFF_P_  (.D(_00014_),
    .Q(\w_value1[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[23]$_DFF_P_  (.D(_00015_),
    .Q(\w_value1[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[24]$_DFF_P_  (.D(_00016_),
    .Q(\w_value1[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[25]$_DFF_P_  (.D(_00017_),
    .Q(\w_value1[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[26]$_DFF_P_  (.D(_00018_),
    .Q(\w_value1[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[27]$_DFF_P_  (.D(_00019_),
    .Q(\w_value1[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[28]$_DFF_P_  (.D(_00020_),
    .Q(\w_value1[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[29]$_DFF_P_  (.D(_00021_),
    .Q(\w_value1[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[2]$_DFF_P_  (.D(_00022_),
    .Q(\w_value1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[30]$_DFF_P_  (.D(_00023_),
    .Q(\w_value1[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[31]$_DFF_P_  (.D(_00024_),
    .Q(\w_value1[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[3]$_DFF_P_  (.D(_00025_),
    .Q(\w_value1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[4]$_DFF_P_  (.D(_00026_),
    .Q(\w_value1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[5]$_DFF_P_  (.D(_00027_),
    .Q(\w_value1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[6]$_DFF_P_  (.D(_00028_),
    .Q(\w_value1[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[7]$_DFF_P_  (.D(_00029_),
    .Q(\w_value1[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[8]$_DFF_P_  (.D(_00030_),
    .Q(\w_value1[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[9]$_DFF_P_  (.D(_00031_),
    .Q(\w_value1[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[0]$_DFF_P_  (.D(_00032_),
    .Q(\w_value2[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[10]$_DFF_P_  (.D(_00033_),
    .Q(\w_value2[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[11]$_DFF_P_  (.D(_00034_),
    .Q(\w_value2[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[12]$_DFF_P_  (.D(_00035_),
    .Q(\w_value2[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[13]$_DFF_P_  (.D(_00036_),
    .Q(\w_value2[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[14]$_DFF_P_  (.D(_00037_),
    .Q(\w_value2[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[15]$_DFF_P_  (.D(_00038_),
    .Q(\w_value2[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[16]$_DFF_P_  (.D(_00039_),
    .Q(\w_value2[16] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[17]$_DFF_P_  (.D(_00040_),
    .Q(\w_value2[17] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[18]$_DFF_P_  (.D(_00041_),
    .Q(\w_value2[18] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[19]$_DFF_P_  (.D(_00042_),
    .Q(\w_value2[19] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[1]$_DFF_P_  (.D(_00043_),
    .Q(\w_value2[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[20]$_DFF_P_  (.D(_00044_),
    .Q(\w_value2[20] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[21]$_DFF_P_  (.D(_00045_),
    .Q(\w_value2[21] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[22]$_DFF_P_  (.D(_00046_),
    .Q(\w_value2[22] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[23]$_DFF_P_  (.D(_00047_),
    .Q(\w_value2[23] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[24]$_DFF_P_  (.D(_00048_),
    .Q(\w_value2[24] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[25]$_DFF_P_  (.D(_00049_),
    .Q(\w_value2[25] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[26]$_DFF_P_  (.D(_00050_),
    .Q(\w_value2[26] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[27]$_DFF_P_  (.D(_00051_),
    .Q(\w_value2[27] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[28]$_DFF_P_  (.D(_00052_),
    .Q(\w_value2[28] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[29]$_DFF_P_  (.D(_00053_),
    .Q(\w_value2[29] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[2]$_DFF_P_  (.D(_00054_),
    .Q(\w_value2[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[30]$_DFF_P_  (.D(_00055_),
    .Q(\w_value2[30] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[31]$_DFF_P_  (.D(_00056_),
    .Q(\w_value2[31] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[3]$_DFF_P_  (.D(_00057_),
    .Q(\w_value2[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[4]$_DFF_P_  (.D(_00058_),
    .Q(\w_value2[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[5]$_DFF_P_  (.D(_00059_),
    .Q(\w_value2[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[6]$_DFF_P_  (.D(_00060_),
    .Q(\w_value2[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[7]$_DFF_P_  (.D(_00061_),
    .Q(\w_value2[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[8]$_DFF_P_  (.D(_00062_),
    .Q(\w_value2[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[9]$_DFF_P_  (.D(_00063_),
    .Q(\w_value2[9] ),
    .CLK(clk));
endmodule
