module sha256_unrolled_pipelined (clk,
    ready,
    reset,
    hashvalue,
    message);
 input clk;
 output ready;
 input reset;
 output [255:0] hashvalue;
 input [0:511] message;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire net376;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire net10;
 wire net9;
 wire _02682_;
 wire net8;
 wire net7;
 wire _02685_;
 wire net6;
 wire net5;
 wire _02688_;
 wire net4;
 wire net3;
 wire _02691_;
 wire net2;
 wire net1;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire net701;
 wire net700;
 wire _02699_;
 wire net699;
 wire net698;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire net697;
 wire net696;
 wire _02708_;
 wire net695;
 wire net694;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire net693;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire net692;
 wire net691;
 wire net690;
 wire net689;
 wire net688;
 wire net687;
 wire net686;
 wire net685;
 wire net684;
 wire _02886_;
 wire net683;
 wire net682;
 wire _02889_;
 wire _02890_;
 wire net681;
 wire net680;
 wire net679;
 wire _02894_;
 wire net678;
 wire net677;
 wire net676;
 wire net675;
 wire net674;
 wire _02900_;
 wire _02901_;
 wire net673;
 wire net672;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire net671;
 wire net670;
 wire _02910_;
 wire net669;
 wire net668;
 wire net667;
 wire _02914_;
 wire net666;
 wire net665;
 wire _02917_;
 wire net664;
 wire net663;
 wire _02920_;
 wire net662;
 wire _02922_;
 wire net661;
 wire net660;
 wire _02925_;
 wire net659;
 wire _02927_;
 wire net658;
 wire net657;
 wire _02930_;
 wire net656;
 wire net655;
 wire _02933_;
 wire net654;
 wire net653;
 wire _02936_;
 wire net652;
 wire net651;
 wire _02939_;
 wire net650;
 wire _02941_;
 wire net649;
 wire _02943_;
 wire net648;
 wire net647;
 wire _02946_;
 wire _02947_;
 wire net646;
 wire net645;
 wire _02950_;
 wire net644;
 wire net643;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire net642;
 wire net641;
 wire net640;
 wire net639;
 wire net638;
 wire net637;
 wire net636;
 wire net635;
 wire net634;
 wire _02970_;
 wire net633;
 wire net632;
 wire net631;
 wire net630;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire net629;
 wire net628;
 wire net627;
 wire net626;
 wire net625;
 wire _02983_;
 wire _02984_;
 wire net624;
 wire net623;
 wire net622;
 wire net621;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire net620;
 wire net619;
 wire _02995_;
 wire net618;
 wire net617;
 wire _02998_;
 wire net616;
 wire net615;
 wire _03001_;
 wire net614;
 wire net613;
 wire _03004_;
 wire net612;
 wire net611;
 wire _03007_;
 wire net610;
 wire net609;
 wire _03010_;
 wire _03011_;
 wire net608;
 wire _03013_;
 wire net607;
 wire net606;
 wire _03016_;
 wire net605;
 wire net604;
 wire _03019_;
 wire net603;
 wire net602;
 wire _03022_;
 wire net601;
 wire _03024_;
 wire net600;
 wire net599;
 wire _03027_;
 wire net598;
 wire net597;
 wire _03030_;
 wire net596;
 wire _03032_;
 wire net595;
 wire _03034_;
 wire net594;
 wire net593;
 wire _03037_;
 wire net592;
 wire net591;
 wire _03040_;
 wire net590;
 wire net589;
 wire _03043_;
 wire net588;
 wire net587;
 wire _03046_;
 wire net586;
 wire net585;
 wire _03049_;
 wire net584;
 wire net583;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire net582;
 wire net581;
 wire net580;
 wire net579;
 wire net578;
 wire net577;
 wire net576;
 wire net575;
 wire _03063_;
 wire net574;
 wire net573;
 wire net572;
 wire net571;
 wire _03068_;
 wire net570;
 wire net569;
 wire _03071_;
 wire net568;
 wire net567;
 wire net566;
 wire _03075_;
 wire net565;
 wire net564;
 wire net563;
 wire net562;
 wire net561;
 wire _03081_;
 wire net560;
 wire net559;
 wire _03084_;
 wire net558;
 wire net557;
 wire _03087_;
 wire net556;
 wire net555;
 wire _03090_;
 wire net554;
 wire net553;
 wire _03093_;
 wire net552;
 wire net551;
 wire _03096_;
 wire net550;
 wire net549;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire net548;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire net547;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire net546;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire net545;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire net544;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire net543;
 wire net542;
 wire _03158_;
 wire net541;
 wire net540;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire net539;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire net538;
 wire net537;
 wire net536;
 wire net535;
 wire net534;
 wire net533;
 wire net532;
 wire net531;
 wire _03195_;
 wire net530;
 wire net529;
 wire net528;
 wire net527;
 wire _03200_;
 wire net526;
 wire net525;
 wire _03203_;
 wire net524;
 wire net523;
 wire net522;
 wire _03207_;
 wire net521;
 wire net520;
 wire net519;
 wire net518;
 wire net517;
 wire _03213_;
 wire net516;
 wire net515;
 wire _03216_;
 wire net514;
 wire net513;
 wire _03219_;
 wire net512;
 wire net511;
 wire _03222_;
 wire net510;
 wire net509;
 wire _03225_;
 wire net508;
 wire net507;
 wire _03228_;
 wire net506;
 wire net505;
 wire net504;
 wire _03232_;
 wire net503;
 wire net502;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire net501;
 wire net500;
 wire _03244_;
 wire net499;
 wire _03246_;
 wire net498;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire net497;
 wire net496;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire net495;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire net494;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire net493;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire net492;
 wire net491;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire net490;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire net489;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire net488;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire net487;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire net486;
 wire _03455_;
 wire _03456_;
 wire net485;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire net484;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire net483;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire net482;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire net481;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire net480;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire net479;
 wire _03597_;
 wire net478;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire net477;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire net476;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire net475;
 wire _03656_;
 wire net474;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire net473;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire net472;
 wire _03709_;
 wire net471;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire net470;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire net469;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire net468;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire net467;
 wire _03776_;
 wire net466;
 wire _03778_;
 wire net465;
 wire _03780_;
 wire net464;
 wire _03782_;
 wire net463;
 wire _03784_;
 wire net462;
 wire _03786_;
 wire net461;
 wire _03788_;
 wire net460;
 wire _03790_;
 wire net459;
 wire _03792_;
 wire net458;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire net457;
 wire net456;
 wire _03842_;
 wire net455;
 wire _03844_;
 wire net454;
 wire _03846_;
 wire net453;
 wire _03848_;
 wire _03849_;
 wire _03851_;
 wire _03853_;
 wire net1169;
 wire _03855_;
 wire net1168;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire net1167;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire net1166;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire net1165;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire net1164;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire net1163;
 wire net1162;
 wire _03953_;
 wire net1161;
 wire net1160;
 wire _03956_;
 wire net1159;
 wire net1152;
 wire _03959_;
 wire net1151;
 wire net1150;
 wire _03962_;
 wire net1115;
 wire net1114;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire net1109;
 wire net1106;
 wire _03970_;
 wire net1142;
 wire net1141;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire net1140;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire net1139;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire net1138;
 wire _04025_;
 wire net1137;
 wire net1136;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire net1135;
 wire _04044_;
 wire _04045_;
 wire net1134;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire net1133;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire net1132;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire net1131;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire net1130;
 wire _04140_;
 wire net1129;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire net1128;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire net1127;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire net1126;
 wire _04177_;
 wire net1125;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire net1124;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire net1123;
 wire _04208_;
 wire net1122;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire net1121;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire net1120;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire net1119;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire net1118;
 wire _04253_;
 wire net1113;
 wire _04255_;
 wire net1112;
 wire _04257_;
 wire net1157;
 wire _04259_;
 wire net1110;
 wire _04261_;
 wire net1105;
 wire _04263_;
 wire net1104;
 wire _04265_;
 wire net1158;
 wire _04267_;
 wire net1102;
 wire _04269_;
 wire net1101;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire net1100;
 wire net1099;
 wire _04297_;
 wire net1098;
 wire _04299_;
 wire net1097;
 wire _04301_;
 wire net1096;
 wire _04303_;
 wire _04304_;
 wire net1095;
 wire _04306_;
 wire net1094;
 wire _04308_;
 wire net1093;
 wire _04310_;
 wire net1092;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire net1091;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire net1090;
 wire net1089;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire net1088;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire net1087;
 wire net1086;
 wire net1085;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire net1084;
 wire net1083;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire net1082;
 wire _04565_;
 wire net1081;
 wire _04567_;
 wire net1080;
 wire net1079;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire net1078;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire net1077;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire net1076;
 wire net1075;
 wire net1074;
 wire _04616_;
 wire net1073;
 wire net1072;
 wire net1071;
 wire _04620_;
 wire net1070;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire net1069;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire net1068;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire net1067;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire net1066;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire net1065;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire net1064;
 wire _04984_;
 wire net1063;
 wire net1062;
 wire net1149;
 wire _04988_;
 wire net1107;
 wire net1108;
 wire _04991_;
 wire _04992_;
 wire net1058;
 wire _04994_;
 wire _04995_;
 wire net1057;
 wire _04997_;
 wire net1056;
 wire net1055;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire net1054;
 wire _05005_;
 wire net1053;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire net1052;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire net1051;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire net1050;
 wire _05031_;
 wire _05032_;
 wire net1049;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire net1048;
 wire _05041_;
 wire net1047;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire net1046;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire net1045;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire net1044;
 wire net1043;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire net1042;
 wire _05079_;
 wire net1041;
 wire net1040;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire net1039;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire net1038;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire net1037;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire net1036;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire net1035;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire net1034;
 wire _05130_;
 wire net1033;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire net1032;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire net1031;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire net1030;
 wire net1029;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire net1028;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire net1027;
 wire _05186_;
 wire net1026;
 wire net1025;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire net1024;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire net1156;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire net1022;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire net1021;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire net1020;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire clknet_5_31__leaf_clk;
 wire _05243_;
 wire clknet_5_30__leaf_clk;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire clknet_5_29__leaf_clk;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire clknet_5_28__leaf_clk;
 wire _05262_;
 wire _05263_;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire clknet_5_23__leaf_clk;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire clknet_5_22__leaf_clk;
 wire _05280_;
 wire _05281_;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire clknet_5_17__leaf_clk;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire clknet_5_16__leaf_clk;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire clknet_5_15__leaf_clk;
 wire _05312_;
 wire _05313_;
 wire clknet_5_14__leaf_clk;
 wire _05315_;
 wire clknet_5_13__leaf_clk;
 wire _05317_;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire _05320_;
 wire _05321_;
 wire clknet_5_10__leaf_clk;
 wire _05323_;
 wire _05324_;
 wire clknet_5_9__leaf_clk;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire clknet_5_8__leaf_clk;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire clknet_5_7__leaf_clk;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire clknet_5_6__leaf_clk;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire clknet_5_5__leaf_clk;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire clknet_5_4__leaf_clk;
 wire _05362_;
 wire clknet_5_3__leaf_clk;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire clknet_5_2__leaf_clk;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire clknet_5_1__leaf_clk;
 wire _05382_;
 wire clknet_5_0__leaf_clk;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire clknet_2_3_0_clk;
 wire clknet_2_2_0_clk;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire clknet_2_1_0_clk;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire clknet_2_0_0_clk;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire clknet_0_clk;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire clknet_leaf_284_clk;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire clknet_leaf_283_clk;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire clknet_leaf_282_clk;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire clknet_leaf_281_clk;
 wire _05455_;
 wire clknet_leaf_280_clk;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire clknet_leaf_279_clk;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire clknet_leaf_278_clk;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_276_clk;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire clknet_leaf_275_clk;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire clknet_leaf_274_clk;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire clknet_leaf_273_clk;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire clknet_leaf_272_clk;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire clknet_leaf_271_clk;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire clknet_leaf_270_clk;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire clknet_leaf_269_clk;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire clknet_leaf_268_clk;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire clknet_leaf_267_clk;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire clknet_leaf_266_clk;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire clknet_leaf_265_clk;
 wire _05613_;
 wire _05614_;
 wire clknet_leaf_264_clk;
 wire _05616_;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_262_clk;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire clknet_leaf_261_clk;
 wire _05628_;
 wire _05629_;
 wire clknet_leaf_260_clk;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire clknet_leaf_259_clk;
 wire _05640_;
 wire _05641_;
 wire clknet_leaf_258_clk;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire clknet_leaf_257_clk;
 wire _05657_;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_255_clk;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire clknet_leaf_254_clk;
 wire _05669_;
 wire _05670_;
 wire clknet_leaf_253_clk;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire clknet_leaf_252_clk;
 wire _05681_;
 wire _05682_;
 wire clknet_leaf_251_clk;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire clknet_leaf_250_clk;
 wire _05698_;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_248_clk;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire clknet_leaf_247_clk;
 wire _05710_;
 wire _05711_;
 wire clknet_leaf_246_clk;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire clknet_leaf_245_clk;
 wire _05722_;
 wire _05723_;
 wire clknet_leaf_244_clk;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire clknet_leaf_243_clk;
 wire _05739_;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_241_clk;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire clknet_leaf_240_clk;
 wire _05751_;
 wire _05752_;
 wire clknet_leaf_239_clk;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire clknet_leaf_238_clk;
 wire _05763_;
 wire _05764_;
 wire clknet_leaf_237_clk;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire clknet_leaf_236_clk;
 wire _05780_;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_234_clk;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire clknet_leaf_233_clk;
 wire _05792_;
 wire _05793_;
 wire clknet_leaf_232_clk;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire clknet_leaf_231_clk;
 wire _05804_;
 wire _05805_;
 wire clknet_leaf_230_clk;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_228_clk;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire clknet_leaf_227_clk;
 wire _05833_;
 wire _05834_;
 wire clknet_leaf_226_clk;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire clknet_leaf_225_clk;
 wire _05845_;
 wire _05846_;
 wire clknet_leaf_224_clk;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_222_clk;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire clknet_leaf_221_clk;
 wire _05872_;
 wire _05873_;
 wire clknet_leaf_220_clk;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire clknet_leaf_219_clk;
 wire _05884_;
 wire _05885_;
 wire clknet_leaf_218_clk;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_216_clk;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire clknet_leaf_215_clk;
 wire _05911_;
 wire _05912_;
 wire clknet_leaf_214_clk;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire clknet_leaf_213_clk;
 wire _05923_;
 wire _05924_;
 wire clknet_leaf_212_clk;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_210_clk;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire clknet_leaf_209_clk;
 wire _05950_;
 wire _05951_;
 wire clknet_leaf_208_clk;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire clknet_leaf_207_clk;
 wire _05962_;
 wire _05963_;
 wire clknet_leaf_206_clk;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_204_clk;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire clknet_leaf_203_clk;
 wire _05989_;
 wire _05990_;
 wire clknet_leaf_202_clk;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire clknet_leaf_201_clk;
 wire _06001_;
 wire _06002_;
 wire clknet_leaf_200_clk;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_198_clk;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire clknet_leaf_197_clk;
 wire _06028_;
 wire _06029_;
 wire clknet_leaf_196_clk;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire clknet_leaf_195_clk;
 wire _06040_;
 wire _06041_;
 wire clknet_leaf_194_clk;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_192_clk;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire clknet_leaf_191_clk;
 wire _06067_;
 wire _06068_;
 wire clknet_leaf_190_clk;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire clknet_leaf_189_clk;
 wire _06079_;
 wire _06080_;
 wire clknet_leaf_188_clk;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_186_clk;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire clknet_leaf_185_clk;
 wire _06106_;
 wire _06107_;
 wire clknet_leaf_184_clk;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire clknet_leaf_183_clk;
 wire _06118_;
 wire _06119_;
 wire clknet_leaf_182_clk;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_180_clk;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire clknet_leaf_179_clk;
 wire _06146_;
 wire _06147_;
 wire clknet_leaf_178_clk;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire clknet_leaf_177_clk;
 wire _06158_;
 wire _06159_;
 wire clknet_leaf_176_clk;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_173_clk;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire clknet_leaf_172_clk;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire clknet_leaf_171_clk;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire clknet_leaf_170_clk;
 wire _06209_;
 wire _06210_;
 wire clknet_leaf_169_clk;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire clknet_leaf_168_clk;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire clknet_leaf_167_clk;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire clknet_leaf_166_clk;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire clknet_leaf_165_clk;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_163_clk;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_160_clk;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_157_clk;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_154_clk;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire clknet_leaf_153_clk;
 wire _06351_;
 wire _06352_;
 wire clknet_leaf_152_clk;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire clknet_leaf_151_clk;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire clknet_leaf_150_clk;
 wire _06431_;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_147_clk;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_145_clk;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire clknet_leaf_144_clk;
 wire _06469_;
 wire _06470_;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_141_clk;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire clknet_leaf_136_clk;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire clknet_leaf_135_clk;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire clknet_leaf_134_clk;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire clknet_leaf_133_clk;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire clknet_leaf_132_clk;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire clknet_leaf_131_clk;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire clknet_leaf_130_clk;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire clknet_leaf_129_clk;
 wire _06616_;
 wire _06617_;
 wire clknet_leaf_128_clk;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire clknet_leaf_127_clk;
 wire _06631_;
 wire _06632_;
 wire clknet_leaf_126_clk;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire clknet_leaf_125_clk;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire clknet_leaf_124_clk;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire clknet_leaf_123_clk;
 wire _06647_;
 wire clknet_leaf_122_clk;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire clknet_leaf_121_clk;
 wire _06654_;
 wire _06655_;
 wire clknet_leaf_120_clk;
 wire _06657_;
 wire _06658_;
 wire clknet_leaf_119_clk;
 wire _06660_;
 wire clknet_leaf_118_clk;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire clknet_leaf_117_clk;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire clknet_leaf_115_clk;
 wire _06676_;
 wire clknet_leaf_114_clk;
 wire _06678_;
 wire _06679_;
 wire clknet_leaf_113_clk;
 wire _06681_;
 wire clknet_leaf_112_clk;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire clknet_leaf_111_clk;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire clknet_leaf_108_clk;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire clknet_leaf_107_clk;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire clknet_leaf_105_clk;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire clknet_leaf_104_clk;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire clknet_leaf_103_clk;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire clknet_leaf_102_clk;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_99_clk;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire clknet_leaf_98_clk;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_94_clk;
 wire _07359_;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_90_clk;
 wire _07364_;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_88_clk;
 wire _07367_;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_85_clk;
 wire _07371_;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_81_clk;
 wire _07376_;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_79_clk;
 wire _07379_;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_77_clk;
 wire _07382_;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_75_clk;
 wire _07385_;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_73_clk;
 wire _07388_;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_71_clk;
 wire _07391_;
 wire clknet_leaf_70_clk;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire clknet_leaf_69_clk;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire clknet_leaf_68_clk;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire clknet_leaf_67_clk;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire clknet_leaf_66_clk;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire clknet_leaf_65_clk;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire clknet_leaf_64_clk;
 wire _07434_;
 wire _07435_;
 wire clknet_leaf_63_clk;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire clknet_leaf_62_clk;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire clknet_leaf_61_clk;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire clknet_leaf_60_clk;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire clknet_leaf_59_clk;
 wire _07462_;
 wire clknet_leaf_58_clk;
 wire _07464_;
 wire clknet_leaf_57_clk;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire clknet_leaf_56_clk;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire clknet_leaf_55_clk;
 wire _07476_;
 wire clknet_leaf_54_clk;
 wire _07478_;
 wire clknet_leaf_53_clk;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire clknet_leaf_52_clk;
 wire _07484_;
 wire clknet_leaf_51_clk;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire clknet_leaf_50_clk;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire clknet_leaf_49_clk;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire clknet_leaf_48_clk;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire clknet_leaf_47_clk;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire clknet_leaf_46_clk;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire clknet_leaf_45_clk;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire clknet_leaf_44_clk;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire clknet_leaf_43_clk;
 wire _07555_;
 wire _07556_;
 wire clknet_leaf_42_clk;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire clknet_leaf_41_clk;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire clknet_leaf_40_clk;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire clknet_leaf_39_clk;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire clknet_leaf_38_clk;
 wire _07583_;
 wire clknet_leaf_37_clk;
 wire _07585_;
 wire clknet_leaf_36_clk;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire clknet_leaf_35_clk;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire clknet_leaf_34_clk;
 wire _07597_;
 wire clknet_leaf_33_clk;
 wire _07599_;
 wire clknet_leaf_32_clk;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire clknet_leaf_31_clk;
 wire _07605_;
 wire clknet_leaf_30_clk;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire clknet_leaf_29_clk;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire clknet_leaf_28_clk;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire clknet_leaf_27_clk;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_23_clk;
 wire _07740_;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_19_clk;
 wire _07745_;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_17_clk;
 wire _07748_;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire _07752_;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_10_clk;
 wire _07757_;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_8_clk;
 wire _07760_;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_6_clk;
 wire _07763_;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_4_clk;
 wire _07766_;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_2_clk;
 wire _07769_;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_0_clk;
 wire _07772_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07815_;
 wire _07816_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07843_;
 wire _07845_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07857_;
 wire _07859_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07865_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07936_;
 wire _07937_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07964_;
 wire _07966_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07978_;
 wire _07980_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07986_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08467_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08534_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08575_;
 wire _08578_;
 wire _08579_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08747_;
 wire _08749_;
 wire _08750_;
 wire _08752_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08760_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08770_;
 wire _08772_;
 wire _08773_;
 wire _08775_;
 wire _08776_;
 wire _08778_;
 wire _08780_;
 wire _08782_;
 wire _08783_;
 wire _08785_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08808_;
 wire _08809_;
 wire _08811_;
 wire _08813_;
 wire _08814_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09020_;
 wire _09056_;
 wire _09091_;
 wire _09095_;
 wire _09099_;
 wire _09103_;
 wire _09107_;
 wire _09111_;
 wire _09116_;
 wire _09120_;
 wire _09124_;
 wire _09128_;
 wire _09132_;
 wire _09136_;
 wire _09140_;
 wire _09144_;
 wire _09148_;
 wire _09152_;
 wire _09156_;
 wire _09160_;
 wire _09165_;
 wire net762;
 wire net761;
 wire net760;
 wire net759;
 wire net758;
 wire net757;
 wire _09201_;
 wire net756;
 wire net755;
 wire net754;
 wire net753;
 wire net752;
 wire net751;
 wire net750;
 wire net749;
 wire net748;
 wire net747;
 wire net746;
 wire net745;
 wire net744;
 wire net743;
 wire net742;
 wire net741;
 wire net740;
 wire net739;
 wire net738;
 wire net737;
 wire net736;
 wire net735;
 wire net734;
 wire net733;
 wire net732;
 wire net731;
 wire net730;
 wire net729;
 wire net728;
 wire net727;
 wire net726;
 wire net725;
 wire net724;
 wire net723;
 wire _09236_;
 wire net722;
 wire net721;
 wire net720;
 wire _09240_;
 wire net719;
 wire net718;
 wire net717;
 wire _09244_;
 wire net716;
 wire net715;
 wire net714;
 wire _09248_;
 wire net713;
 wire net712;
 wire net711;
 wire _09252_;
 wire net710;
 wire net709;
 wire net708;
 wire _09256_;
 wire net707;
 wire net706;
 wire net705;
 wire _09260_;
 wire net704;
 wire net703;
 wire net702;
 wire _09264_;
 wire net452;
 wire net451;
 wire net450;
 wire _09268_;
 wire net449;
 wire net448;
 wire net447;
 wire _09272_;
 wire net446;
 wire net445;
 wire net444;
 wire _09276_;
 wire net443;
 wire net442;
 wire net441;
 wire _09280_;
 wire net440;
 wire net439;
 wire net438;
 wire _09284_;
 wire net437;
 wire net436;
 wire net435;
 wire _09288_;
 wire net434;
 wire net433;
 wire net432;
 wire _09292_;
 wire net431;
 wire net430;
 wire net429;
 wire _09296_;
 wire net428;
 wire net427;
 wire net426;
 wire _09300_;
 wire net425;
 wire net424;
 wire net423;
 wire _09304_;
 wire net422;
 wire net421;
 wire net420;
 wire net419;
 wire _09309_;
 wire net418;
 wire net417;
 wire net416;
 wire _09313_;
 wire net415;
 wire net414;
 wire net413;
 wire _09317_;
 wire net412;
 wire net411;
 wire net410;
 wire _09321_;
 wire net409;
 wire net408;
 wire net407;
 wire _09325_;
 wire net406;
 wire net405;
 wire net404;
 wire _09329_;
 wire net403;
 wire net402;
 wire net401;
 wire _09333_;
 wire net400;
 wire net399;
 wire net398;
 wire _09337_;
 wire net397;
 wire net396;
 wire net395;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire net394;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire net393;
 wire net392;
 wire net391;
 wire net390;
 wire net389;
 wire net388;
 wire net387;
 wire net386;
 wire net385;
 wire net384;
 wire net383;
 wire net382;
 wire net381;
 wire net380;
 wire net379;
 wire _09889_;
 wire _09890_;
 wire net378;
 wire net377;
 wire _09893_;
 wire net375;
 wire net374;
 wire net373;
 wire _09897_;
 wire _09898_;
 wire net372;
 wire net371;
 wire _09901_;
 wire _09902_;
 wire net370;
 wire _09904_;
 wire net369;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire net368;
 wire net367;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire net366;
 wire _09928_;
 wire _09929_;
 wire net365;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire net364;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire net363;
 wire _09942_;
 wire net362;
 wire net361;
 wire net360;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire net359;
 wire net358;
 wire _09951_;
 wire net357;
 wire _09953_;
 wire net356;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire net355;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire net354;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire net353;
 wire _09997_;
 wire net352;
 wire net351;
 wire net350;
 wire net349;
 wire net348;
 wire net347;
 wire _10004_;
 wire net346;
 wire net345;
 wire _10007_;
 wire _10008_;
 wire net344;
 wire net343;
 wire _10011_;
 wire net342;
 wire _10013_;
 wire net341;
 wire _10015_;
 wire _10016_;
 wire net340;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire net339;
 wire net338;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire net337;
 wire net336;
 wire _10030_;
 wire net335;
 wire net334;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire net333;
 wire net332;
 wire net331;
 wire net330;
 wire _10040_;
 wire net329;
 wire net328;
 wire net327;
 wire net326;
 wire _10045_;
 wire net325;
 wire net324;
 wire _10048_;
 wire net323;
 wire net322;
 wire _10051_;
 wire net321;
 wire net320;
 wire _10054_;
 wire net319;
 wire net318;
 wire net317;
 wire _10058_;
 wire net316;
 wire net315;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire net314;
 wire net313;
 wire _10066_;
 wire net312;
 wire net311;
 wire _10069_;
 wire net310;
 wire _10071_;
 wire _10072_;
 wire net309;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire net308;
 wire net307;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire net306;
 wire net305;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire net304;
 wire net303;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire net302;
 wire net301;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire net300;
 wire net299;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire net298;
 wire net297;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire net296;
 wire _10158_;
 wire net295;
 wire net294;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire net293;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire net292;
 wire net291;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire net290;
 wire net289;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire net288;
 wire net287;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire net286;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire net285;
 wire net284;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire net283;
 wire net282;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire net281;
 wire net280;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire net279;
 wire net278;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire net277;
 wire net276;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire net275;
 wire net274;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire net273;
 wire _10301_;
 wire net272;
 wire net271;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire net270;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire net269;
 wire net268;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire net267;
 wire net266;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire net265;
 wire net264;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire net263;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire net262;
 wire net261;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire net260;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire net259;
 wire net258;
 wire net257;
 wire net256;
 wire net255;
 wire net254;
 wire net253;
 wire _10490_;
 wire net252;
 wire net251;
 wire _10493_;
 wire _10494_;
 wire net250;
 wire net249;
 wire net248;
 wire _10498_;
 wire _10499_;
 wire net247;
 wire net246;
 wire _10502_;
 wire _10503_;
 wire net245;
 wire net244;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire net243;
 wire net242;
 wire net241;
 wire _10512_;
 wire _10513_;
 wire net240;
 wire net239;
 wire net238;
 wire net237;
 wire net236;
 wire net235;
 wire net234;
 wire _10521_;
 wire _10522_;
 wire net233;
 wire net232;
 wire net231;
 wire net230;
 wire net229;
 wire net228;
 wire net227;
 wire net226;
 wire _10531_;
 wire _10532_;
 wire net225;
 wire net224;
 wire _10535_;
 wire _10536_;
 wire net223;
 wire net222;
 wire net221;
 wire _10540_;
 wire _10541_;
 wire net220;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire net219;
 wire _10552_;
 wire _10553_;
 wire net218;
 wire net217;
 wire _10556_;
 wire net216;
 wire _10558_;
 wire net215;
 wire _10560_;
 wire _10561_;
 wire net214;
 wire _10563_;
 wire _10564_;
 wire net213;
 wire net212;
 wire net211;
 wire _10568_;
 wire _10569_;
 wire net210;
 wire _10571_;
 wire net209;
 wire _10573_;
 wire net208;
 wire _10575_;
 wire net207;
 wire net206;
 wire net205;
 wire net204;
 wire _10580_;
 wire net203;
 wire net202;
 wire _10583_;
 wire net201;
 wire _10585_;
 wire net200;
 wire net199;
 wire net198;
 wire net197;
 wire _10590_;
 wire net196;
 wire net195;
 wire net194;
 wire _10594_;
 wire _10595_;
 wire net193;
 wire net192;
 wire net191;
 wire _10599_;
 wire _10600_;
 wire net190;
 wire _10602_;
 wire net189;
 wire _10604_;
 wire net188;
 wire net187;
 wire net186;
 wire net185;
 wire _10609_;
 wire net184;
 wire net183;
 wire net182;
 wire _10613_;
 wire _10614_;
 wire net181;
 wire _10616_;
 wire _10617_;
 wire net180;
 wire _10619_;
 wire net179;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire net178;
 wire _10625_;
 wire _10626_;
 wire net177;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire net176;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire net175;
 wire _10645_;
 wire net174;
 wire _10647_;
 wire _10648_;
 wire net173;
 wire net172;
 wire _10651_;
 wire net171;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire net170;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire net169;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire net168;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire net167;
 wire _10712_;
 wire _10713_;
 wire net166;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire net165;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire net164;
 wire _10754_;
 wire net163;
 wire net162;
 wire _10757_;
 wire net161;
 wire _10759_;
 wire net160;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire net159;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire net158;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire net157;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire net156;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire net155;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire net154;
 wire _10835_;
 wire _10836_;
 wire net153;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire net152;
 wire _10845_;
 wire _10846_;
 wire net151;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire net150;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire net149;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire net148;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire net147;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire net146;
 wire net145;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire net144;
 wire net143;
 wire net142;
 wire net141;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire net136;
 wire _11155_;
 wire net135;
 wire net134;
 wire net133;
 wire net132;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire net131;
 wire net130;
 wire net129;
 wire net128;
 wire net127;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire net126;
 wire net125;
 wire _11176_;
 wire net124;
 wire net123;
 wire net122;
 wire _11180_;
 wire net121;
 wire net120;
 wire _11183_;
 wire net119;
 wire net118;
 wire _11186_;
 wire net117;
 wire net116;
 wire _11189_;
 wire net115;
 wire net114;
 wire _11192_;
 wire net113;
 wire _11194_;
 wire net112;
 wire net111;
 wire _11197_;
 wire net110;
 wire net109;
 wire _11200_;
 wire net108;
 wire net107;
 wire _11203_;
 wire net106;
 wire net105;
 wire _11206_;
 wire net104;
 wire _11208_;
 wire net103;
 wire net102;
 wire _11211_;
 wire net101;
 wire _11213_;
 wire net100;
 wire net99;
 wire _11216_;
 wire _11217_;
 wire net98;
 wire _11219_;
 wire net97;
 wire net96;
 wire _11222_;
 wire net95;
 wire net94;
 wire _11225_;
 wire net93;
 wire _11227_;
 wire net92;
 wire net91;
 wire _11230_;
 wire net90;
 wire net89;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire net88;
 wire _11250_;
 wire _11251_;
 wire net87;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire net86;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire _11283_;
 wire net75;
 wire net74;
 wire _11286_;
 wire _11287_;
 wire net73;
 wire net72;
 wire _11290_;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire _11296_;
 wire _11297_;
 wire net66;
 wire net65;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire net64;
 wire net63;
 wire _11306_;
 wire net62;
 wire net61;
 wire net60;
 wire _11310_;
 wire net59;
 wire net58;
 wire _11313_;
 wire net57;
 wire net56;
 wire _11316_;
 wire net55;
 wire net54;
 wire _11319_;
 wire net53;
 wire net52;
 wire _11322_;
 wire net51;
 wire net50;
 wire _11325_;
 wire net49;
 wire _11327_;
 wire net48;
 wire net47;
 wire _11330_;
 wire net46;
 wire net45;
 wire _11333_;
 wire net44;
 wire net43;
 wire _11336_;
 wire net42;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire net41;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire net40;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire net39;
 wire _11399_;
 wire _11400_;
 wire net38;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire net37;
 wire _11410_;
 wire _11411_;
 wire net36;
 wire _11413_;
 wire net35;
 wire _11415_;
 wire _11416_;
 wire net34;
 wire net33;
 wire _11419_;
 wire net32;
 wire net31;
 wire _11422_;
 wire _11423_;
 wire net30;
 wire net29;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire net28;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire net27;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire net26;
 wire net25;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire net24;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire net23;
 wire net22;
 wire _11479_;
 wire _11480_;
 wire net21;
 wire _11482_;
 wire net20;
 wire _11484_;
 wire net19;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire net18;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire net17;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire net16;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire net15;
 wire _11555_;
 wire _11556_;
 wire net14;
 wire net13;
 wire _11559_;
 wire net12;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire net11;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire clknet_leaf_138_clk;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire \count15_1[1] ;
 wire \count15_1[2] ;
 wire \count15_1[3] ;
 wire \count15_1[4] ;
 wire \count15_1[5] ;
 wire \count15_2[1] ;
 wire \count15_2[2] ;
 wire \count15_2[3] ;
 wire \count15_2[4] ;
 wire \count15_2[5] ;
 wire \count16_1[1] ;
 wire \count16_1[2] ;
 wire \count16_1[3] ;
 wire \count16_1[4] ;
 wire \count16_1[5] ;
 wire \count16_2[1] ;
 wire \count16_2[2] ;
 wire \count16_2[3] ;
 wire \count16_2[4] ;
 wire \count16_2[5] ;
 wire \count2_1[1] ;
 wire \count2_1[2] ;
 wire \count2_1[3] ;
 wire \count2_1[4] ;
 wire \count2_1[5] ;
 wire \count2_2[1] ;
 wire \count2_2[2] ;
 wire \count2_2[3] ;
 wire \count2_2[4] ;
 wire \count2_2[5] ;
 wire \count7_1[1] ;
 wire \count7_1[2] ;
 wire \count7_1[3] ;
 wire \count7_1[4] ;
 wire \count7_1[5] ;
 wire \count7_2[1] ;
 wire \count7_2[2] ;
 wire \count7_2[3] ;
 wire \count7_2[4] ;
 wire \count7_2[5] ;
 wire \count_1[1] ;
 wire \count_1[2] ;
 wire \count_1[3] ;
 wire \count_1[4] ;
 wire \count_1[5] ;
 wire \count_2[1] ;
 wire \count_2[2] ;
 wire \count_2[3] ;
 wire \count_2[4] ;
 wire \count_2[5] ;
 wire \count_2[6] ;
 wire \count_hash1[1] ;
 wire \count_hash1[2] ;
 wire \count_hash1[3] ;
 wire \count_hash1[4] ;
 wire \count_hash1[5] ;
 wire \count_hash1[6] ;
 wire \count_hash2[1] ;
 wire \count_hash2[2] ;
 wire \count_hash2[3] ;
 wire \count_hash2[4] ;
 wire \count_hash2[5] ;
 wire done;
 wire \hash.CA1.S0.X[0] ;
 wire \hash.CA1.S0.X[10] ;
 wire \hash.CA1.S0.X[11] ;
 wire \hash.CA1.S0.X[12] ;
 wire \hash.CA1.S0.X[13] ;
 wire \hash.CA1.S0.X[14] ;
 wire \hash.CA1.S0.X[15] ;
 wire \hash.CA1.S0.X[16] ;
 wire \hash.CA1.S0.X[17] ;
 wire clknet_leaf_159_clk;
 wire \hash.CA1.S0.X[19] ;
 wire \hash.CA1.S0.X[1] ;
 wire \hash.CA1.S0.X[20] ;
 wire clknet_leaf_156_clk;
 wire \hash.CA1.S0.X[22] ;
 wire \hash.CA1.S0.X[23] ;
 wire \hash.CA1.S0.X[24] ;
 wire \hash.CA1.S0.X[25] ;
 wire \hash.CA1.S0.X[26] ;
 wire \hash.CA1.S0.X[27] ;
 wire \hash.CA1.S0.X[28] ;
 wire \hash.CA1.S0.X[29] ;
 wire \hash.CA1.S0.X[2] ;
 wire \hash.CA1.S0.X[30] ;
 wire \hash.CA1.S0.X[31] ;
 wire \hash.CA1.S0.X[3] ;
 wire \hash.CA1.S0.X[4] ;
 wire \hash.CA1.S0.X[5] ;
 wire \hash.CA1.S0.X[6] ;
 wire \hash.CA1.S0.X[7] ;
 wire \hash.CA1.S0.X[8] ;
 wire \hash.CA1.S0.X[9] ;
 wire \hash.CA1.S1.X[0] ;
 wire \hash.CA1.S1.X[10] ;
 wire \hash.CA1.S1.X[11] ;
 wire \hash.CA1.S1.X[12] ;
 wire \hash.CA1.S1.X[13] ;
 wire \hash.CA1.S1.X[14] ;
 wire \hash.CA1.S1.X[15] ;
 wire clknet_leaf_110_clk;
 wire \hash.CA1.S1.X[17] ;
 wire \hash.CA1.S1.X[18] ;
 wire \hash.CA1.S1.X[19] ;
 wire \hash.CA1.S1.X[1] ;
 wire \hash.CA1.S1.X[20] ;
 wire \hash.CA1.S1.X[21] ;
 wire clknet_leaf_109_clk;
 wire \hash.CA1.S1.X[23] ;
 wire \hash.CA1.S1.X[24] ;
 wire \hash.CA1.S1.X[25] ;
 wire \hash.CA1.S1.X[26] ;
 wire \hash.CA1.S1.X[27] ;
 wire \hash.CA1.S1.X[28] ;
 wire \hash.CA1.S1.X[29] ;
 wire \hash.CA1.S1.X[2] ;
 wire \hash.CA1.S1.X[30] ;
 wire clknet_leaf_106_clk;
 wire \hash.CA1.S1.X[3] ;
 wire \hash.CA1.S1.X[4] ;
 wire \hash.CA1.S1.X[5] ;
 wire \hash.CA1.S1.X[6] ;
 wire \hash.CA1.S1.X[7] ;
 wire \hash.CA1.S1.X[8] ;
 wire \hash.CA1.S1.X[9] ;
 wire \hash.CA1.b[0] ;
 wire \hash.CA1.b[10] ;
 wire \hash.CA1.b[11] ;
 wire \hash.CA1.b[12] ;
 wire \hash.CA1.b[13] ;
 wire \hash.CA1.b[14] ;
 wire \hash.CA1.b[15] ;
 wire \hash.CA1.b[16] ;
 wire \hash.CA1.b[17] ;
 wire \hash.CA1.b[18] ;
 wire \hash.CA1.b[19] ;
 wire \hash.CA1.b[1] ;
 wire \hash.CA1.b[20] ;
 wire clknet_leaf_140_clk;
 wire \hash.CA1.b[22] ;
 wire clknet_leaf_139_clk;
 wire \hash.CA1.b[24] ;
 wire \hash.CA1.b[25] ;
 wire \hash.CA1.b[26] ;
 wire clknet_leaf_137_clk;
 wire \hash.CA1.b[28] ;
 wire \hash.CA1.b[29] ;
 wire \hash.CA1.b[2] ;
 wire \hash.CA1.b[30] ;
 wire \hash.CA1.b[31] ;
 wire \hash.CA1.b[3] ;
 wire \hash.CA1.b[4] ;
 wire \hash.CA1.b[5] ;
 wire \hash.CA1.b[6] ;
 wire \hash.CA1.b[7] ;
 wire \hash.CA1.b[8] ;
 wire \hash.CA1.b[9] ;
 wire \hash.CA1.c[0] ;
 wire \hash.CA1.d[0] ;
 wire \hash.CA1.f[0] ;
 wire \hash.CA1.f[10] ;
 wire \hash.CA1.f[11] ;
 wire \hash.CA1.f[12] ;
 wire \hash.CA1.f[13] ;
 wire \hash.CA1.f[14] ;
 wire \hash.CA1.f[15] ;
 wire \hash.CA1.f[16] ;
 wire \hash.CA1.f[17] ;
 wire \hash.CA1.f[18] ;
 wire \hash.CA1.f[19] ;
 wire \hash.CA1.f[1] ;
 wire \hash.CA1.f[20] ;
 wire \hash.CA1.f[21] ;
 wire \hash.CA1.f[22] ;
 wire \hash.CA1.f[23] ;
 wire clknet_leaf_116_clk;
 wire \hash.CA1.f[25] ;
 wire \hash.CA1.f[26] ;
 wire \hash.CA1.f[27] ;
 wire \hash.CA1.f[28] ;
 wire \hash.CA1.f[29] ;
 wire \hash.CA1.f[2] ;
 wire \hash.CA1.f[30] ;
 wire \hash.CA1.f[31] ;
 wire \hash.CA1.f[3] ;
 wire \hash.CA1.f[4] ;
 wire \hash.CA1.f[5] ;
 wire \hash.CA1.f[6] ;
 wire \hash.CA1.f[7] ;
 wire \hash.CA1.f[8] ;
 wire \hash.CA1.f[9] ;
 wire \hash.CA1.k_i1[0] ;
 wire \hash.CA1.k_i1[10] ;
 wire \hash.CA1.k_i1[11] ;
 wire \hash.CA1.k_i1[12] ;
 wire \hash.CA1.k_i1[13] ;
 wire \hash.CA1.k_i1[14] ;
 wire \hash.CA1.k_i1[15] ;
 wire \hash.CA1.k_i1[16] ;
 wire \hash.CA1.k_i1[17] ;
 wire \hash.CA1.k_i1[18] ;
 wire \hash.CA1.k_i1[19] ;
 wire \hash.CA1.k_i1[1] ;
 wire \hash.CA1.k_i1[20] ;
 wire \hash.CA1.k_i1[21] ;
 wire \hash.CA1.k_i1[22] ;
 wire \hash.CA1.k_i1[23] ;
 wire \hash.CA1.k_i1[24] ;
 wire \hash.CA1.k_i1[25] ;
 wire \hash.CA1.k_i1[26] ;
 wire \hash.CA1.k_i1[27] ;
 wire \hash.CA1.k_i1[28] ;
 wire \hash.CA1.k_i1[29] ;
 wire \hash.CA1.k_i1[2] ;
 wire \hash.CA1.k_i1[30] ;
 wire \hash.CA1.k_i1[31] ;
 wire \hash.CA1.k_i1[3] ;
 wire \hash.CA1.k_i1[4] ;
 wire \hash.CA1.k_i1[5] ;
 wire \hash.CA1.k_i1[6] ;
 wire \hash.CA1.k_i1[7] ;
 wire \hash.CA1.k_i1[8] ;
 wire \hash.CA1.k_i1[9] ;
 wire \hash.CA1.k_i2[0] ;
 wire \hash.CA1.k_i2[10] ;
 wire \hash.CA1.k_i2[11] ;
 wire \hash.CA1.k_i2[12] ;
 wire \hash.CA1.k_i2[13] ;
 wire \hash.CA1.k_i2[14] ;
 wire \hash.CA1.k_i2[15] ;
 wire \hash.CA1.k_i2[16] ;
 wire \hash.CA1.k_i2[17] ;
 wire \hash.CA1.k_i2[18] ;
 wire \hash.CA1.k_i2[19] ;
 wire \hash.CA1.k_i2[1] ;
 wire \hash.CA1.k_i2[20] ;
 wire \hash.CA1.k_i2[21] ;
 wire \hash.CA1.k_i2[22] ;
 wire \hash.CA1.k_i2[23] ;
 wire \hash.CA1.k_i2[24] ;
 wire \hash.CA1.k_i2[25] ;
 wire \hash.CA1.k_i2[26] ;
 wire \hash.CA1.k_i2[27] ;
 wire \hash.CA1.k_i2[28] ;
 wire \hash.CA1.k_i2[29] ;
 wire \hash.CA1.k_i2[2] ;
 wire \hash.CA1.k_i2[30] ;
 wire \hash.CA1.k_i2[31] ;
 wire \hash.CA1.k_i2[3] ;
 wire \hash.CA1.k_i2[4] ;
 wire \hash.CA1.k_i2[5] ;
 wire \hash.CA1.k_i2[6] ;
 wire \hash.CA1.k_i2[7] ;
 wire \hash.CA1.k_i2[8] ;
 wire \hash.CA1.k_i2[9] ;
 wire \hash.CA1.p1[0] ;
 wire \hash.CA1.p1[10] ;
 wire \hash.CA1.p1[11] ;
 wire \hash.CA1.p1[12] ;
 wire \hash.CA1.p1[13] ;
 wire \hash.CA1.p1[14] ;
 wire \hash.CA1.p1[15] ;
 wire \hash.CA1.p1[16] ;
 wire \hash.CA1.p1[17] ;
 wire \hash.CA1.p1[18] ;
 wire \hash.CA1.p1[19] ;
 wire \hash.CA1.p1[1] ;
 wire \hash.CA1.p1[20] ;
 wire \hash.CA1.p1[21] ;
 wire \hash.CA1.p1[22] ;
 wire \hash.CA1.p1[23] ;
 wire \hash.CA1.p1[24] ;
 wire \hash.CA1.p1[25] ;
 wire \hash.CA1.p1[26] ;
 wire \hash.CA1.p1[27] ;
 wire \hash.CA1.p1[28] ;
 wire \hash.CA1.p1[29] ;
 wire \hash.CA1.p1[2] ;
 wire \hash.CA1.p1[30] ;
 wire \hash.CA1.p1[31] ;
 wire \hash.CA1.p1[3] ;
 wire \hash.CA1.p1[4] ;
 wire \hash.CA1.p1[5] ;
 wire \hash.CA1.p1[6] ;
 wire \hash.CA1.p1[7] ;
 wire \hash.CA1.p1[8] ;
 wire \hash.CA1.p1[9] ;
 wire \hash.CA1.p2[0] ;
 wire \hash.CA1.p2[10] ;
 wire \hash.CA1.p2[11] ;
 wire \hash.CA1.p2[12] ;
 wire \hash.CA1.p2[13] ;
 wire \hash.CA1.p2[14] ;
 wire \hash.CA1.p2[15] ;
 wire \hash.CA1.p2[16] ;
 wire \hash.CA1.p2[17] ;
 wire \hash.CA1.p2[18] ;
 wire \hash.CA1.p2[19] ;
 wire \hash.CA1.p2[1] ;
 wire \hash.CA1.p2[20] ;
 wire \hash.CA1.p2[21] ;
 wire \hash.CA1.p2[22] ;
 wire \hash.CA1.p2[23] ;
 wire \hash.CA1.p2[24] ;
 wire \hash.CA1.p2[25] ;
 wire \hash.CA1.p2[26] ;
 wire \hash.CA1.p2[27] ;
 wire \hash.CA1.p2[28] ;
 wire \hash.CA1.p2[29] ;
 wire \hash.CA1.p2[2] ;
 wire \hash.CA1.p2[30] ;
 wire \hash.CA1.p2[31] ;
 wire \hash.CA1.p2[3] ;
 wire \hash.CA1.p2[4] ;
 wire \hash.CA1.p2[5] ;
 wire \hash.CA1.p2[6] ;
 wire \hash.CA1.p2[7] ;
 wire \hash.CA1.p2[8] ;
 wire \hash.CA1.p2[9] ;
 wire \hash.CA1.p3[0] ;
 wire \hash.CA1.p3[10] ;
 wire \hash.CA1.p3[11] ;
 wire \hash.CA1.p3[12] ;
 wire \hash.CA1.p3[13] ;
 wire \hash.CA1.p3[14] ;
 wire \hash.CA1.p3[15] ;
 wire \hash.CA1.p3[16] ;
 wire \hash.CA1.p3[17] ;
 wire \hash.CA1.p3[18] ;
 wire \hash.CA1.p3[19] ;
 wire \hash.CA1.p3[1] ;
 wire \hash.CA1.p3[20] ;
 wire \hash.CA1.p3[21] ;
 wire \hash.CA1.p3[22] ;
 wire \hash.CA1.p3[23] ;
 wire \hash.CA1.p3[24] ;
 wire \hash.CA1.p3[25] ;
 wire \hash.CA1.p3[26] ;
 wire \hash.CA1.p3[27] ;
 wire \hash.CA1.p3[28] ;
 wire \hash.CA1.p3[29] ;
 wire \hash.CA1.p3[2] ;
 wire \hash.CA1.p3[30] ;
 wire \hash.CA1.p3[31] ;
 wire \hash.CA1.p3[3] ;
 wire \hash.CA1.p3[4] ;
 wire \hash.CA1.p3[5] ;
 wire \hash.CA1.p3[6] ;
 wire \hash.CA1.p3[7] ;
 wire \hash.CA1.p3[8] ;
 wire \hash.CA1.p3[9] ;
 wire \hash.CA1.p4[0] ;
 wire \hash.CA1.p4[10] ;
 wire \hash.CA1.p4[11] ;
 wire \hash.CA1.p4[12] ;
 wire \hash.CA1.p4[13] ;
 wire \hash.CA1.p4[14] ;
 wire \hash.CA1.p4[15] ;
 wire \hash.CA1.p4[16] ;
 wire \hash.CA1.p4[17] ;
 wire \hash.CA1.p4[18] ;
 wire \hash.CA1.p4[19] ;
 wire \hash.CA1.p4[1] ;
 wire \hash.CA1.p4[20] ;
 wire \hash.CA1.p4[21] ;
 wire \hash.CA1.p4[22] ;
 wire \hash.CA1.p4[23] ;
 wire \hash.CA1.p4[24] ;
 wire \hash.CA1.p4[25] ;
 wire \hash.CA1.p4[26] ;
 wire \hash.CA1.p4[27] ;
 wire \hash.CA1.p4[28] ;
 wire \hash.CA1.p4[29] ;
 wire \hash.CA1.p4[2] ;
 wire \hash.CA1.p4[30] ;
 wire \hash.CA1.p4[31] ;
 wire \hash.CA1.p4[3] ;
 wire \hash.CA1.p4[4] ;
 wire \hash.CA1.p4[5] ;
 wire \hash.CA1.p4[6] ;
 wire \hash.CA1.p4[7] ;
 wire \hash.CA1.p4[8] ;
 wire \hash.CA1.p4[9] ;
 wire \hash.CA1.p5[0] ;
 wire \hash.CA1.p5[10] ;
 wire \hash.CA1.p5[11] ;
 wire \hash.CA1.p5[12] ;
 wire \hash.CA1.p5[13] ;
 wire \hash.CA1.p5[14] ;
 wire \hash.CA1.p5[15] ;
 wire \hash.CA1.p5[16] ;
 wire \hash.CA1.p5[17] ;
 wire \hash.CA1.p5[18] ;
 wire \hash.CA1.p5[19] ;
 wire \hash.CA1.p5[1] ;
 wire \hash.CA1.p5[20] ;
 wire \hash.CA1.p5[21] ;
 wire \hash.CA1.p5[22] ;
 wire \hash.CA1.p5[23] ;
 wire \hash.CA1.p5[24] ;
 wire \hash.CA1.p5[25] ;
 wire \hash.CA1.p5[26] ;
 wire \hash.CA1.p5[27] ;
 wire \hash.CA1.p5[28] ;
 wire \hash.CA1.p5[29] ;
 wire \hash.CA1.p5[2] ;
 wire \hash.CA1.p5[30] ;
 wire \hash.CA1.p5[31] ;
 wire \hash.CA1.p5[3] ;
 wire \hash.CA1.p5[4] ;
 wire \hash.CA1.p5[5] ;
 wire \hash.CA1.p5[6] ;
 wire \hash.CA1.p5[7] ;
 wire \hash.CA1.p5[8] ;
 wire \hash.CA1.p5[9] ;
 wire \hash.CA1.w_i1[0] ;
 wire \hash.CA1.w_i1[10] ;
 wire \hash.CA1.w_i1[11] ;
 wire \hash.CA1.w_i1[12] ;
 wire \hash.CA1.w_i1[13] ;
 wire \hash.CA1.w_i1[14] ;
 wire \hash.CA1.w_i1[15] ;
 wire \hash.CA1.w_i1[16] ;
 wire \hash.CA1.w_i1[17] ;
 wire \hash.CA1.w_i1[18] ;
 wire \hash.CA1.w_i1[19] ;
 wire \hash.CA1.w_i1[1] ;
 wire \hash.CA1.w_i1[20] ;
 wire \hash.CA1.w_i1[21] ;
 wire \hash.CA1.w_i1[22] ;
 wire \hash.CA1.w_i1[23] ;
 wire \hash.CA1.w_i1[24] ;
 wire \hash.CA1.w_i1[25] ;
 wire \hash.CA1.w_i1[26] ;
 wire \hash.CA1.w_i1[27] ;
 wire \hash.CA1.w_i1[28] ;
 wire \hash.CA1.w_i1[29] ;
 wire \hash.CA1.w_i1[2] ;
 wire \hash.CA1.w_i1[30] ;
 wire \hash.CA1.w_i1[31] ;
 wire \hash.CA1.w_i1[3] ;
 wire \hash.CA1.w_i1[4] ;
 wire \hash.CA1.w_i1[5] ;
 wire \hash.CA1.w_i1[6] ;
 wire \hash.CA1.w_i1[7] ;
 wire \hash.CA1.w_i1[8] ;
 wire \hash.CA1.w_i1[9] ;
 wire \hash.CA1.w_i2[0] ;
 wire \hash.CA1.w_i2[10] ;
 wire \hash.CA1.w_i2[11] ;
 wire \hash.CA1.w_i2[12] ;
 wire \hash.CA1.w_i2[13] ;
 wire \hash.CA1.w_i2[14] ;
 wire \hash.CA1.w_i2[15] ;
 wire \hash.CA1.w_i2[16] ;
 wire \hash.CA1.w_i2[17] ;
 wire \hash.CA1.w_i2[18] ;
 wire \hash.CA1.w_i2[19] ;
 wire \hash.CA1.w_i2[1] ;
 wire \hash.CA1.w_i2[20] ;
 wire \hash.CA1.w_i2[21] ;
 wire \hash.CA1.w_i2[22] ;
 wire \hash.CA1.w_i2[23] ;
 wire \hash.CA1.w_i2[24] ;
 wire \hash.CA1.w_i2[25] ;
 wire \hash.CA1.w_i2[26] ;
 wire \hash.CA1.w_i2[27] ;
 wire \hash.CA1.w_i2[28] ;
 wire \hash.CA1.w_i2[29] ;
 wire \hash.CA1.w_i2[2] ;
 wire \hash.CA1.w_i2[30] ;
 wire \hash.CA1.w_i2[31] ;
 wire \hash.CA1.w_i2[3] ;
 wire \hash.CA1.w_i2[4] ;
 wire \hash.CA1.w_i2[5] ;
 wire \hash.CA1.w_i2[6] ;
 wire \hash.CA1.w_i2[7] ;
 wire \hash.CA1.w_i2[8] ;
 wire \hash.CA1.w_i2[9] ;
 wire \hash.CA2.S1.X[0] ;
 wire \hash.CA2.S1.X[10] ;
 wire \hash.CA2.S1.X[11] ;
 wire \hash.CA2.S1.X[12] ;
 wire \hash.CA2.S1.X[13] ;
 wire \hash.CA2.S1.X[14] ;
 wire \hash.CA2.S1.X[15] ;
 wire \hash.CA2.S1.X[16] ;
 wire \hash.CA2.S1.X[17] ;
 wire \hash.CA2.S1.X[18] ;
 wire \hash.CA2.S1.X[19] ;
 wire \hash.CA2.S1.X[1] ;
 wire \hash.CA2.S1.X[20] ;
 wire \hash.CA2.S1.X[21] ;
 wire \hash.CA2.S1.X[22] ;
 wire \hash.CA2.S1.X[23] ;
 wire \hash.CA2.S1.X[24] ;
 wire \hash.CA2.S1.X[25] ;
 wire \hash.CA2.S1.X[26] ;
 wire \hash.CA2.S1.X[27] ;
 wire \hash.CA2.S1.X[28] ;
 wire \hash.CA2.S1.X[29] ;
 wire \hash.CA2.S1.X[2] ;
 wire \hash.CA2.S1.X[30] ;
 wire \hash.CA2.S1.X[31] ;
 wire \hash.CA2.S1.X[3] ;
 wire \hash.CA2.S1.X[4] ;
 wire \hash.CA2.S1.X[5] ;
 wire \hash.CA2.S1.X[6] ;
 wire \hash.CA2.S1.X[7] ;
 wire \hash.CA2.S1.X[8] ;
 wire \hash.CA2.S1.X[9] ;
 wire \hash.CA2.a_dash[0] ;
 wire \hash.CA2.a_dash[10] ;
 wire \hash.CA2.a_dash[11] ;
 wire \hash.CA2.a_dash[12] ;
 wire \hash.CA2.a_dash[13] ;
 wire \hash.CA2.a_dash[14] ;
 wire \hash.CA2.a_dash[15] ;
 wire \hash.CA2.a_dash[16] ;
 wire \hash.CA2.a_dash[17] ;
 wire \hash.CA2.a_dash[18] ;
 wire \hash.CA2.a_dash[19] ;
 wire \hash.CA2.a_dash[1] ;
 wire \hash.CA2.a_dash[20] ;
 wire \hash.CA2.a_dash[21] ;
 wire \hash.CA2.a_dash[22] ;
 wire \hash.CA2.a_dash[23] ;
 wire \hash.CA2.a_dash[24] ;
 wire \hash.CA2.a_dash[25] ;
 wire \hash.CA2.a_dash[26] ;
 wire \hash.CA2.a_dash[27] ;
 wire \hash.CA2.a_dash[28] ;
 wire \hash.CA2.a_dash[29] ;
 wire \hash.CA2.a_dash[2] ;
 wire \hash.CA2.a_dash[30] ;
 wire \hash.CA2.a_dash[31] ;
 wire \hash.CA2.a_dash[3] ;
 wire \hash.CA2.a_dash[4] ;
 wire \hash.CA2.a_dash[5] ;
 wire \hash.CA2.a_dash[6] ;
 wire \hash.CA2.a_dash[7] ;
 wire \hash.CA2.a_dash[8] ;
 wire \hash.CA2.a_dash[9] ;
 wire \hash.CA2.b_dash[0] ;
 wire \hash.CA2.b_dash[10] ;
 wire \hash.CA2.b_dash[11] ;
 wire \hash.CA2.b_dash[12] ;
 wire \hash.CA2.b_dash[13] ;
 wire \hash.CA2.b_dash[14] ;
 wire \hash.CA2.b_dash[15] ;
 wire \hash.CA2.b_dash[16] ;
 wire \hash.CA2.b_dash[17] ;
 wire \hash.CA2.b_dash[18] ;
 wire \hash.CA2.b_dash[19] ;
 wire \hash.CA2.b_dash[1] ;
 wire \hash.CA2.b_dash[20] ;
 wire \hash.CA2.b_dash[21] ;
 wire \hash.CA2.b_dash[22] ;
 wire \hash.CA2.b_dash[23] ;
 wire \hash.CA2.b_dash[24] ;
 wire \hash.CA2.b_dash[25] ;
 wire \hash.CA2.b_dash[26] ;
 wire \hash.CA2.b_dash[27] ;
 wire \hash.CA2.b_dash[28] ;
 wire \hash.CA2.b_dash[29] ;
 wire \hash.CA2.b_dash[2] ;
 wire \hash.CA2.b_dash[30] ;
 wire \hash.CA2.b_dash[31] ;
 wire \hash.CA2.b_dash[3] ;
 wire \hash.CA2.b_dash[4] ;
 wire \hash.CA2.b_dash[5] ;
 wire \hash.CA2.b_dash[6] ;
 wire \hash.CA2.b_dash[7] ;
 wire \hash.CA2.b_dash[8] ;
 wire \hash.CA2.b_dash[9] ;
 wire \hash.CA2.e_dash[0] ;
 wire \hash.CA2.e_dash[10] ;
 wire \hash.CA2.e_dash[11] ;
 wire \hash.CA2.e_dash[12] ;
 wire \hash.CA2.e_dash[13] ;
 wire \hash.CA2.e_dash[14] ;
 wire \hash.CA2.e_dash[15] ;
 wire \hash.CA2.e_dash[16] ;
 wire \hash.CA2.e_dash[17] ;
 wire \hash.CA2.e_dash[18] ;
 wire \hash.CA2.e_dash[19] ;
 wire \hash.CA2.e_dash[1] ;
 wire \hash.CA2.e_dash[20] ;
 wire \hash.CA2.e_dash[21] ;
 wire \hash.CA2.e_dash[22] ;
 wire \hash.CA2.e_dash[23] ;
 wire \hash.CA2.e_dash[24] ;
 wire \hash.CA2.e_dash[25] ;
 wire \hash.CA2.e_dash[26] ;
 wire \hash.CA2.e_dash[27] ;
 wire \hash.CA2.e_dash[28] ;
 wire \hash.CA2.e_dash[29] ;
 wire \hash.CA2.e_dash[2] ;
 wire \hash.CA2.e_dash[30] ;
 wire \hash.CA2.e_dash[31] ;
 wire \hash.CA2.e_dash[3] ;
 wire \hash.CA2.e_dash[4] ;
 wire \hash.CA2.e_dash[5] ;
 wire \hash.CA2.e_dash[6] ;
 wire \hash.CA2.e_dash[7] ;
 wire \hash.CA2.e_dash[8] ;
 wire \hash.CA2.e_dash[9] ;
 wire \hash.CA2.f_dash[0] ;
 wire \hash.CA2.f_dash[10] ;
 wire \hash.CA2.f_dash[11] ;
 wire \hash.CA2.f_dash[12] ;
 wire \hash.CA2.f_dash[13] ;
 wire \hash.CA2.f_dash[14] ;
 wire \hash.CA2.f_dash[15] ;
 wire \hash.CA2.f_dash[16] ;
 wire \hash.CA2.f_dash[17] ;
 wire \hash.CA2.f_dash[18] ;
 wire \hash.CA2.f_dash[19] ;
 wire \hash.CA2.f_dash[1] ;
 wire \hash.CA2.f_dash[20] ;
 wire \hash.CA2.f_dash[21] ;
 wire \hash.CA2.f_dash[22] ;
 wire \hash.CA2.f_dash[23] ;
 wire \hash.CA2.f_dash[24] ;
 wire \hash.CA2.f_dash[25] ;
 wire \hash.CA2.f_dash[26] ;
 wire \hash.CA2.f_dash[27] ;
 wire \hash.CA2.f_dash[28] ;
 wire \hash.CA2.f_dash[29] ;
 wire \hash.CA2.f_dash[2] ;
 wire \hash.CA2.f_dash[30] ;
 wire \hash.CA2.f_dash[31] ;
 wire \hash.CA2.f_dash[3] ;
 wire \hash.CA2.f_dash[4] ;
 wire \hash.CA2.f_dash[5] ;
 wire \hash.CA2.f_dash[6] ;
 wire \hash.CA2.f_dash[7] ;
 wire \hash.CA2.f_dash[8] ;
 wire \hash.CA2.f_dash[9] ;
 wire \hash.CA2.p1[0] ;
 wire \hash.CA2.p1[10] ;
 wire \hash.CA2.p1[11] ;
 wire \hash.CA2.p1[12] ;
 wire \hash.CA2.p1[13] ;
 wire \hash.CA2.p1[14] ;
 wire \hash.CA2.p1[15] ;
 wire \hash.CA2.p1[16] ;
 wire \hash.CA2.p1[17] ;
 wire \hash.CA2.p1[18] ;
 wire \hash.CA2.p1[19] ;
 wire \hash.CA2.p1[1] ;
 wire \hash.CA2.p1[20] ;
 wire \hash.CA2.p1[21] ;
 wire \hash.CA2.p1[22] ;
 wire \hash.CA2.p1[23] ;
 wire \hash.CA2.p1[24] ;
 wire \hash.CA2.p1[25] ;
 wire \hash.CA2.p1[26] ;
 wire \hash.CA2.p1[27] ;
 wire \hash.CA2.p1[28] ;
 wire \hash.CA2.p1[29] ;
 wire \hash.CA2.p1[2] ;
 wire \hash.CA2.p1[30] ;
 wire \hash.CA2.p1[31] ;
 wire \hash.CA2.p1[3] ;
 wire \hash.CA2.p1[4] ;
 wire \hash.CA2.p1[5] ;
 wire \hash.CA2.p1[6] ;
 wire \hash.CA2.p1[7] ;
 wire \hash.CA2.p1[8] ;
 wire \hash.CA2.p1[9] ;
 wire \hash.CA2.p3[0] ;
 wire \hash.CA2.p3[10] ;
 wire \hash.CA2.p3[11] ;
 wire \hash.CA2.p3[12] ;
 wire \hash.CA2.p3[13] ;
 wire \hash.CA2.p3[14] ;
 wire \hash.CA2.p3[15] ;
 wire \hash.CA2.p3[16] ;
 wire \hash.CA2.p3[17] ;
 wire \hash.CA2.p3[18] ;
 wire \hash.CA2.p3[19] ;
 wire \hash.CA2.p3[1] ;
 wire \hash.CA2.p3[20] ;
 wire \hash.CA2.p3[21] ;
 wire \hash.CA2.p3[22] ;
 wire \hash.CA2.p3[23] ;
 wire \hash.CA2.p3[24] ;
 wire \hash.CA2.p3[25] ;
 wire \hash.CA2.p3[26] ;
 wire \hash.CA2.p3[27] ;
 wire \hash.CA2.p3[28] ;
 wire \hash.CA2.p3[29] ;
 wire \hash.CA2.p3[2] ;
 wire \hash.CA2.p3[30] ;
 wire \hash.CA2.p3[31] ;
 wire \hash.CA2.p3[3] ;
 wire \hash.CA2.p3[4] ;
 wire \hash.CA2.p3[5] ;
 wire \hash.CA2.p3[6] ;
 wire \hash.CA2.p3[7] ;
 wire \hash.CA2.p3[8] ;
 wire \hash.CA2.p3[9] ;
 wire \hash.CA2.p4[0] ;
 wire \hash.CA2.p4[10] ;
 wire \hash.CA2.p4[11] ;
 wire \hash.CA2.p4[12] ;
 wire \hash.CA2.p4[13] ;
 wire \hash.CA2.p4[14] ;
 wire \hash.CA2.p4[15] ;
 wire \hash.CA2.p4[16] ;
 wire \hash.CA2.p4[17] ;
 wire \hash.CA2.p4[18] ;
 wire \hash.CA2.p4[19] ;
 wire \hash.CA2.p4[1] ;
 wire \hash.CA2.p4[20] ;
 wire \hash.CA2.p4[21] ;
 wire \hash.CA2.p4[22] ;
 wire \hash.CA2.p4[23] ;
 wire \hash.CA2.p4[24] ;
 wire \hash.CA2.p4[25] ;
 wire \hash.CA2.p4[26] ;
 wire \hash.CA2.p4[27] ;
 wire \hash.CA2.p4[28] ;
 wire \hash.CA2.p4[29] ;
 wire \hash.CA2.p4[2] ;
 wire \hash.CA2.p4[30] ;
 wire \hash.CA2.p4[31] ;
 wire \hash.CA2.p4[3] ;
 wire \hash.CA2.p4[4] ;
 wire \hash.CA2.p4[5] ;
 wire \hash.CA2.p4[6] ;
 wire \hash.CA2.p4[7] ;
 wire \hash.CA2.p4[8] ;
 wire \hash.CA2.p4[9] ;
 wire \hash.CA2.p5[0] ;
 wire \hash.CA2.p5[10] ;
 wire \hash.CA2.p5[11] ;
 wire \hash.CA2.p5[12] ;
 wire \hash.CA2.p5[13] ;
 wire \hash.CA2.p5[14] ;
 wire \hash.CA2.p5[15] ;
 wire \hash.CA2.p5[16] ;
 wire \hash.CA2.p5[17] ;
 wire \hash.CA2.p5[18] ;
 wire \hash.CA2.p5[19] ;
 wire \hash.CA2.p5[1] ;
 wire \hash.CA2.p5[20] ;
 wire \hash.CA2.p5[21] ;
 wire \hash.CA2.p5[22] ;
 wire \hash.CA2.p5[23] ;
 wire \hash.CA2.p5[24] ;
 wire \hash.CA2.p5[25] ;
 wire \hash.CA2.p5[26] ;
 wire \hash.CA2.p5[27] ;
 wire \hash.CA2.p5[28] ;
 wire \hash.CA2.p5[29] ;
 wire \hash.CA2.p5[2] ;
 wire \hash.CA2.p5[30] ;
 wire \hash.CA2.p5[31] ;
 wire \hash.CA2.p5[3] ;
 wire \hash.CA2.p5[4] ;
 wire \hash.CA2.p5[5] ;
 wire \hash.CA2.p5[6] ;
 wire \hash.CA2.p5[7] ;
 wire \hash.CA2.p5[8] ;
 wire \hash.CA2.p5[9] ;
 wire \hash.reset ;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire ready_dash;
 wire reset_hash;
 wire \w[0][0] ;
 wire \w[0][10] ;
 wire \w[0][11] ;
 wire \w[0][12] ;
 wire \w[0][13] ;
 wire \w[0][14] ;
 wire \w[0][15] ;
 wire \w[0][16] ;
 wire \w[0][17] ;
 wire \w[0][18] ;
 wire \w[0][19] ;
 wire \w[0][1] ;
 wire \w[0][20] ;
 wire \w[0][21] ;
 wire \w[0][22] ;
 wire \w[0][23] ;
 wire \w[0][24] ;
 wire \w[0][25] ;
 wire \w[0][26] ;
 wire \w[0][27] ;
 wire \w[0][28] ;
 wire \w[0][29] ;
 wire \w[0][2] ;
 wire \w[0][30] ;
 wire \w[0][31] ;
 wire \w[0][3] ;
 wire \w[0][4] ;
 wire \w[0][5] ;
 wire \w[0][6] ;
 wire \w[0][7] ;
 wire \w[0][8] ;
 wire \w[0][9] ;
 wire \w[10][0] ;
 wire \w[10][10] ;
 wire \w[10][11] ;
 wire \w[10][12] ;
 wire \w[10][13] ;
 wire \w[10][14] ;
 wire \w[10][15] ;
 wire \w[10][16] ;
 wire \w[10][17] ;
 wire \w[10][18] ;
 wire \w[10][19] ;
 wire \w[10][1] ;
 wire \w[10][20] ;
 wire \w[10][21] ;
 wire \w[10][22] ;
 wire \w[10][23] ;
 wire \w[10][24] ;
 wire \w[10][25] ;
 wire \w[10][26] ;
 wire \w[10][27] ;
 wire \w[10][28] ;
 wire \w[10][29] ;
 wire \w[10][2] ;
 wire \w[10][30] ;
 wire \w[10][31] ;
 wire \w[10][3] ;
 wire \w[10][4] ;
 wire \w[10][5] ;
 wire \w[10][6] ;
 wire \w[10][7] ;
 wire \w[10][8] ;
 wire \w[10][9] ;
 wire \w[11][0] ;
 wire \w[11][10] ;
 wire \w[11][11] ;
 wire \w[11][12] ;
 wire \w[11][13] ;
 wire \w[11][14] ;
 wire \w[11][15] ;
 wire \w[11][16] ;
 wire \w[11][17] ;
 wire \w[11][18] ;
 wire \w[11][19] ;
 wire \w[11][1] ;
 wire \w[11][20] ;
 wire \w[11][21] ;
 wire \w[11][22] ;
 wire \w[11][23] ;
 wire \w[11][24] ;
 wire \w[11][25] ;
 wire \w[11][26] ;
 wire \w[11][27] ;
 wire \w[11][28] ;
 wire \w[11][29] ;
 wire \w[11][2] ;
 wire \w[11][30] ;
 wire \w[11][31] ;
 wire \w[11][3] ;
 wire \w[11][4] ;
 wire \w[11][5] ;
 wire \w[11][6] ;
 wire \w[11][7] ;
 wire \w[11][8] ;
 wire \w[11][9] ;
 wire \w[12][0] ;
 wire \w[12][10] ;
 wire \w[12][11] ;
 wire \w[12][12] ;
 wire \w[12][13] ;
 wire \w[12][14] ;
 wire \w[12][15] ;
 wire \w[12][16] ;
 wire \w[12][17] ;
 wire \w[12][18] ;
 wire \w[12][19] ;
 wire \w[12][1] ;
 wire \w[12][20] ;
 wire \w[12][21] ;
 wire \w[12][22] ;
 wire \w[12][23] ;
 wire \w[12][24] ;
 wire \w[12][25] ;
 wire \w[12][26] ;
 wire \w[12][27] ;
 wire \w[12][28] ;
 wire \w[12][29] ;
 wire \w[12][2] ;
 wire \w[12][30] ;
 wire \w[12][31] ;
 wire \w[12][3] ;
 wire \w[12][4] ;
 wire \w[12][5] ;
 wire \w[12][6] ;
 wire \w[12][7] ;
 wire \w[12][8] ;
 wire \w[12][9] ;
 wire \w[13][0] ;
 wire \w[13][10] ;
 wire \w[13][11] ;
 wire \w[13][12] ;
 wire \w[13][13] ;
 wire \w[13][14] ;
 wire \w[13][15] ;
 wire \w[13][16] ;
 wire \w[13][17] ;
 wire \w[13][18] ;
 wire \w[13][19] ;
 wire \w[13][1] ;
 wire \w[13][20] ;
 wire \w[13][21] ;
 wire \w[13][22] ;
 wire \w[13][23] ;
 wire \w[13][24] ;
 wire \w[13][25] ;
 wire \w[13][26] ;
 wire \w[13][27] ;
 wire \w[13][28] ;
 wire \w[13][29] ;
 wire \w[13][2] ;
 wire \w[13][30] ;
 wire \w[13][31] ;
 wire \w[13][3] ;
 wire \w[13][4] ;
 wire \w[13][5] ;
 wire \w[13][6] ;
 wire \w[13][7] ;
 wire \w[13][8] ;
 wire \w[13][9] ;
 wire \w[14][0] ;
 wire \w[14][10] ;
 wire \w[14][11] ;
 wire \w[14][12] ;
 wire \w[14][13] ;
 wire \w[14][14] ;
 wire \w[14][15] ;
 wire \w[14][16] ;
 wire \w[14][17] ;
 wire \w[14][18] ;
 wire \w[14][19] ;
 wire \w[14][1] ;
 wire \w[14][20] ;
 wire \w[14][21] ;
 wire \w[14][22] ;
 wire \w[14][23] ;
 wire \w[14][24] ;
 wire \w[14][25] ;
 wire \w[14][26] ;
 wire \w[14][27] ;
 wire \w[14][28] ;
 wire \w[14][29] ;
 wire \w[14][2] ;
 wire \w[14][30] ;
 wire \w[14][31] ;
 wire \w[14][3] ;
 wire \w[14][4] ;
 wire \w[14][5] ;
 wire \w[14][6] ;
 wire \w[14][7] ;
 wire \w[14][8] ;
 wire \w[14][9] ;
 wire \w[15][0] ;
 wire \w[15][10] ;
 wire \w[15][11] ;
 wire \w[15][12] ;
 wire \w[15][13] ;
 wire \w[15][14] ;
 wire \w[15][15] ;
 wire \w[15][16] ;
 wire \w[15][17] ;
 wire \w[15][18] ;
 wire \w[15][19] ;
 wire \w[15][1] ;
 wire \w[15][20] ;
 wire \w[15][21] ;
 wire \w[15][22] ;
 wire \w[15][23] ;
 wire \w[15][24] ;
 wire \w[15][25] ;
 wire \w[15][26] ;
 wire \w[15][27] ;
 wire \w[15][28] ;
 wire \w[15][29] ;
 wire \w[15][2] ;
 wire \w[15][30] ;
 wire \w[15][31] ;
 wire \w[15][3] ;
 wire \w[15][4] ;
 wire \w[15][5] ;
 wire \w[15][6] ;
 wire \w[15][7] ;
 wire \w[15][8] ;
 wire \w[15][9] ;
 wire \w[16][0] ;
 wire \w[16][10] ;
 wire \w[16][11] ;
 wire \w[16][12] ;
 wire \w[16][13] ;
 wire \w[16][14] ;
 wire \w[16][15] ;
 wire \w[16][16] ;
 wire \w[16][17] ;
 wire \w[16][18] ;
 wire \w[16][19] ;
 wire \w[16][1] ;
 wire \w[16][20] ;
 wire \w[16][21] ;
 wire \w[16][22] ;
 wire \w[16][23] ;
 wire \w[16][24] ;
 wire \w[16][25] ;
 wire \w[16][26] ;
 wire \w[16][27] ;
 wire \w[16][28] ;
 wire \w[16][29] ;
 wire \w[16][2] ;
 wire \w[16][30] ;
 wire \w[16][31] ;
 wire \w[16][3] ;
 wire \w[16][4] ;
 wire \w[16][5] ;
 wire \w[16][6] ;
 wire \w[16][7] ;
 wire \w[16][8] ;
 wire \w[16][9] ;
 wire \w[17][0] ;
 wire \w[17][10] ;
 wire \w[17][11] ;
 wire \w[17][12] ;
 wire \w[17][13] ;
 wire \w[17][14] ;
 wire \w[17][15] ;
 wire \w[17][16] ;
 wire \w[17][17] ;
 wire \w[17][18] ;
 wire \w[17][19] ;
 wire \w[17][1] ;
 wire \w[17][20] ;
 wire \w[17][21] ;
 wire \w[17][22] ;
 wire \w[17][23] ;
 wire \w[17][24] ;
 wire \w[17][25] ;
 wire \w[17][26] ;
 wire \w[17][27] ;
 wire \w[17][28] ;
 wire \w[17][29] ;
 wire \w[17][2] ;
 wire \w[17][30] ;
 wire \w[17][31] ;
 wire \w[17][3] ;
 wire \w[17][4] ;
 wire \w[17][5] ;
 wire \w[17][6] ;
 wire \w[17][7] ;
 wire \w[17][8] ;
 wire \w[17][9] ;
 wire \w[18][0] ;
 wire \w[18][10] ;
 wire \w[18][11] ;
 wire \w[18][12] ;
 wire \w[18][13] ;
 wire \w[18][14] ;
 wire \w[18][15] ;
 wire \w[18][16] ;
 wire \w[18][17] ;
 wire \w[18][18] ;
 wire \w[18][19] ;
 wire \w[18][1] ;
 wire \w[18][20] ;
 wire \w[18][21] ;
 wire \w[18][22] ;
 wire \w[18][23] ;
 wire \w[18][24] ;
 wire \w[18][25] ;
 wire \w[18][26] ;
 wire \w[18][27] ;
 wire \w[18][28] ;
 wire \w[18][29] ;
 wire \w[18][2] ;
 wire \w[18][30] ;
 wire \w[18][31] ;
 wire \w[18][3] ;
 wire \w[18][4] ;
 wire \w[18][5] ;
 wire \w[18][6] ;
 wire \w[18][7] ;
 wire \w[18][8] ;
 wire \w[18][9] ;
 wire \w[19][0] ;
 wire \w[19][10] ;
 wire \w[19][11] ;
 wire \w[19][12] ;
 wire \w[19][13] ;
 wire \w[19][14] ;
 wire \w[19][15] ;
 wire \w[19][16] ;
 wire \w[19][17] ;
 wire \w[19][18] ;
 wire \w[19][19] ;
 wire \w[19][1] ;
 wire \w[19][20] ;
 wire \w[19][21] ;
 wire \w[19][22] ;
 wire \w[19][23] ;
 wire \w[19][24] ;
 wire \w[19][25] ;
 wire \w[19][26] ;
 wire \w[19][27] ;
 wire \w[19][28] ;
 wire \w[19][29] ;
 wire \w[19][2] ;
 wire \w[19][30] ;
 wire \w[19][31] ;
 wire \w[19][3] ;
 wire \w[19][4] ;
 wire \w[19][5] ;
 wire \w[19][6] ;
 wire \w[19][7] ;
 wire \w[19][8] ;
 wire \w[19][9] ;
 wire \w[1][0] ;
 wire \w[1][10] ;
 wire \w[1][11] ;
 wire \w[1][12] ;
 wire \w[1][13] ;
 wire \w[1][14] ;
 wire \w[1][15] ;
 wire \w[1][16] ;
 wire \w[1][17] ;
 wire \w[1][18] ;
 wire \w[1][19] ;
 wire \w[1][1] ;
 wire \w[1][20] ;
 wire \w[1][21] ;
 wire \w[1][22] ;
 wire \w[1][23] ;
 wire \w[1][24] ;
 wire \w[1][25] ;
 wire \w[1][26] ;
 wire \w[1][27] ;
 wire \w[1][28] ;
 wire \w[1][29] ;
 wire \w[1][2] ;
 wire \w[1][30] ;
 wire \w[1][31] ;
 wire \w[1][3] ;
 wire \w[1][4] ;
 wire \w[1][5] ;
 wire \w[1][6] ;
 wire \w[1][7] ;
 wire \w[1][8] ;
 wire \w[1][9] ;
 wire \w[20][0] ;
 wire \w[20][10] ;
 wire \w[20][11] ;
 wire \w[20][12] ;
 wire \w[20][13] ;
 wire \w[20][14] ;
 wire \w[20][15] ;
 wire \w[20][16] ;
 wire \w[20][17] ;
 wire \w[20][18] ;
 wire \w[20][19] ;
 wire \w[20][1] ;
 wire \w[20][20] ;
 wire \w[20][21] ;
 wire \w[20][22] ;
 wire \w[20][23] ;
 wire \w[20][24] ;
 wire \w[20][25] ;
 wire \w[20][26] ;
 wire \w[20][27] ;
 wire \w[20][28] ;
 wire \w[20][29] ;
 wire \w[20][2] ;
 wire \w[20][30] ;
 wire \w[20][31] ;
 wire \w[20][3] ;
 wire \w[20][4] ;
 wire \w[20][5] ;
 wire \w[20][6] ;
 wire \w[20][7] ;
 wire \w[20][8] ;
 wire \w[20][9] ;
 wire \w[21][0] ;
 wire \w[21][10] ;
 wire \w[21][11] ;
 wire \w[21][12] ;
 wire \w[21][13] ;
 wire \w[21][14] ;
 wire \w[21][15] ;
 wire \w[21][16] ;
 wire \w[21][17] ;
 wire \w[21][18] ;
 wire \w[21][19] ;
 wire \w[21][1] ;
 wire \w[21][20] ;
 wire \w[21][21] ;
 wire \w[21][22] ;
 wire \w[21][23] ;
 wire \w[21][24] ;
 wire \w[21][25] ;
 wire \w[21][26] ;
 wire \w[21][27] ;
 wire \w[21][28] ;
 wire \w[21][29] ;
 wire \w[21][2] ;
 wire \w[21][30] ;
 wire \w[21][31] ;
 wire \w[21][3] ;
 wire \w[21][4] ;
 wire \w[21][5] ;
 wire \w[21][6] ;
 wire \w[21][7] ;
 wire \w[21][8] ;
 wire \w[21][9] ;
 wire \w[22][0] ;
 wire \w[22][10] ;
 wire \w[22][11] ;
 wire \w[22][12] ;
 wire \w[22][13] ;
 wire \w[22][14] ;
 wire \w[22][15] ;
 wire \w[22][16] ;
 wire \w[22][17] ;
 wire \w[22][18] ;
 wire \w[22][19] ;
 wire \w[22][1] ;
 wire \w[22][20] ;
 wire \w[22][21] ;
 wire \w[22][22] ;
 wire \w[22][23] ;
 wire \w[22][24] ;
 wire \w[22][25] ;
 wire \w[22][26] ;
 wire \w[22][27] ;
 wire \w[22][28] ;
 wire \w[22][29] ;
 wire \w[22][2] ;
 wire \w[22][30] ;
 wire \w[22][31] ;
 wire \w[22][3] ;
 wire \w[22][4] ;
 wire \w[22][5] ;
 wire \w[22][6] ;
 wire \w[22][7] ;
 wire \w[22][8] ;
 wire \w[22][9] ;
 wire \w[23][0] ;
 wire \w[23][10] ;
 wire \w[23][11] ;
 wire \w[23][12] ;
 wire \w[23][13] ;
 wire \w[23][14] ;
 wire \w[23][15] ;
 wire \w[23][16] ;
 wire \w[23][17] ;
 wire \w[23][18] ;
 wire \w[23][19] ;
 wire \w[23][1] ;
 wire \w[23][20] ;
 wire \w[23][21] ;
 wire \w[23][22] ;
 wire \w[23][23] ;
 wire \w[23][24] ;
 wire \w[23][25] ;
 wire \w[23][26] ;
 wire \w[23][27] ;
 wire \w[23][28] ;
 wire \w[23][29] ;
 wire \w[23][2] ;
 wire \w[23][30] ;
 wire \w[23][31] ;
 wire \w[23][3] ;
 wire \w[23][4] ;
 wire \w[23][5] ;
 wire \w[23][6] ;
 wire \w[23][7] ;
 wire \w[23][8] ;
 wire \w[23][9] ;
 wire \w[24][0] ;
 wire \w[24][10] ;
 wire \w[24][11] ;
 wire \w[24][12] ;
 wire \w[24][13] ;
 wire \w[24][14] ;
 wire \w[24][15] ;
 wire \w[24][16] ;
 wire \w[24][17] ;
 wire \w[24][18] ;
 wire \w[24][19] ;
 wire \w[24][1] ;
 wire \w[24][20] ;
 wire \w[24][21] ;
 wire \w[24][22] ;
 wire \w[24][23] ;
 wire \w[24][24] ;
 wire \w[24][25] ;
 wire \w[24][26] ;
 wire \w[24][27] ;
 wire \w[24][28] ;
 wire \w[24][29] ;
 wire \w[24][2] ;
 wire \w[24][30] ;
 wire \w[24][31] ;
 wire \w[24][3] ;
 wire \w[24][4] ;
 wire \w[24][5] ;
 wire \w[24][6] ;
 wire \w[24][7] ;
 wire \w[24][8] ;
 wire \w[24][9] ;
 wire \w[25][0] ;
 wire \w[25][10] ;
 wire \w[25][11] ;
 wire \w[25][12] ;
 wire \w[25][13] ;
 wire \w[25][14] ;
 wire \w[25][15] ;
 wire \w[25][16] ;
 wire \w[25][17] ;
 wire \w[25][18] ;
 wire \w[25][19] ;
 wire \w[25][1] ;
 wire \w[25][20] ;
 wire \w[25][21] ;
 wire \w[25][22] ;
 wire \w[25][23] ;
 wire \w[25][24] ;
 wire \w[25][25] ;
 wire \w[25][26] ;
 wire \w[25][27] ;
 wire \w[25][28] ;
 wire \w[25][29] ;
 wire \w[25][2] ;
 wire \w[25][30] ;
 wire \w[25][31] ;
 wire \w[25][3] ;
 wire \w[25][4] ;
 wire \w[25][5] ;
 wire \w[25][6] ;
 wire \w[25][7] ;
 wire \w[25][8] ;
 wire \w[25][9] ;
 wire \w[26][0] ;
 wire \w[26][10] ;
 wire \w[26][11] ;
 wire \w[26][12] ;
 wire \w[26][13] ;
 wire \w[26][14] ;
 wire \w[26][15] ;
 wire \w[26][16] ;
 wire \w[26][17] ;
 wire \w[26][18] ;
 wire \w[26][19] ;
 wire \w[26][1] ;
 wire \w[26][20] ;
 wire \w[26][21] ;
 wire \w[26][22] ;
 wire \w[26][23] ;
 wire \w[26][24] ;
 wire \w[26][25] ;
 wire \w[26][26] ;
 wire \w[26][27] ;
 wire \w[26][28] ;
 wire \w[26][29] ;
 wire \w[26][2] ;
 wire \w[26][30] ;
 wire \w[26][31] ;
 wire \w[26][3] ;
 wire \w[26][4] ;
 wire \w[26][5] ;
 wire \w[26][6] ;
 wire \w[26][7] ;
 wire \w[26][8] ;
 wire \w[26][9] ;
 wire \w[27][0] ;
 wire \w[27][10] ;
 wire \w[27][11] ;
 wire \w[27][12] ;
 wire \w[27][13] ;
 wire \w[27][14] ;
 wire \w[27][15] ;
 wire \w[27][16] ;
 wire \w[27][17] ;
 wire \w[27][18] ;
 wire \w[27][19] ;
 wire \w[27][1] ;
 wire \w[27][20] ;
 wire \w[27][21] ;
 wire \w[27][22] ;
 wire \w[27][23] ;
 wire \w[27][24] ;
 wire \w[27][25] ;
 wire \w[27][26] ;
 wire \w[27][27] ;
 wire \w[27][28] ;
 wire \w[27][29] ;
 wire \w[27][2] ;
 wire \w[27][30] ;
 wire \w[27][31] ;
 wire \w[27][3] ;
 wire \w[27][4] ;
 wire \w[27][5] ;
 wire \w[27][6] ;
 wire \w[27][7] ;
 wire \w[27][8] ;
 wire \w[27][9] ;
 wire \w[28][0] ;
 wire \w[28][10] ;
 wire \w[28][11] ;
 wire \w[28][12] ;
 wire \w[28][13] ;
 wire \w[28][14] ;
 wire \w[28][15] ;
 wire \w[28][16] ;
 wire \w[28][17] ;
 wire \w[28][18] ;
 wire \w[28][19] ;
 wire \w[28][1] ;
 wire \w[28][20] ;
 wire \w[28][21] ;
 wire \w[28][22] ;
 wire \w[28][23] ;
 wire \w[28][24] ;
 wire \w[28][25] ;
 wire \w[28][26] ;
 wire \w[28][27] ;
 wire \w[28][28] ;
 wire \w[28][29] ;
 wire \w[28][2] ;
 wire \w[28][30] ;
 wire \w[28][31] ;
 wire \w[28][3] ;
 wire \w[28][4] ;
 wire \w[28][5] ;
 wire \w[28][6] ;
 wire \w[28][7] ;
 wire \w[28][8] ;
 wire \w[28][9] ;
 wire \w[29][0] ;
 wire \w[29][10] ;
 wire \w[29][11] ;
 wire \w[29][12] ;
 wire \w[29][13] ;
 wire \w[29][14] ;
 wire \w[29][15] ;
 wire \w[29][16] ;
 wire \w[29][17] ;
 wire \w[29][18] ;
 wire \w[29][19] ;
 wire \w[29][1] ;
 wire \w[29][20] ;
 wire \w[29][21] ;
 wire \w[29][22] ;
 wire \w[29][23] ;
 wire \w[29][24] ;
 wire \w[29][25] ;
 wire \w[29][26] ;
 wire \w[29][27] ;
 wire \w[29][28] ;
 wire \w[29][29] ;
 wire \w[29][2] ;
 wire \w[29][30] ;
 wire \w[29][31] ;
 wire \w[29][3] ;
 wire \w[29][4] ;
 wire \w[29][5] ;
 wire \w[29][6] ;
 wire \w[29][7] ;
 wire \w[29][8] ;
 wire \w[29][9] ;
 wire \w[2][0] ;
 wire \w[2][10] ;
 wire \w[2][11] ;
 wire \w[2][12] ;
 wire \w[2][13] ;
 wire \w[2][14] ;
 wire \w[2][15] ;
 wire \w[2][16] ;
 wire \w[2][17] ;
 wire \w[2][18] ;
 wire \w[2][19] ;
 wire \w[2][1] ;
 wire \w[2][20] ;
 wire \w[2][21] ;
 wire \w[2][22] ;
 wire \w[2][23] ;
 wire \w[2][24] ;
 wire \w[2][25] ;
 wire \w[2][26] ;
 wire \w[2][27] ;
 wire \w[2][28] ;
 wire \w[2][29] ;
 wire \w[2][2] ;
 wire \w[2][30] ;
 wire \w[2][31] ;
 wire \w[2][3] ;
 wire \w[2][4] ;
 wire \w[2][5] ;
 wire \w[2][6] ;
 wire \w[2][7] ;
 wire \w[2][8] ;
 wire \w[2][9] ;
 wire \w[30][0] ;
 wire \w[30][10] ;
 wire \w[30][11] ;
 wire \w[30][12] ;
 wire \w[30][13] ;
 wire \w[30][14] ;
 wire \w[30][15] ;
 wire \w[30][16] ;
 wire \w[30][17] ;
 wire \w[30][18] ;
 wire \w[30][19] ;
 wire \w[30][1] ;
 wire \w[30][20] ;
 wire \w[30][21] ;
 wire \w[30][22] ;
 wire \w[30][23] ;
 wire \w[30][24] ;
 wire \w[30][25] ;
 wire \w[30][26] ;
 wire \w[30][27] ;
 wire \w[30][28] ;
 wire \w[30][29] ;
 wire \w[30][2] ;
 wire \w[30][30] ;
 wire \w[30][31] ;
 wire \w[30][3] ;
 wire \w[30][4] ;
 wire \w[30][5] ;
 wire \w[30][6] ;
 wire \w[30][7] ;
 wire \w[30][8] ;
 wire \w[30][9] ;
 wire \w[31][0] ;
 wire \w[31][10] ;
 wire \w[31][11] ;
 wire \w[31][12] ;
 wire \w[31][13] ;
 wire \w[31][14] ;
 wire \w[31][15] ;
 wire \w[31][16] ;
 wire \w[31][17] ;
 wire \w[31][18] ;
 wire \w[31][19] ;
 wire \w[31][1] ;
 wire \w[31][20] ;
 wire \w[31][21] ;
 wire \w[31][22] ;
 wire \w[31][23] ;
 wire \w[31][24] ;
 wire \w[31][25] ;
 wire \w[31][26] ;
 wire \w[31][27] ;
 wire \w[31][28] ;
 wire \w[31][29] ;
 wire \w[31][2] ;
 wire \w[31][30] ;
 wire \w[31][31] ;
 wire \w[31][3] ;
 wire \w[31][4] ;
 wire \w[31][5] ;
 wire \w[31][6] ;
 wire \w[31][7] ;
 wire \w[31][8] ;
 wire \w[31][9] ;
 wire \w[32][0] ;
 wire \w[32][10] ;
 wire \w[32][11] ;
 wire \w[32][12] ;
 wire \w[32][13] ;
 wire \w[32][14] ;
 wire \w[32][15] ;
 wire \w[32][16] ;
 wire \w[32][17] ;
 wire \w[32][18] ;
 wire \w[32][19] ;
 wire \w[32][1] ;
 wire \w[32][20] ;
 wire \w[32][21] ;
 wire \w[32][22] ;
 wire \w[32][23] ;
 wire \w[32][24] ;
 wire \w[32][25] ;
 wire \w[32][26] ;
 wire \w[32][27] ;
 wire \w[32][28] ;
 wire \w[32][29] ;
 wire \w[32][2] ;
 wire \w[32][30] ;
 wire \w[32][31] ;
 wire \w[32][3] ;
 wire \w[32][4] ;
 wire \w[32][5] ;
 wire \w[32][6] ;
 wire \w[32][7] ;
 wire \w[32][8] ;
 wire \w[32][9] ;
 wire \w[33][0] ;
 wire \w[33][10] ;
 wire \w[33][11] ;
 wire \w[33][12] ;
 wire \w[33][13] ;
 wire \w[33][14] ;
 wire \w[33][15] ;
 wire \w[33][16] ;
 wire \w[33][17] ;
 wire \w[33][18] ;
 wire \w[33][19] ;
 wire \w[33][1] ;
 wire \w[33][20] ;
 wire \w[33][21] ;
 wire \w[33][22] ;
 wire \w[33][23] ;
 wire \w[33][24] ;
 wire \w[33][25] ;
 wire \w[33][26] ;
 wire \w[33][27] ;
 wire \w[33][28] ;
 wire \w[33][29] ;
 wire \w[33][2] ;
 wire \w[33][30] ;
 wire \w[33][31] ;
 wire \w[33][3] ;
 wire \w[33][4] ;
 wire \w[33][5] ;
 wire \w[33][6] ;
 wire \w[33][7] ;
 wire \w[33][8] ;
 wire \w[33][9] ;
 wire \w[34][0] ;
 wire \w[34][10] ;
 wire \w[34][11] ;
 wire \w[34][12] ;
 wire \w[34][13] ;
 wire \w[34][14] ;
 wire \w[34][15] ;
 wire \w[34][16] ;
 wire \w[34][17] ;
 wire \w[34][18] ;
 wire \w[34][19] ;
 wire \w[34][1] ;
 wire \w[34][20] ;
 wire \w[34][21] ;
 wire \w[34][22] ;
 wire \w[34][23] ;
 wire \w[34][24] ;
 wire \w[34][25] ;
 wire \w[34][26] ;
 wire \w[34][27] ;
 wire \w[34][28] ;
 wire \w[34][29] ;
 wire \w[34][2] ;
 wire \w[34][30] ;
 wire \w[34][31] ;
 wire \w[34][3] ;
 wire \w[34][4] ;
 wire \w[34][5] ;
 wire \w[34][6] ;
 wire \w[34][7] ;
 wire \w[34][8] ;
 wire \w[34][9] ;
 wire \w[35][0] ;
 wire \w[35][10] ;
 wire \w[35][11] ;
 wire \w[35][12] ;
 wire \w[35][13] ;
 wire \w[35][14] ;
 wire \w[35][15] ;
 wire \w[35][16] ;
 wire \w[35][17] ;
 wire \w[35][18] ;
 wire \w[35][19] ;
 wire \w[35][1] ;
 wire \w[35][20] ;
 wire \w[35][21] ;
 wire \w[35][22] ;
 wire \w[35][23] ;
 wire \w[35][24] ;
 wire \w[35][25] ;
 wire \w[35][26] ;
 wire \w[35][27] ;
 wire \w[35][28] ;
 wire \w[35][29] ;
 wire \w[35][2] ;
 wire \w[35][30] ;
 wire \w[35][31] ;
 wire \w[35][3] ;
 wire \w[35][4] ;
 wire \w[35][5] ;
 wire \w[35][6] ;
 wire \w[35][7] ;
 wire \w[35][8] ;
 wire \w[35][9] ;
 wire \w[36][0] ;
 wire \w[36][10] ;
 wire \w[36][11] ;
 wire \w[36][12] ;
 wire \w[36][13] ;
 wire \w[36][14] ;
 wire \w[36][15] ;
 wire \w[36][16] ;
 wire \w[36][17] ;
 wire \w[36][18] ;
 wire \w[36][19] ;
 wire \w[36][1] ;
 wire \w[36][20] ;
 wire \w[36][21] ;
 wire \w[36][22] ;
 wire \w[36][23] ;
 wire \w[36][24] ;
 wire \w[36][25] ;
 wire \w[36][26] ;
 wire \w[36][27] ;
 wire \w[36][28] ;
 wire \w[36][29] ;
 wire \w[36][2] ;
 wire \w[36][30] ;
 wire \w[36][31] ;
 wire \w[36][3] ;
 wire \w[36][4] ;
 wire \w[36][5] ;
 wire \w[36][6] ;
 wire \w[36][7] ;
 wire \w[36][8] ;
 wire \w[36][9] ;
 wire \w[37][0] ;
 wire \w[37][10] ;
 wire \w[37][11] ;
 wire \w[37][12] ;
 wire \w[37][13] ;
 wire \w[37][14] ;
 wire \w[37][15] ;
 wire \w[37][16] ;
 wire \w[37][17] ;
 wire \w[37][18] ;
 wire \w[37][19] ;
 wire \w[37][1] ;
 wire \w[37][20] ;
 wire \w[37][21] ;
 wire \w[37][22] ;
 wire \w[37][23] ;
 wire \w[37][24] ;
 wire \w[37][25] ;
 wire \w[37][26] ;
 wire \w[37][27] ;
 wire \w[37][28] ;
 wire \w[37][29] ;
 wire \w[37][2] ;
 wire \w[37][30] ;
 wire \w[37][31] ;
 wire \w[37][3] ;
 wire \w[37][4] ;
 wire \w[37][5] ;
 wire \w[37][6] ;
 wire \w[37][7] ;
 wire \w[37][8] ;
 wire \w[37][9] ;
 wire \w[38][0] ;
 wire \w[38][10] ;
 wire \w[38][11] ;
 wire \w[38][12] ;
 wire \w[38][13] ;
 wire \w[38][14] ;
 wire \w[38][15] ;
 wire \w[38][16] ;
 wire \w[38][17] ;
 wire \w[38][18] ;
 wire \w[38][19] ;
 wire \w[38][1] ;
 wire \w[38][20] ;
 wire \w[38][21] ;
 wire \w[38][22] ;
 wire \w[38][23] ;
 wire \w[38][24] ;
 wire \w[38][25] ;
 wire \w[38][26] ;
 wire \w[38][27] ;
 wire \w[38][28] ;
 wire \w[38][29] ;
 wire \w[38][2] ;
 wire \w[38][30] ;
 wire \w[38][31] ;
 wire \w[38][3] ;
 wire \w[38][4] ;
 wire \w[38][5] ;
 wire \w[38][6] ;
 wire \w[38][7] ;
 wire \w[38][8] ;
 wire \w[38][9] ;
 wire \w[39][0] ;
 wire \w[39][10] ;
 wire \w[39][11] ;
 wire \w[39][12] ;
 wire \w[39][13] ;
 wire \w[39][14] ;
 wire \w[39][15] ;
 wire \w[39][16] ;
 wire \w[39][17] ;
 wire \w[39][18] ;
 wire \w[39][19] ;
 wire \w[39][1] ;
 wire \w[39][20] ;
 wire \w[39][21] ;
 wire \w[39][22] ;
 wire \w[39][23] ;
 wire \w[39][24] ;
 wire \w[39][25] ;
 wire \w[39][26] ;
 wire \w[39][27] ;
 wire \w[39][28] ;
 wire \w[39][29] ;
 wire \w[39][2] ;
 wire \w[39][30] ;
 wire \w[39][31] ;
 wire \w[39][3] ;
 wire \w[39][4] ;
 wire \w[39][5] ;
 wire \w[39][6] ;
 wire \w[39][7] ;
 wire \w[39][8] ;
 wire \w[39][9] ;
 wire \w[3][0] ;
 wire \w[3][10] ;
 wire \w[3][11] ;
 wire \w[3][12] ;
 wire \w[3][13] ;
 wire \w[3][14] ;
 wire \w[3][15] ;
 wire \w[3][16] ;
 wire \w[3][17] ;
 wire \w[3][18] ;
 wire \w[3][19] ;
 wire \w[3][1] ;
 wire \w[3][20] ;
 wire \w[3][21] ;
 wire \w[3][22] ;
 wire \w[3][23] ;
 wire \w[3][24] ;
 wire \w[3][25] ;
 wire \w[3][26] ;
 wire \w[3][27] ;
 wire \w[3][28] ;
 wire \w[3][29] ;
 wire \w[3][2] ;
 wire \w[3][30] ;
 wire \w[3][31] ;
 wire \w[3][3] ;
 wire \w[3][4] ;
 wire \w[3][5] ;
 wire \w[3][6] ;
 wire \w[3][7] ;
 wire \w[3][8] ;
 wire \w[3][9] ;
 wire \w[40][0] ;
 wire \w[40][10] ;
 wire \w[40][11] ;
 wire \w[40][12] ;
 wire \w[40][13] ;
 wire \w[40][14] ;
 wire \w[40][15] ;
 wire \w[40][16] ;
 wire \w[40][17] ;
 wire \w[40][18] ;
 wire \w[40][19] ;
 wire \w[40][1] ;
 wire \w[40][20] ;
 wire \w[40][21] ;
 wire \w[40][22] ;
 wire \w[40][23] ;
 wire \w[40][24] ;
 wire \w[40][25] ;
 wire \w[40][26] ;
 wire \w[40][27] ;
 wire \w[40][28] ;
 wire \w[40][29] ;
 wire \w[40][2] ;
 wire \w[40][30] ;
 wire \w[40][31] ;
 wire \w[40][3] ;
 wire \w[40][4] ;
 wire \w[40][5] ;
 wire \w[40][6] ;
 wire \w[40][7] ;
 wire \w[40][8] ;
 wire \w[40][9] ;
 wire \w[41][0] ;
 wire \w[41][10] ;
 wire \w[41][11] ;
 wire \w[41][12] ;
 wire \w[41][13] ;
 wire \w[41][14] ;
 wire \w[41][15] ;
 wire \w[41][16] ;
 wire \w[41][17] ;
 wire \w[41][18] ;
 wire \w[41][19] ;
 wire \w[41][1] ;
 wire \w[41][20] ;
 wire \w[41][21] ;
 wire \w[41][22] ;
 wire \w[41][23] ;
 wire \w[41][24] ;
 wire \w[41][25] ;
 wire \w[41][26] ;
 wire \w[41][27] ;
 wire \w[41][28] ;
 wire \w[41][29] ;
 wire \w[41][2] ;
 wire \w[41][30] ;
 wire \w[41][31] ;
 wire \w[41][3] ;
 wire \w[41][4] ;
 wire \w[41][5] ;
 wire \w[41][6] ;
 wire \w[41][7] ;
 wire \w[41][8] ;
 wire \w[41][9] ;
 wire \w[42][0] ;
 wire \w[42][10] ;
 wire \w[42][11] ;
 wire \w[42][12] ;
 wire \w[42][13] ;
 wire \w[42][14] ;
 wire \w[42][15] ;
 wire \w[42][16] ;
 wire \w[42][17] ;
 wire \w[42][18] ;
 wire \w[42][19] ;
 wire \w[42][1] ;
 wire \w[42][20] ;
 wire \w[42][21] ;
 wire \w[42][22] ;
 wire \w[42][23] ;
 wire \w[42][24] ;
 wire \w[42][25] ;
 wire \w[42][26] ;
 wire \w[42][27] ;
 wire \w[42][28] ;
 wire \w[42][29] ;
 wire \w[42][2] ;
 wire \w[42][30] ;
 wire \w[42][31] ;
 wire \w[42][3] ;
 wire \w[42][4] ;
 wire \w[42][5] ;
 wire \w[42][6] ;
 wire \w[42][7] ;
 wire \w[42][8] ;
 wire \w[42][9] ;
 wire \w[43][0] ;
 wire \w[43][10] ;
 wire \w[43][11] ;
 wire \w[43][12] ;
 wire \w[43][13] ;
 wire \w[43][14] ;
 wire \w[43][15] ;
 wire \w[43][16] ;
 wire \w[43][17] ;
 wire \w[43][18] ;
 wire \w[43][19] ;
 wire \w[43][1] ;
 wire \w[43][20] ;
 wire \w[43][21] ;
 wire \w[43][22] ;
 wire \w[43][23] ;
 wire \w[43][24] ;
 wire \w[43][25] ;
 wire \w[43][26] ;
 wire \w[43][27] ;
 wire \w[43][28] ;
 wire \w[43][29] ;
 wire \w[43][2] ;
 wire \w[43][30] ;
 wire \w[43][31] ;
 wire \w[43][3] ;
 wire \w[43][4] ;
 wire \w[43][5] ;
 wire \w[43][6] ;
 wire \w[43][7] ;
 wire \w[43][8] ;
 wire \w[43][9] ;
 wire \w[44][0] ;
 wire \w[44][10] ;
 wire \w[44][11] ;
 wire \w[44][12] ;
 wire \w[44][13] ;
 wire \w[44][14] ;
 wire \w[44][15] ;
 wire \w[44][16] ;
 wire \w[44][17] ;
 wire \w[44][18] ;
 wire \w[44][19] ;
 wire \w[44][1] ;
 wire \w[44][20] ;
 wire \w[44][21] ;
 wire \w[44][22] ;
 wire \w[44][23] ;
 wire \w[44][24] ;
 wire \w[44][25] ;
 wire \w[44][26] ;
 wire \w[44][27] ;
 wire \w[44][28] ;
 wire \w[44][29] ;
 wire \w[44][2] ;
 wire \w[44][30] ;
 wire \w[44][31] ;
 wire \w[44][3] ;
 wire \w[44][4] ;
 wire \w[44][5] ;
 wire \w[44][6] ;
 wire \w[44][7] ;
 wire \w[44][8] ;
 wire \w[44][9] ;
 wire \w[45][0] ;
 wire \w[45][10] ;
 wire \w[45][11] ;
 wire \w[45][12] ;
 wire \w[45][13] ;
 wire \w[45][14] ;
 wire \w[45][15] ;
 wire \w[45][16] ;
 wire \w[45][17] ;
 wire \w[45][18] ;
 wire \w[45][19] ;
 wire \w[45][1] ;
 wire \w[45][20] ;
 wire \w[45][21] ;
 wire \w[45][22] ;
 wire \w[45][23] ;
 wire \w[45][24] ;
 wire \w[45][25] ;
 wire \w[45][26] ;
 wire \w[45][27] ;
 wire \w[45][28] ;
 wire \w[45][29] ;
 wire \w[45][2] ;
 wire \w[45][30] ;
 wire \w[45][31] ;
 wire \w[45][3] ;
 wire \w[45][4] ;
 wire \w[45][5] ;
 wire \w[45][6] ;
 wire \w[45][7] ;
 wire \w[45][8] ;
 wire \w[45][9] ;
 wire \w[46][0] ;
 wire \w[46][10] ;
 wire \w[46][11] ;
 wire \w[46][12] ;
 wire \w[46][13] ;
 wire \w[46][14] ;
 wire \w[46][15] ;
 wire \w[46][16] ;
 wire \w[46][17] ;
 wire \w[46][18] ;
 wire \w[46][19] ;
 wire \w[46][1] ;
 wire \w[46][20] ;
 wire \w[46][21] ;
 wire \w[46][22] ;
 wire \w[46][23] ;
 wire \w[46][24] ;
 wire \w[46][25] ;
 wire \w[46][26] ;
 wire \w[46][27] ;
 wire \w[46][28] ;
 wire \w[46][29] ;
 wire \w[46][2] ;
 wire \w[46][30] ;
 wire \w[46][31] ;
 wire \w[46][3] ;
 wire \w[46][4] ;
 wire \w[46][5] ;
 wire \w[46][6] ;
 wire \w[46][7] ;
 wire \w[46][8] ;
 wire \w[46][9] ;
 wire \w[47][0] ;
 wire \w[47][10] ;
 wire \w[47][11] ;
 wire \w[47][12] ;
 wire \w[47][13] ;
 wire \w[47][14] ;
 wire \w[47][15] ;
 wire \w[47][16] ;
 wire \w[47][17] ;
 wire \w[47][18] ;
 wire \w[47][19] ;
 wire \w[47][1] ;
 wire \w[47][20] ;
 wire \w[47][21] ;
 wire \w[47][22] ;
 wire \w[47][23] ;
 wire \w[47][24] ;
 wire \w[47][25] ;
 wire \w[47][26] ;
 wire \w[47][27] ;
 wire \w[47][28] ;
 wire \w[47][29] ;
 wire \w[47][2] ;
 wire \w[47][30] ;
 wire \w[47][31] ;
 wire \w[47][3] ;
 wire \w[47][4] ;
 wire \w[47][5] ;
 wire \w[47][6] ;
 wire \w[47][7] ;
 wire \w[47][8] ;
 wire \w[47][9] ;
 wire \w[48][0] ;
 wire \w[48][10] ;
 wire \w[48][11] ;
 wire \w[48][12] ;
 wire \w[48][13] ;
 wire \w[48][14] ;
 wire \w[48][15] ;
 wire \w[48][16] ;
 wire \w[48][17] ;
 wire \w[48][18] ;
 wire \w[48][19] ;
 wire \w[48][1] ;
 wire \w[48][20] ;
 wire \w[48][21] ;
 wire \w[48][22] ;
 wire \w[48][23] ;
 wire \w[48][24] ;
 wire \w[48][25] ;
 wire \w[48][26] ;
 wire \w[48][27] ;
 wire \w[48][28] ;
 wire \w[48][29] ;
 wire \w[48][2] ;
 wire \w[48][30] ;
 wire \w[48][31] ;
 wire \w[48][3] ;
 wire \w[48][4] ;
 wire \w[48][5] ;
 wire \w[48][6] ;
 wire \w[48][7] ;
 wire \w[48][8] ;
 wire \w[48][9] ;
 wire \w[49][0] ;
 wire \w[49][10] ;
 wire \w[49][11] ;
 wire \w[49][12] ;
 wire \w[49][13] ;
 wire \w[49][14] ;
 wire \w[49][15] ;
 wire \w[49][16] ;
 wire \w[49][17] ;
 wire \w[49][18] ;
 wire \w[49][19] ;
 wire \w[49][1] ;
 wire \w[49][20] ;
 wire \w[49][21] ;
 wire \w[49][22] ;
 wire \w[49][23] ;
 wire \w[49][24] ;
 wire \w[49][25] ;
 wire \w[49][26] ;
 wire \w[49][27] ;
 wire \w[49][28] ;
 wire \w[49][29] ;
 wire \w[49][2] ;
 wire \w[49][30] ;
 wire \w[49][31] ;
 wire \w[49][3] ;
 wire \w[49][4] ;
 wire \w[49][5] ;
 wire \w[49][6] ;
 wire \w[49][7] ;
 wire \w[49][8] ;
 wire \w[49][9] ;
 wire \w[4][0] ;
 wire \w[4][10] ;
 wire \w[4][11] ;
 wire \w[4][12] ;
 wire \w[4][13] ;
 wire \w[4][14] ;
 wire \w[4][15] ;
 wire \w[4][16] ;
 wire \w[4][17] ;
 wire \w[4][18] ;
 wire \w[4][19] ;
 wire \w[4][1] ;
 wire \w[4][20] ;
 wire \w[4][21] ;
 wire \w[4][22] ;
 wire \w[4][23] ;
 wire \w[4][24] ;
 wire \w[4][25] ;
 wire \w[4][26] ;
 wire \w[4][27] ;
 wire \w[4][28] ;
 wire \w[4][29] ;
 wire \w[4][2] ;
 wire \w[4][30] ;
 wire \w[4][31] ;
 wire \w[4][3] ;
 wire \w[4][4] ;
 wire \w[4][5] ;
 wire \w[4][6] ;
 wire \w[4][7] ;
 wire \w[4][8] ;
 wire \w[4][9] ;
 wire \w[50][0] ;
 wire \w[50][10] ;
 wire \w[50][11] ;
 wire \w[50][12] ;
 wire \w[50][13] ;
 wire \w[50][14] ;
 wire \w[50][15] ;
 wire \w[50][16] ;
 wire \w[50][17] ;
 wire \w[50][18] ;
 wire \w[50][19] ;
 wire \w[50][1] ;
 wire \w[50][20] ;
 wire \w[50][21] ;
 wire \w[50][22] ;
 wire \w[50][23] ;
 wire \w[50][24] ;
 wire \w[50][25] ;
 wire \w[50][26] ;
 wire \w[50][27] ;
 wire \w[50][28] ;
 wire \w[50][29] ;
 wire \w[50][2] ;
 wire \w[50][30] ;
 wire \w[50][31] ;
 wire \w[50][3] ;
 wire \w[50][4] ;
 wire \w[50][5] ;
 wire \w[50][6] ;
 wire \w[50][7] ;
 wire \w[50][8] ;
 wire \w[50][9] ;
 wire \w[51][0] ;
 wire \w[51][10] ;
 wire \w[51][11] ;
 wire \w[51][12] ;
 wire \w[51][13] ;
 wire \w[51][14] ;
 wire \w[51][15] ;
 wire \w[51][16] ;
 wire \w[51][17] ;
 wire \w[51][18] ;
 wire \w[51][19] ;
 wire \w[51][1] ;
 wire \w[51][20] ;
 wire \w[51][21] ;
 wire \w[51][22] ;
 wire \w[51][23] ;
 wire \w[51][24] ;
 wire \w[51][25] ;
 wire \w[51][26] ;
 wire \w[51][27] ;
 wire \w[51][28] ;
 wire \w[51][29] ;
 wire \w[51][2] ;
 wire \w[51][30] ;
 wire \w[51][31] ;
 wire \w[51][3] ;
 wire \w[51][4] ;
 wire \w[51][5] ;
 wire \w[51][6] ;
 wire \w[51][7] ;
 wire \w[51][8] ;
 wire \w[51][9] ;
 wire \w[52][0] ;
 wire \w[52][10] ;
 wire \w[52][11] ;
 wire \w[52][12] ;
 wire \w[52][13] ;
 wire \w[52][14] ;
 wire \w[52][15] ;
 wire \w[52][16] ;
 wire \w[52][17] ;
 wire \w[52][18] ;
 wire \w[52][19] ;
 wire \w[52][1] ;
 wire \w[52][20] ;
 wire \w[52][21] ;
 wire \w[52][22] ;
 wire \w[52][23] ;
 wire \w[52][24] ;
 wire \w[52][25] ;
 wire \w[52][26] ;
 wire \w[52][27] ;
 wire \w[52][28] ;
 wire \w[52][29] ;
 wire \w[52][2] ;
 wire \w[52][30] ;
 wire \w[52][31] ;
 wire \w[52][3] ;
 wire \w[52][4] ;
 wire \w[52][5] ;
 wire \w[52][6] ;
 wire \w[52][7] ;
 wire \w[52][8] ;
 wire \w[52][9] ;
 wire \w[53][0] ;
 wire \w[53][10] ;
 wire \w[53][11] ;
 wire \w[53][12] ;
 wire \w[53][13] ;
 wire \w[53][14] ;
 wire \w[53][15] ;
 wire \w[53][16] ;
 wire \w[53][17] ;
 wire \w[53][18] ;
 wire \w[53][19] ;
 wire \w[53][1] ;
 wire \w[53][20] ;
 wire \w[53][21] ;
 wire \w[53][22] ;
 wire \w[53][23] ;
 wire \w[53][24] ;
 wire \w[53][25] ;
 wire \w[53][26] ;
 wire \w[53][27] ;
 wire \w[53][28] ;
 wire \w[53][29] ;
 wire \w[53][2] ;
 wire \w[53][30] ;
 wire \w[53][31] ;
 wire \w[53][3] ;
 wire \w[53][4] ;
 wire \w[53][5] ;
 wire \w[53][6] ;
 wire \w[53][7] ;
 wire \w[53][8] ;
 wire \w[53][9] ;
 wire \w[54][0] ;
 wire \w[54][10] ;
 wire \w[54][11] ;
 wire \w[54][12] ;
 wire \w[54][13] ;
 wire \w[54][14] ;
 wire \w[54][15] ;
 wire \w[54][16] ;
 wire \w[54][17] ;
 wire \w[54][18] ;
 wire \w[54][19] ;
 wire \w[54][1] ;
 wire \w[54][20] ;
 wire \w[54][21] ;
 wire \w[54][22] ;
 wire \w[54][23] ;
 wire \w[54][24] ;
 wire \w[54][25] ;
 wire \w[54][26] ;
 wire \w[54][27] ;
 wire \w[54][28] ;
 wire \w[54][29] ;
 wire \w[54][2] ;
 wire \w[54][30] ;
 wire \w[54][31] ;
 wire \w[54][3] ;
 wire \w[54][4] ;
 wire \w[54][5] ;
 wire \w[54][6] ;
 wire \w[54][7] ;
 wire \w[54][8] ;
 wire \w[54][9] ;
 wire \w[55][0] ;
 wire \w[55][10] ;
 wire \w[55][11] ;
 wire \w[55][12] ;
 wire \w[55][13] ;
 wire \w[55][14] ;
 wire \w[55][15] ;
 wire \w[55][16] ;
 wire \w[55][17] ;
 wire \w[55][18] ;
 wire \w[55][19] ;
 wire \w[55][1] ;
 wire \w[55][20] ;
 wire \w[55][21] ;
 wire \w[55][22] ;
 wire \w[55][23] ;
 wire \w[55][24] ;
 wire \w[55][25] ;
 wire \w[55][26] ;
 wire \w[55][27] ;
 wire \w[55][28] ;
 wire \w[55][29] ;
 wire \w[55][2] ;
 wire \w[55][30] ;
 wire \w[55][31] ;
 wire \w[55][3] ;
 wire \w[55][4] ;
 wire \w[55][5] ;
 wire \w[55][6] ;
 wire \w[55][7] ;
 wire \w[55][8] ;
 wire \w[55][9] ;
 wire \w[56][0] ;
 wire \w[56][10] ;
 wire \w[56][11] ;
 wire \w[56][12] ;
 wire \w[56][13] ;
 wire \w[56][14] ;
 wire \w[56][15] ;
 wire \w[56][16] ;
 wire \w[56][17] ;
 wire \w[56][18] ;
 wire \w[56][19] ;
 wire \w[56][1] ;
 wire \w[56][20] ;
 wire \w[56][21] ;
 wire \w[56][22] ;
 wire \w[56][23] ;
 wire \w[56][24] ;
 wire \w[56][25] ;
 wire \w[56][26] ;
 wire \w[56][27] ;
 wire \w[56][28] ;
 wire \w[56][29] ;
 wire \w[56][2] ;
 wire \w[56][30] ;
 wire \w[56][31] ;
 wire \w[56][3] ;
 wire \w[56][4] ;
 wire \w[56][5] ;
 wire \w[56][6] ;
 wire \w[56][7] ;
 wire \w[56][8] ;
 wire \w[56][9] ;
 wire \w[57][0] ;
 wire \w[57][10] ;
 wire \w[57][11] ;
 wire \w[57][12] ;
 wire \w[57][13] ;
 wire \w[57][14] ;
 wire \w[57][15] ;
 wire \w[57][16] ;
 wire \w[57][17] ;
 wire \w[57][18] ;
 wire \w[57][19] ;
 wire \w[57][1] ;
 wire \w[57][20] ;
 wire \w[57][21] ;
 wire \w[57][22] ;
 wire \w[57][23] ;
 wire \w[57][24] ;
 wire \w[57][25] ;
 wire \w[57][26] ;
 wire \w[57][27] ;
 wire \w[57][28] ;
 wire \w[57][29] ;
 wire \w[57][2] ;
 wire \w[57][30] ;
 wire \w[57][31] ;
 wire \w[57][3] ;
 wire \w[57][4] ;
 wire \w[57][5] ;
 wire \w[57][6] ;
 wire \w[57][7] ;
 wire \w[57][8] ;
 wire \w[57][9] ;
 wire \w[58][0] ;
 wire \w[58][10] ;
 wire \w[58][11] ;
 wire \w[58][12] ;
 wire \w[58][13] ;
 wire \w[58][14] ;
 wire \w[58][15] ;
 wire \w[58][16] ;
 wire \w[58][17] ;
 wire \w[58][18] ;
 wire \w[58][19] ;
 wire \w[58][1] ;
 wire \w[58][20] ;
 wire \w[58][21] ;
 wire \w[58][22] ;
 wire \w[58][23] ;
 wire \w[58][24] ;
 wire \w[58][25] ;
 wire \w[58][26] ;
 wire \w[58][27] ;
 wire \w[58][28] ;
 wire \w[58][29] ;
 wire \w[58][2] ;
 wire \w[58][30] ;
 wire \w[58][31] ;
 wire \w[58][3] ;
 wire \w[58][4] ;
 wire \w[58][5] ;
 wire \w[58][6] ;
 wire \w[58][7] ;
 wire \w[58][8] ;
 wire \w[58][9] ;
 wire \w[59][0] ;
 wire \w[59][10] ;
 wire \w[59][11] ;
 wire \w[59][12] ;
 wire \w[59][13] ;
 wire \w[59][14] ;
 wire \w[59][15] ;
 wire \w[59][16] ;
 wire \w[59][17] ;
 wire \w[59][18] ;
 wire \w[59][19] ;
 wire \w[59][1] ;
 wire \w[59][20] ;
 wire \w[59][21] ;
 wire \w[59][22] ;
 wire \w[59][23] ;
 wire \w[59][24] ;
 wire \w[59][25] ;
 wire \w[59][26] ;
 wire \w[59][27] ;
 wire \w[59][28] ;
 wire \w[59][29] ;
 wire \w[59][2] ;
 wire \w[59][30] ;
 wire \w[59][31] ;
 wire \w[59][3] ;
 wire \w[59][4] ;
 wire \w[59][5] ;
 wire \w[59][6] ;
 wire \w[59][7] ;
 wire \w[59][8] ;
 wire \w[59][9] ;
 wire \w[5][0] ;
 wire \w[5][10] ;
 wire \w[5][11] ;
 wire \w[5][12] ;
 wire \w[5][13] ;
 wire \w[5][14] ;
 wire \w[5][15] ;
 wire \w[5][16] ;
 wire \w[5][17] ;
 wire \w[5][18] ;
 wire \w[5][19] ;
 wire \w[5][1] ;
 wire \w[5][20] ;
 wire \w[5][21] ;
 wire \w[5][22] ;
 wire \w[5][23] ;
 wire \w[5][24] ;
 wire \w[5][25] ;
 wire \w[5][26] ;
 wire \w[5][27] ;
 wire \w[5][28] ;
 wire \w[5][29] ;
 wire \w[5][2] ;
 wire \w[5][30] ;
 wire \w[5][31] ;
 wire \w[5][3] ;
 wire \w[5][4] ;
 wire \w[5][5] ;
 wire \w[5][6] ;
 wire \w[5][7] ;
 wire \w[5][8] ;
 wire \w[5][9] ;
 wire \w[60][0] ;
 wire \w[60][10] ;
 wire \w[60][11] ;
 wire \w[60][12] ;
 wire \w[60][13] ;
 wire \w[60][14] ;
 wire \w[60][15] ;
 wire \w[60][16] ;
 wire \w[60][17] ;
 wire \w[60][18] ;
 wire \w[60][19] ;
 wire \w[60][1] ;
 wire \w[60][20] ;
 wire \w[60][21] ;
 wire \w[60][22] ;
 wire \w[60][23] ;
 wire \w[60][24] ;
 wire \w[60][25] ;
 wire \w[60][26] ;
 wire \w[60][27] ;
 wire \w[60][28] ;
 wire \w[60][29] ;
 wire \w[60][2] ;
 wire \w[60][30] ;
 wire \w[60][31] ;
 wire \w[60][3] ;
 wire \w[60][4] ;
 wire \w[60][5] ;
 wire \w[60][6] ;
 wire \w[60][7] ;
 wire \w[60][8] ;
 wire \w[60][9] ;
 wire \w[61][0] ;
 wire \w[61][10] ;
 wire \w[61][11] ;
 wire \w[61][12] ;
 wire \w[61][13] ;
 wire \w[61][14] ;
 wire \w[61][15] ;
 wire \w[61][16] ;
 wire \w[61][17] ;
 wire \w[61][18] ;
 wire \w[61][19] ;
 wire \w[61][1] ;
 wire \w[61][20] ;
 wire \w[61][21] ;
 wire \w[61][22] ;
 wire \w[61][23] ;
 wire \w[61][24] ;
 wire \w[61][25] ;
 wire \w[61][26] ;
 wire \w[61][27] ;
 wire \w[61][28] ;
 wire \w[61][29] ;
 wire \w[61][2] ;
 wire \w[61][30] ;
 wire \w[61][31] ;
 wire \w[61][3] ;
 wire \w[61][4] ;
 wire \w[61][5] ;
 wire \w[61][6] ;
 wire \w[61][7] ;
 wire \w[61][8] ;
 wire \w[61][9] ;
 wire \w[62][0] ;
 wire \w[62][10] ;
 wire \w[62][11] ;
 wire \w[62][12] ;
 wire \w[62][13] ;
 wire \w[62][14] ;
 wire \w[62][15] ;
 wire \w[62][16] ;
 wire \w[62][17] ;
 wire \w[62][18] ;
 wire \w[62][19] ;
 wire \w[62][1] ;
 wire \w[62][20] ;
 wire \w[62][21] ;
 wire \w[62][22] ;
 wire \w[62][23] ;
 wire \w[62][24] ;
 wire \w[62][25] ;
 wire \w[62][26] ;
 wire \w[62][27] ;
 wire \w[62][28] ;
 wire \w[62][29] ;
 wire \w[62][2] ;
 wire \w[62][30] ;
 wire \w[62][31] ;
 wire \w[62][3] ;
 wire \w[62][4] ;
 wire \w[62][5] ;
 wire \w[62][6] ;
 wire \w[62][7] ;
 wire \w[62][8] ;
 wire \w[62][9] ;
 wire \w[63][0] ;
 wire \w[63][10] ;
 wire \w[63][11] ;
 wire \w[63][12] ;
 wire \w[63][13] ;
 wire \w[63][14] ;
 wire \w[63][15] ;
 wire \w[63][16] ;
 wire \w[63][17] ;
 wire \w[63][18] ;
 wire \w[63][19] ;
 wire \w[63][1] ;
 wire \w[63][20] ;
 wire \w[63][21] ;
 wire \w[63][22] ;
 wire \w[63][23] ;
 wire \w[63][24] ;
 wire \w[63][25] ;
 wire \w[63][26] ;
 wire \w[63][27] ;
 wire \w[63][28] ;
 wire \w[63][29] ;
 wire \w[63][2] ;
 wire \w[63][30] ;
 wire \w[63][31] ;
 wire \w[63][3] ;
 wire \w[63][4] ;
 wire \w[63][5] ;
 wire \w[63][6] ;
 wire \w[63][7] ;
 wire \w[63][8] ;
 wire \w[63][9] ;
 wire \w[6][0] ;
 wire \w[6][10] ;
 wire \w[6][11] ;
 wire \w[6][12] ;
 wire \w[6][13] ;
 wire \w[6][14] ;
 wire \w[6][15] ;
 wire \w[6][16] ;
 wire \w[6][17] ;
 wire \w[6][18] ;
 wire \w[6][19] ;
 wire \w[6][1] ;
 wire \w[6][20] ;
 wire \w[6][21] ;
 wire \w[6][22] ;
 wire \w[6][23] ;
 wire \w[6][24] ;
 wire \w[6][25] ;
 wire \w[6][26] ;
 wire \w[6][27] ;
 wire \w[6][28] ;
 wire \w[6][29] ;
 wire \w[6][2] ;
 wire \w[6][30] ;
 wire \w[6][31] ;
 wire \w[6][3] ;
 wire \w[6][4] ;
 wire \w[6][5] ;
 wire \w[6][6] ;
 wire \w[6][7] ;
 wire \w[6][8] ;
 wire \w[6][9] ;
 wire \w[7][0] ;
 wire \w[7][10] ;
 wire \w[7][11] ;
 wire \w[7][12] ;
 wire \w[7][13] ;
 wire \w[7][14] ;
 wire \w[7][15] ;
 wire \w[7][16] ;
 wire \w[7][17] ;
 wire \w[7][18] ;
 wire \w[7][19] ;
 wire \w[7][1] ;
 wire \w[7][20] ;
 wire \w[7][21] ;
 wire \w[7][22] ;
 wire \w[7][23] ;
 wire \w[7][24] ;
 wire \w[7][25] ;
 wire \w[7][26] ;
 wire \w[7][27] ;
 wire \w[7][28] ;
 wire \w[7][29] ;
 wire \w[7][2] ;
 wire \w[7][30] ;
 wire \w[7][31] ;
 wire \w[7][3] ;
 wire \w[7][4] ;
 wire \w[7][5] ;
 wire \w[7][6] ;
 wire \w[7][7] ;
 wire \w[7][8] ;
 wire \w[7][9] ;
 wire \w[8][0] ;
 wire \w[8][10] ;
 wire \w[8][11] ;
 wire \w[8][12] ;
 wire \w[8][13] ;
 wire \w[8][14] ;
 wire \w[8][15] ;
 wire \w[8][16] ;
 wire \w[8][17] ;
 wire \w[8][18] ;
 wire \w[8][19] ;
 wire \w[8][1] ;
 wire \w[8][20] ;
 wire \w[8][21] ;
 wire \w[8][22] ;
 wire \w[8][23] ;
 wire \w[8][24] ;
 wire \w[8][25] ;
 wire \w[8][26] ;
 wire \w[8][27] ;
 wire \w[8][28] ;
 wire \w[8][29] ;
 wire \w[8][2] ;
 wire \w[8][30] ;
 wire \w[8][31] ;
 wire \w[8][3] ;
 wire \w[8][4] ;
 wire \w[8][5] ;
 wire \w[8][6] ;
 wire \w[8][7] ;
 wire \w[8][8] ;
 wire \w[8][9] ;
 wire \w[9][0] ;
 wire \w[9][10] ;
 wire \w[9][11] ;
 wire \w[9][12] ;
 wire \w[9][13] ;
 wire \w[9][14] ;
 wire \w[9][15] ;
 wire \w[9][16] ;
 wire \w[9][17] ;
 wire \w[9][18] ;
 wire \w[9][19] ;
 wire \w[9][1] ;
 wire \w[9][20] ;
 wire \w[9][21] ;
 wire \w[9][22] ;
 wire \w[9][23] ;
 wire \w[9][24] ;
 wire \w[9][25] ;
 wire \w[9][26] ;
 wire \w[9][27] ;
 wire \w[9][28] ;
 wire \w[9][29] ;
 wire \w[9][2] ;
 wire \w[9][30] ;
 wire \w[9][31] ;
 wire \w[9][3] ;
 wire \w[9][4] ;
 wire \w[9][5] ;
 wire \w[9][6] ;
 wire \w[9][7] ;
 wire \w[9][8] ;
 wire \w[9][9] ;
 wire net1170;

 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1475 ();
 sky130_fd_sc_hd__mux4_1 _14381_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03855_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1474 ();
 sky130_fd_sc_hd__mux4_1 _14383_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03857_));
 sky130_fd_sc_hd__mux4_1 _14384_ (.A0(_03851_),
    .A1(_03853_),
    .A2(_03855_),
    .A3(_03857_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_03858_));
 sky130_fd_sc_hd__mux2i_4 _14385_ (.A0(_03849_),
    .A1(_03858_),
    .S(net630),
    .Y(_12083_));
 sky130_fd_sc_hd__mux4_1 _14386_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03859_));
 sky130_fd_sc_hd__mux4_1 _14387_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03860_));
 sky130_fd_sc_hd__mux4_1 _14388_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03861_));
 sky130_fd_sc_hd__mux4_1 _14389_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03862_));
 sky130_fd_sc_hd__mux4_2 _14390_ (.A0(_03859_),
    .A1(_03860_),
    .A2(_03861_),
    .A3(_03862_),
    .S0(net596),
    .S1(net595),
    .X(_03863_));
 sky130_fd_sc_hd__mux4_1 _14391_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03864_));
 sky130_fd_sc_hd__mux4_1 _14392_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03865_));
 sky130_fd_sc_hd__mux4_1 _14393_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03866_));
 sky130_fd_sc_hd__mux4_1 _14394_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net602),
    .S1(net605),
    .X(_03867_));
 sky130_fd_sc_hd__mux4_1 _14395_ (.A0(_03864_),
    .A1(_03865_),
    .A2(_03866_),
    .A3(_03867_),
    .S0(net596),
    .S1(net595),
    .X(_03868_));
 sky130_fd_sc_hd__mux2i_4 _14396_ (.A0(_03863_),
    .A1(_03868_),
    .S(net593),
    .Y(_03869_));
 sky130_fd_sc_hd__xnor2_1 _14397_ (.A(_03739_),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__xnor2_1 _14398_ (.A(_03259_),
    .B(_03870_),
    .Y(_12088_));
 sky130_fd_sc_hd__mux4_1 _14399_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net673),
    .S1(net680),
    .X(_03871_));
 sky130_fd_sc_hd__mux4_1 _14400_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net673),
    .S1(net680),
    .X(_03872_));
 sky130_fd_sc_hd__mux4_1 _14401_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net673),
    .S1(net680),
    .X(_03873_));
 sky130_fd_sc_hd__mux4_1 _14402_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net673),
    .S1(net680),
    .X(_03874_));
 sky130_fd_sc_hd__mux4_4 _14403_ (.A0(_03871_),
    .A1(_03872_),
    .A2(_03873_),
    .A3(_03874_),
    .S0(net669),
    .S1(net667),
    .X(_03875_));
 sky130_fd_sc_hd__mux4_1 _14404_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net672),
    .S1(\count15_2[1] ),
    .X(_03876_));
 sky130_fd_sc_hd__mux4_1 _14405_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net672),
    .S1(\count15_2[1] ),
    .X(_03877_));
 sky130_fd_sc_hd__mux4_1 _14406_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net672),
    .S1(\count15_2[1] ),
    .X(_03878_));
 sky130_fd_sc_hd__mux4_1 _14407_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net672),
    .S1(\count15_2[1] ),
    .X(_03879_));
 sky130_fd_sc_hd__mux4_1 _14408_ (.A0(_03876_),
    .A1(_03877_),
    .A2(_03878_),
    .A3(_03879_),
    .S0(net671),
    .S1(net668),
    .X(_03880_));
 sky130_fd_sc_hd__mux2i_4 _14409_ (.A0(_03875_),
    .A1(_03880_),
    .S(net665),
    .Y(_03881_));
 sky130_fd_sc_hd__xnor2_1 _14410_ (.A(_03643_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__xnor2_2 _14411_ (.A(_03053_),
    .B(_03882_),
    .Y(_12087_));
 sky130_fd_sc_hd__mux4_1 _14412_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net560),
    .S1(net570),
    .X(_03883_));
 sky130_fd_sc_hd__mux4_1 _14413_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net560),
    .S1(net570),
    .X(_03884_));
 sky130_fd_sc_hd__mux4_1 _14414_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net560),
    .S1(net570),
    .X(_03885_));
 sky130_fd_sc_hd__mux4_1 _14415_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net560),
    .S1(net570),
    .X(_03886_));
 sky130_fd_sc_hd__mux4_4 _14416_ (.A0(_03883_),
    .A1(_03884_),
    .A2(_03885_),
    .A3(_03886_),
    .S0(net557),
    .S1(net555),
    .X(_03887_));
 sky130_fd_sc_hd__mux4_1 _14417_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net560),
    .S1(net569),
    .X(_03888_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1473 ();
 sky130_fd_sc_hd__mux4_1 _14419_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net560),
    .S1(net569),
    .X(_03890_));
 sky130_fd_sc_hd__mux4_1 _14420_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net560),
    .S1(net569),
    .X(_03891_));
 sky130_fd_sc_hd__mux4_1 _14421_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net560),
    .S1(net569),
    .X(_03892_));
 sky130_fd_sc_hd__mux4_1 _14422_ (.A0(_03888_),
    .A1(_03890_),
    .A2(_03891_),
    .A3(_03892_),
    .S0(net557),
    .S1(net555),
    .X(_03893_));
 sky130_fd_sc_hd__mux2i_4 _14423_ (.A0(_03887_),
    .A1(_03893_),
    .S(net553),
    .Y(_12086_));
 sky130_fd_sc_hd__mux4_1 _14424_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net640),
    .S1(net642),
    .X(_03894_));
 sky130_fd_sc_hd__mux4_1 _14425_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net640),
    .S1(net642),
    .X(_03895_));
 sky130_fd_sc_hd__mux4_1 _14426_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net640),
    .S1(net642),
    .X(_03896_));
 sky130_fd_sc_hd__mux4_1 _14427_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net640),
    .S1(net642),
    .X(_03897_));
 sky130_fd_sc_hd__mux4_2 _14428_ (.A0(_03894_),
    .A1(_03895_),
    .A2(_03896_),
    .A3(_03897_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_03898_));
 sky130_fd_sc_hd__mux4_1 _14429_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net640),
    .S1(net642),
    .X(_03899_));
 sky130_fd_sc_hd__mux4_1 _14430_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_03900_));
 sky130_fd_sc_hd__mux4_1 _14431_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_03901_));
 sky130_fd_sc_hd__mux4_1 _14432_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_03902_));
 sky130_fd_sc_hd__mux4_1 _14433_ (.A0(_03899_),
    .A1(_03900_),
    .A2(_03901_),
    .A3(_03902_),
    .S0(net634),
    .S1(net632),
    .X(_03903_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1472 ();
 sky130_fd_sc_hd__mux2i_2 _14435_ (.A0(_03898_),
    .A1(_03903_),
    .S(net630),
    .Y(_12091_));
 sky130_fd_sc_hd__mux4_1 _14436_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net603),
    .S1(net607),
    .X(_03905_));
 sky130_fd_sc_hd__mux4_1 _14437_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net603),
    .S1(net607),
    .X(_03906_));
 sky130_fd_sc_hd__mux4_1 _14438_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net603),
    .S1(net607),
    .X(_03907_));
 sky130_fd_sc_hd__mux4_1 _14439_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net603),
    .S1(net607),
    .X(_03908_));
 sky130_fd_sc_hd__mux4_4 _14440_ (.A0(_03905_),
    .A1(_03906_),
    .A2(_03907_),
    .A3(_03908_),
    .S0(net596),
    .S1(net595),
    .X(_03909_));
 sky130_fd_sc_hd__mux4_1 _14441_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net603),
    .S1(net605),
    .X(_03910_));
 sky130_fd_sc_hd__mux4_1 _14442_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net603),
    .S1(net605),
    .X(_03911_));
 sky130_fd_sc_hd__mux4_1 _14443_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net603),
    .S1(net605),
    .X(_03912_));
 sky130_fd_sc_hd__mux4_1 _14444_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net603),
    .S1(net605),
    .X(_03913_));
 sky130_fd_sc_hd__mux4_1 _14445_ (.A0(_03910_),
    .A1(_03911_),
    .A2(_03912_),
    .A3(_03913_),
    .S0(net596),
    .S1(net595),
    .X(_03914_));
 sky130_fd_sc_hd__mux2i_4 _14446_ (.A0(_03909_),
    .A1(_03914_),
    .S(net593),
    .Y(_03915_));
 sky130_fd_sc_hd__xnor2_1 _14447_ (.A(_03805_),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__xnor2_1 _14448_ (.A(_03340_),
    .B(_03916_),
    .Y(_12096_));
 sky130_fd_sc_hd__mux4_1 _14449_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03917_));
 sky130_fd_sc_hd__mux4_1 _14450_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03918_));
 sky130_fd_sc_hd__mux4_1 _14451_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03919_));
 sky130_fd_sc_hd__mux4_1 _14452_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03920_));
 sky130_fd_sc_hd__mux4_4 _14453_ (.A0(_03917_),
    .A1(_03918_),
    .A2(_03919_),
    .A3(_03920_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03921_));
 sky130_fd_sc_hd__mux4_1 _14454_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net674),
    .S1(net678),
    .X(_03922_));
 sky130_fd_sc_hd__mux4_1 _14455_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net674),
    .S1(net678),
    .X(_03923_));
 sky130_fd_sc_hd__mux4_1 _14456_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net674),
    .S1(net678),
    .X(_03924_));
 sky130_fd_sc_hd__mux4_1 _14457_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net674),
    .S1(net678),
    .X(_03925_));
 sky130_fd_sc_hd__mux4_1 _14458_ (.A0(_03922_),
    .A1(_03923_),
    .A2(_03924_),
    .A3(_03925_),
    .S0(net669),
    .S1(net667),
    .X(_03926_));
 sky130_fd_sc_hd__mux2i_4 _14459_ (.A0(_03921_),
    .A1(_03926_),
    .S(net666),
    .Y(_03927_));
 sky130_fd_sc_hd__xnor2_2 _14460_ (.A(_03691_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__xnor2_4 _14461_ (.A(_03174_),
    .B(_03928_),
    .Y(_12095_));
 sky130_fd_sc_hd__mux4_1 _14462_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net561),
    .S1(net572),
    .X(_03929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1471 ();
 sky130_fd_sc_hd__mux4_1 _14464_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net561),
    .S1(net572),
    .X(_03931_));
 sky130_fd_sc_hd__mux4_1 _14465_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net561),
    .S1(net572),
    .X(_03932_));
 sky130_fd_sc_hd__mux4_1 _14466_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net561),
    .S1(net572),
    .X(_03933_));
 sky130_fd_sc_hd__mux4_4 _14467_ (.A0(_03929_),
    .A1(_03931_),
    .A2(_03932_),
    .A3(_03933_),
    .S0(net559),
    .S1(net555),
    .X(_03934_));
 sky130_fd_sc_hd__mux4_1 _14468_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net561),
    .S1(net572),
    .X(_03935_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1470 ();
 sky130_fd_sc_hd__mux4_1 _14470_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net566),
    .S1(net572),
    .X(_03937_));
 sky130_fd_sc_hd__mux4_1 _14471_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net561),
    .S1(net572),
    .X(_03938_));
 sky130_fd_sc_hd__mux4_1 _14472_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net566),
    .S1(net571),
    .X(_03939_));
 sky130_fd_sc_hd__mux4_1 _14473_ (.A0(_03935_),
    .A1(_03937_),
    .A2(_03938_),
    .A3(_03939_),
    .S0(net559),
    .S1(net555),
    .X(_03940_));
 sky130_fd_sc_hd__mux2i_4 _14474_ (.A0(_03934_),
    .A1(_03940_),
    .S(net553),
    .Y(_12094_));
 sky130_fd_sc_hd__mux4_1 _14475_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net636),
    .S1(net646),
    .X(_03941_));
 sky130_fd_sc_hd__mux4_1 _14476_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net636),
    .S1(net647),
    .X(_03942_));
 sky130_fd_sc_hd__mux4_1 _14477_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net636),
    .S1(net646),
    .X(_03943_));
 sky130_fd_sc_hd__mux4_1 _14478_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net636),
    .S1(net646),
    .X(_03944_));
 sky130_fd_sc_hd__mux4_4 _14479_ (.A0(_03941_),
    .A1(_03942_),
    .A2(_03943_),
    .A3(_03944_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03945_));
 sky130_fd_sc_hd__mux4_1 _14480_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net638),
    .S1(net645),
    .X(_03946_));
 sky130_fd_sc_hd__mux4_1 _14481_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net637),
    .S1(net645),
    .X(_03947_));
 sky130_fd_sc_hd__mux4_1 _14482_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net637),
    .S1(net645),
    .X(_03948_));
 sky130_fd_sc_hd__mux4_1 _14483_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net639),
    .S1(net645),
    .X(_03949_));
 sky130_fd_sc_hd__mux4_1 _14484_ (.A0(_03946_),
    .A1(_03947_),
    .A2(_03948_),
    .A3(_03949_),
    .S0(net633),
    .S1(net631),
    .X(_03950_));
 sky130_fd_sc_hd__mux2i_4 _14485_ (.A0(_03945_),
    .A1(_03950_),
    .S(net629),
    .Y(_12099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1468 ();
 sky130_fd_sc_hd__mux4_1 _14488_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03953_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1466 ();
 sky130_fd_sc_hd__mux4_1 _14491_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03956_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1464 ();
 sky130_fd_sc_hd__mux4_1 _14494_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1462 ();
 sky130_fd_sc_hd__mux4_1 _14497_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03962_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1460 ();
 sky130_fd_sc_hd__mux4_4 _14500_ (.A0(_03953_),
    .A1(_03956_),
    .A2(_03959_),
    .A3(_03962_),
    .S0(net597),
    .S1(net594),
    .X(_03965_));
 sky130_fd_sc_hd__mux4_1 _14501_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03966_));
 sky130_fd_sc_hd__mux4_1 _14502_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03967_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1458 ();
 sky130_fd_sc_hd__mux4_1 _14505_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1456 ();
 sky130_fd_sc_hd__mux4_1 _14508_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_03973_));
 sky130_fd_sc_hd__mux4_1 _14509_ (.A0(_03966_),
    .A1(_03967_),
    .A2(_03970_),
    .A3(_03973_),
    .S0(net597),
    .S1(net594),
    .X(_03974_));
 sky130_fd_sc_hd__mux2i_4 _14510_ (.A0(_03965_),
    .A1(_03974_),
    .S(net592),
    .Y(_03975_));
 sky130_fd_sc_hd__xnor2_1 _14511_ (.A(_03869_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__xnor2_1 _14512_ (.A(_03411_),
    .B(_03976_),
    .Y(_12104_));
 sky130_fd_sc_hd__mux4_1 _14513_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net675),
    .S1(net681),
    .X(_03977_));
 sky130_fd_sc_hd__mux4_1 _14514_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net675),
    .S1(net681),
    .X(_03978_));
 sky130_fd_sc_hd__mux4_1 _14515_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net675),
    .S1(net681),
    .X(_03979_));
 sky130_fd_sc_hd__mux4_1 _14516_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net675),
    .S1(net681),
    .X(_03980_));
 sky130_fd_sc_hd__mux4_4 _14517_ (.A0(_03977_),
    .A1(_03978_),
    .A2(_03979_),
    .A3(_03980_),
    .S0(net670),
    .S1(net668),
    .X(_03981_));
 sky130_fd_sc_hd__mux4_2 _14518_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net676),
    .S1(net682),
    .X(_03982_));
 sky130_fd_sc_hd__mux4_1 _14519_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net675),
    .S1(net681),
    .X(_03983_));
 sky130_fd_sc_hd__mux4_1 _14520_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net675),
    .S1(net681),
    .X(_03984_));
 sky130_fd_sc_hd__mux4_1 _14521_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net675),
    .S1(net681),
    .X(_03985_));
 sky130_fd_sc_hd__mux4_1 _14522_ (.A0(_03982_),
    .A1(_03983_),
    .A2(_03984_),
    .A3(_03985_),
    .S0(net671),
    .S1(net668),
    .X(_03986_));
 sky130_fd_sc_hd__mux2i_4 _14523_ (.A0(_03981_),
    .A1(_03986_),
    .S(net665),
    .Y(_03987_));
 sky130_fd_sc_hd__xnor2_2 _14524_ (.A(_03762_),
    .B(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__xnor2_4 _14525_ (.A(_03284_),
    .B(_03988_),
    .Y(_12103_));
 sky130_fd_sc_hd__mux4_1 _14526_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1455 ();
 sky130_fd_sc_hd__mux4_1 _14528_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03991_));
 sky130_fd_sc_hd__mux4_1 _14529_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03992_));
 sky130_fd_sc_hd__mux4_1 _14530_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03993_));
 sky130_fd_sc_hd__mux4_2 _14531_ (.A0(_03989_),
    .A1(_03991_),
    .A2(_03992_),
    .A3(_03993_),
    .S0(net558),
    .S1(net556),
    .X(_03994_));
 sky130_fd_sc_hd__mux4_1 _14532_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03995_));
 sky130_fd_sc_hd__mux4_1 _14533_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03996_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1454 ();
 sky130_fd_sc_hd__mux4_1 _14535_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03998_));
 sky130_fd_sc_hd__mux4_1 _14536_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net563),
    .S1(net568),
    .X(_03999_));
 sky130_fd_sc_hd__mux4_1 _14537_ (.A0(_03995_),
    .A1(_03996_),
    .A2(_03998_),
    .A3(_03999_),
    .S0(net558),
    .S1(net556),
    .X(_04000_));
 sky130_fd_sc_hd__mux2i_4 _14538_ (.A0(_03994_),
    .A1(_04000_),
    .S(net554),
    .Y(_12102_));
 sky130_fd_sc_hd__mux4_1 _14539_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net640),
    .S1(net645),
    .X(_04001_));
 sky130_fd_sc_hd__mux4_1 _14540_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net640),
    .S1(net645),
    .X(_04002_));
 sky130_fd_sc_hd__mux4_1 _14541_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net640),
    .S1(net645),
    .X(_04003_));
 sky130_fd_sc_hd__mux4_1 _14542_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net640),
    .S1(net645),
    .X(_04004_));
 sky130_fd_sc_hd__mux4_4 _14543_ (.A0(_04001_),
    .A1(_04002_),
    .A2(_04003_),
    .A3(_04004_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04005_));
 sky130_fd_sc_hd__mux4_1 _14544_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net640),
    .S1(net642),
    .X(_04006_));
 sky130_fd_sc_hd__mux4_1 _14545_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net640),
    .S1(net642),
    .X(_04007_));
 sky130_fd_sc_hd__mux4_1 _14546_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net640),
    .S1(net642),
    .X(_04008_));
 sky130_fd_sc_hd__mux4_1 _14547_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net640),
    .S1(net642),
    .X(_04009_));
 sky130_fd_sc_hd__mux4_1 _14548_ (.A0(_04006_),
    .A1(_04007_),
    .A2(_04008_),
    .A3(_04009_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04010_));
 sky130_fd_sc_hd__mux2i_4 _14549_ (.A0(_04005_),
    .A1(_04010_),
    .S(net630),
    .Y(_12107_));
 sky130_fd_sc_hd__mux4_1 _14550_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04011_));
 sky130_fd_sc_hd__mux4_1 _14551_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04012_));
 sky130_fd_sc_hd__mux4_1 _14552_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04013_));
 sky130_fd_sc_hd__mux4_1 _14553_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04014_));
 sky130_fd_sc_hd__mux4_4 _14554_ (.A0(_04011_),
    .A1(_04012_),
    .A2(_04013_),
    .A3(_04014_),
    .S0(net597),
    .S1(net594),
    .X(_04015_));
 sky130_fd_sc_hd__mux4_1 _14555_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04016_));
 sky130_fd_sc_hd__mux4_1 _14556_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04017_));
 sky130_fd_sc_hd__mux4_1 _14557_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04018_));
 sky130_fd_sc_hd__mux4_1 _14558_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04019_));
 sky130_fd_sc_hd__mux4_1 _14559_ (.A0(_04016_),
    .A1(_04017_),
    .A2(_04018_),
    .A3(_04019_),
    .S0(net597),
    .S1(net594),
    .X(_04020_));
 sky130_fd_sc_hd__mux2i_4 _14560_ (.A0(_04015_),
    .A1(_04020_),
    .S(net592),
    .Y(_04021_));
 sky130_fd_sc_hd__xnor2_1 _14561_ (.A(_03915_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__xnor2_1 _14562_ (.A(_03492_),
    .B(_04022_),
    .Y(_12112_));
 sky130_fd_sc_hd__mux4_1 _14563_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04023_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1453 ();
 sky130_fd_sc_hd__mux4_1 _14565_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1451 ();
 sky130_fd_sc_hd__mux4_1 _14568_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04028_));
 sky130_fd_sc_hd__mux4_1 _14569_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04029_));
 sky130_fd_sc_hd__mux4_4 _14570_ (.A0(_04023_),
    .A1(_04025_),
    .A2(_04028_),
    .A3(_04029_),
    .S0(net669),
    .S1(net667),
    .X(_04030_));
 sky130_fd_sc_hd__mux4_1 _14571_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04031_));
 sky130_fd_sc_hd__mux4_1 _14572_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04032_));
 sky130_fd_sc_hd__mux4_1 _14573_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04033_));
 sky130_fd_sc_hd__mux4_1 _14574_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net673),
    .S1(net680),
    .X(_04034_));
 sky130_fd_sc_hd__mux4_1 _14575_ (.A0(_04031_),
    .A1(_04032_),
    .A2(_04033_),
    .A3(_04034_),
    .S0(net669),
    .S1(net667),
    .X(_04035_));
 sky130_fd_sc_hd__mux2i_4 _14576_ (.A0(_04030_),
    .A1(_04035_),
    .S(net666),
    .Y(_04036_));
 sky130_fd_sc_hd__xnor2_2 _14577_ (.A(_03817_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__xnor2_4 _14578_ (.A(_03353_),
    .B(_04037_),
    .Y(_12111_));
 sky130_fd_sc_hd__mux4_1 _14579_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04038_));
 sky130_fd_sc_hd__mux4_1 _14580_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04039_));
 sky130_fd_sc_hd__mux4_1 _14581_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04040_));
 sky130_fd_sc_hd__mux4_1 _14582_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04041_));
 sky130_fd_sc_hd__mux4_2 _14583_ (.A0(_04038_),
    .A1(_04039_),
    .A2(_04040_),
    .A3(_04041_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_04042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1450 ();
 sky130_fd_sc_hd__mux4_1 _14585_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04044_));
 sky130_fd_sc_hd__mux4_1 _14586_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1449 ();
 sky130_fd_sc_hd__mux4_1 _14588_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04047_));
 sky130_fd_sc_hd__mux4_1 _14589_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04048_));
 sky130_fd_sc_hd__mux4_1 _14590_ (.A0(_04044_),
    .A1(_04045_),
    .A2(_04047_),
    .A3(_04048_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_04049_));
 sky130_fd_sc_hd__mux2i_4 _14591_ (.A0(_04042_),
    .A1(_04049_),
    .S(\count7_2[5] ),
    .Y(_12110_));
 sky130_fd_sc_hd__mux4_1 _14592_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net636),
    .S1(net646),
    .X(_04050_));
 sky130_fd_sc_hd__mux4_1 _14593_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net636),
    .S1(net646),
    .X(_04051_));
 sky130_fd_sc_hd__mux4_1 _14594_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net636),
    .S1(net646),
    .X(_04052_));
 sky130_fd_sc_hd__mux4_1 _14595_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net636),
    .S1(net646),
    .X(_04053_));
 sky130_fd_sc_hd__mux4_2 _14596_ (.A0(_04050_),
    .A1(_04051_),
    .A2(_04052_),
    .A3(_04053_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04054_));
 sky130_fd_sc_hd__mux4_1 _14597_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net639),
    .S1(net647),
    .X(_04055_));
 sky130_fd_sc_hd__mux4_1 _14598_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net639),
    .S1(net647),
    .X(_04056_));
 sky130_fd_sc_hd__mux4_1 _14599_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net639),
    .S1(net647),
    .X(_04057_));
 sky130_fd_sc_hd__mux4_1 _14600_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net639),
    .S1(net647),
    .X(_04058_));
 sky130_fd_sc_hd__mux4_1 _14601_ (.A0(_04055_),
    .A1(_04056_),
    .A2(_04057_),
    .A3(_04058_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04059_));
 sky130_fd_sc_hd__mux2i_4 _14602_ (.A0(_04054_),
    .A1(_04059_),
    .S(\count16_2[5] ),
    .Y(_12115_));
 sky130_fd_sc_hd__mux4_1 _14603_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04060_));
 sky130_fd_sc_hd__mux4_1 _14604_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04061_));
 sky130_fd_sc_hd__mux4_1 _14605_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04062_));
 sky130_fd_sc_hd__mux4_1 _14606_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04063_));
 sky130_fd_sc_hd__mux4_4 _14607_ (.A0(_04060_),
    .A1(_04061_),
    .A2(_04062_),
    .A3(_04063_),
    .S0(net598),
    .S1(net594),
    .X(_04064_));
 sky130_fd_sc_hd__mux4_1 _14608_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04065_));
 sky130_fd_sc_hd__mux4_1 _14609_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04066_));
 sky130_fd_sc_hd__mux4_1 _14610_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04067_));
 sky130_fd_sc_hd__mux4_1 _14611_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net599),
    .S1(net606),
    .X(_04068_));
 sky130_fd_sc_hd__mux4_1 _14612_ (.A0(_04065_),
    .A1(_04066_),
    .A2(_04067_),
    .A3(_04068_),
    .S0(net598),
    .S1(net594),
    .X(_04069_));
 sky130_fd_sc_hd__mux2i_4 _14613_ (.A0(_04064_),
    .A1(_04069_),
    .S(net592),
    .Y(_04070_));
 sky130_fd_sc_hd__xnor2_1 _14614_ (.A(_03975_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__xnor2_1 _14615_ (.A(_03562_),
    .B(_04071_),
    .Y(_12120_));
 sky130_fd_sc_hd__mux4_1 _14616_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net672),
    .S1(net679),
    .X(_04072_));
 sky130_fd_sc_hd__mux4_1 _14617_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net672),
    .S1(net679),
    .X(_04073_));
 sky130_fd_sc_hd__mux4_1 _14618_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net672),
    .S1(net679),
    .X(_04074_));
 sky130_fd_sc_hd__mux4_1 _14619_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net672),
    .S1(net679),
    .X(_04075_));
 sky130_fd_sc_hd__mux4_4 _14620_ (.A0(_04072_),
    .A1(_04073_),
    .A2(_04074_),
    .A3(_04075_),
    .S0(net669),
    .S1(net667),
    .X(_04076_));
 sky130_fd_sc_hd__mux4_1 _14621_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net677),
    .S1(\count15_2[1] ),
    .X(_04077_));
 sky130_fd_sc_hd__mux4_1 _14622_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net677),
    .S1(\count15_2[1] ),
    .X(_04078_));
 sky130_fd_sc_hd__mux4_1 _14623_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net677),
    .S1(\count15_2[1] ),
    .X(_04079_));
 sky130_fd_sc_hd__mux4_1 _14624_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net677),
    .S1(\count15_2[1] ),
    .X(_04080_));
 sky130_fd_sc_hd__mux4_1 _14625_ (.A0(_04077_),
    .A1(_04078_),
    .A2(_04079_),
    .A3(_04080_),
    .S0(net671),
    .S1(net668),
    .X(_04081_));
 sky130_fd_sc_hd__mux2i_4 _14626_ (.A0(_04076_),
    .A1(_04081_),
    .S(net665),
    .Y(_04082_));
 sky130_fd_sc_hd__xnor2_4 _14627_ (.A(_03436_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__xnor2_4 _14628_ (.A(_03053_),
    .B(_04083_),
    .Y(_12119_));
 sky130_fd_sc_hd__mux4_1 _14629_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04084_));
 sky130_fd_sc_hd__mux4_1 _14630_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1448 ();
 sky130_fd_sc_hd__mux4_1 _14632_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04087_));
 sky130_fd_sc_hd__mux4_1 _14633_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04088_));
 sky130_fd_sc_hd__mux4_4 _14634_ (.A0(_04084_),
    .A1(_04085_),
    .A2(_04087_),
    .A3(_04088_),
    .S0(net559),
    .S1(\count7_2[4] ),
    .X(_04089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1447 ();
 sky130_fd_sc_hd__mux4_1 _14636_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04091_));
 sky130_fd_sc_hd__mux4_1 _14637_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04092_));
 sky130_fd_sc_hd__mux4_1 _14638_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04093_));
 sky130_fd_sc_hd__mux4_1 _14639_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net562),
    .S1(net567),
    .X(_04094_));
 sky130_fd_sc_hd__mux4_1 _14640_ (.A0(_04091_),
    .A1(_04092_),
    .A2(_04093_),
    .A3(_04094_),
    .S0(net559),
    .S1(\count7_2[4] ),
    .X(_04095_));
 sky130_fd_sc_hd__mux2i_4 _14641_ (.A0(_04089_),
    .A1(_04095_),
    .S(\count7_2[5] ),
    .Y(_12118_));
 sky130_fd_sc_hd__mux4_1 _14642_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net636),
    .S1(net646),
    .X(_04096_));
 sky130_fd_sc_hd__mux4_1 _14643_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net636),
    .S1(net647),
    .X(_04097_));
 sky130_fd_sc_hd__mux4_1 _14644_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net636),
    .S1(net646),
    .X(_04098_));
 sky130_fd_sc_hd__mux4_1 _14645_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net636),
    .S1(net646),
    .X(_04099_));
 sky130_fd_sc_hd__mux4_2 _14646_ (.A0(_04096_),
    .A1(_04097_),
    .A2(_04098_),
    .A3(_04099_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04100_));
 sky130_fd_sc_hd__mux4_1 _14647_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net639),
    .S1(net643),
    .X(_04101_));
 sky130_fd_sc_hd__mux4_1 _14648_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net639),
    .S1(net647),
    .X(_04102_));
 sky130_fd_sc_hd__mux4_1 _14649_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net639),
    .S1(net647),
    .X(_04103_));
 sky130_fd_sc_hd__mux4_1 _14650_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net639),
    .S1(net647),
    .X(_04104_));
 sky130_fd_sc_hd__mux4_1 _14651_ (.A0(_04101_),
    .A1(_04102_),
    .A2(_04103_),
    .A3(_04104_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04105_));
 sky130_fd_sc_hd__mux2i_4 _14652_ (.A0(_04100_),
    .A1(_04105_),
    .S(\count16_2[5] ),
    .Y(_12123_));
 sky130_fd_sc_hd__mux4_1 _14653_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04106_));
 sky130_fd_sc_hd__mux4_1 _14654_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04107_));
 sky130_fd_sc_hd__mux4_1 _14655_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04108_));
 sky130_fd_sc_hd__mux4_1 _14656_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net601),
    .S1(net608),
    .X(_04109_));
 sky130_fd_sc_hd__mux4_4 _14657_ (.A0(_04106_),
    .A1(_04107_),
    .A2(_04108_),
    .A3(_04109_),
    .S0(net597),
    .S1(net594),
    .X(_04110_));
 sky130_fd_sc_hd__mux4_1 _14658_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net599),
    .S1(net606),
    .X(_04111_));
 sky130_fd_sc_hd__mux4_1 _14659_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net600),
    .S1(net607),
    .X(_04112_));
 sky130_fd_sc_hd__mux4_1 _14660_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04113_));
 sky130_fd_sc_hd__mux4_1 _14661_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net600),
    .S1(net607),
    .X(_04114_));
 sky130_fd_sc_hd__mux4_1 _14662_ (.A0(_04111_),
    .A1(_04112_),
    .A2(_04113_),
    .A3(_04114_),
    .S0(net598),
    .S1(net594),
    .X(_04115_));
 sky130_fd_sc_hd__mux2i_4 _14663_ (.A0(_04110_),
    .A1(_04115_),
    .S(net592),
    .Y(_04116_));
 sky130_fd_sc_hd__xnor2_1 _14664_ (.A(_04021_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__xnor2_1 _14665_ (.A(_03620_),
    .B(_04117_),
    .Y(_12128_));
 sky130_fd_sc_hd__mux4_1 _14666_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net672),
    .S1(net679),
    .X(_04118_));
 sky130_fd_sc_hd__mux4_1 _14667_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net672),
    .S1(net679),
    .X(_04119_));
 sky130_fd_sc_hd__mux4_1 _14668_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net672),
    .S1(net679),
    .X(_04120_));
 sky130_fd_sc_hd__mux4_1 _14669_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net672),
    .S1(net679),
    .X(_04121_));
 sky130_fd_sc_hd__mux4_4 _14670_ (.A0(_04118_),
    .A1(_04119_),
    .A2(_04120_),
    .A3(_04121_),
    .S0(net669),
    .S1(net667),
    .X(_04122_));
 sky130_fd_sc_hd__mux4_1 _14671_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net677),
    .S1(net679),
    .X(_04123_));
 sky130_fd_sc_hd__mux4_1 _14672_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net677),
    .S1(net679),
    .X(_04124_));
 sky130_fd_sc_hd__mux4_1 _14673_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net677),
    .S1(net679),
    .X(_04125_));
 sky130_fd_sc_hd__mux4_1 _14674_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net677),
    .S1(net679),
    .X(_04126_));
 sky130_fd_sc_hd__mux4_1 _14675_ (.A0(_04123_),
    .A1(_04124_),
    .A2(_04125_),
    .A3(_04126_),
    .S0(net671),
    .S1(net668),
    .X(_04127_));
 sky130_fd_sc_hd__mux2i_4 _14676_ (.A0(_04122_),
    .A1(_04127_),
    .S(net665),
    .Y(_04128_));
 sky130_fd_sc_hd__xnor2_4 _14677_ (.A(_03517_),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__xnor2_4 _14678_ (.A(_03174_),
    .B(_04129_),
    .Y(_12127_));
 sky130_fd_sc_hd__mux4_1 _14679_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net560),
    .S1(net570),
    .X(_04130_));
 sky130_fd_sc_hd__mux4_1 _14680_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net560),
    .S1(net570),
    .X(_04131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1446 ();
 sky130_fd_sc_hd__mux4_1 _14682_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net560),
    .S1(net570),
    .X(_04133_));
 sky130_fd_sc_hd__mux4_1 _14683_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net560),
    .S1(net570),
    .X(_04134_));
 sky130_fd_sc_hd__mux4_2 _14684_ (.A0(_04130_),
    .A1(_04131_),
    .A2(_04133_),
    .A3(_04134_),
    .S0(net557),
    .S1(net555),
    .X(_04135_));
 sky130_fd_sc_hd__mux4_1 _14685_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net560),
    .S1(net569),
    .X(_04136_));
 sky130_fd_sc_hd__mux4_1 _14686_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net560),
    .S1(net569),
    .X(_04137_));
 sky130_fd_sc_hd__mux4_1 _14687_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net560),
    .S1(net569),
    .X(_04138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1445 ();
 sky130_fd_sc_hd__mux4_1 _14689_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net560),
    .S1(net569),
    .X(_04140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1444 ();
 sky130_fd_sc_hd__mux4_1 _14691_ (.A0(_04136_),
    .A1(_04137_),
    .A2(_04138_),
    .A3(_04140_),
    .S0(net557),
    .S1(net555),
    .X(_04142_));
 sky130_fd_sc_hd__mux2i_4 _14692_ (.A0(_04135_),
    .A1(_04142_),
    .S(net553),
    .Y(_12126_));
 sky130_fd_sc_hd__mux4_1 _14693_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net636),
    .S1(net646),
    .X(_04143_));
 sky130_fd_sc_hd__mux4_1 _14694_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net636),
    .S1(net647),
    .X(_04144_));
 sky130_fd_sc_hd__mux4_1 _14695_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net636),
    .S1(net646),
    .X(_04145_));
 sky130_fd_sc_hd__mux4_1 _14696_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net636),
    .S1(net646),
    .X(_04146_));
 sky130_fd_sc_hd__mux4_4 _14697_ (.A0(_04143_),
    .A1(_04144_),
    .A2(_04145_),
    .A3(_04146_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04147_));
 sky130_fd_sc_hd__mux4_1 _14698_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net639),
    .S1(net647),
    .X(_04148_));
 sky130_fd_sc_hd__mux4_1 _14699_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net639),
    .S1(net647),
    .X(_04149_));
 sky130_fd_sc_hd__mux4_1 _14700_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net639),
    .S1(net647),
    .X(_04150_));
 sky130_fd_sc_hd__mux4_1 _14701_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net639),
    .S1(net647),
    .X(_04151_));
 sky130_fd_sc_hd__mux4_1 _14702_ (.A0(_04148_),
    .A1(_04149_),
    .A2(_04150_),
    .A3(_04151_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04152_));
 sky130_fd_sc_hd__mux2i_4 _14703_ (.A0(_04147_),
    .A1(_04152_),
    .S(\count16_2[5] ),
    .Y(_12131_));
 sky130_fd_sc_hd__mux4_1 _14704_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net601),
    .S1(net608),
    .X(_04153_));
 sky130_fd_sc_hd__mux4_1 _14705_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net601),
    .S1(net608),
    .X(_04154_));
 sky130_fd_sc_hd__mux4_1 _14706_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04155_));
 sky130_fd_sc_hd__mux4_1 _14707_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net601),
    .S1(net608),
    .X(_04156_));
 sky130_fd_sc_hd__mux4_4 _14708_ (.A0(_04153_),
    .A1(_04154_),
    .A2(_04155_),
    .A3(_04156_),
    .S0(net597),
    .S1(net594),
    .X(_04157_));
 sky130_fd_sc_hd__mux4_1 _14709_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_04158_));
 sky130_fd_sc_hd__mux4_1 _14710_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_04159_));
 sky130_fd_sc_hd__mux4_1 _14711_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04160_));
 sky130_fd_sc_hd__mux4_1 _14712_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(\count2_2[2] ),
    .S1(net608),
    .X(_04161_));
 sky130_fd_sc_hd__mux4_1 _14713_ (.A0(_04158_),
    .A1(_04159_),
    .A2(_04160_),
    .A3(_04161_),
    .S0(net597),
    .S1(net594),
    .X(_04162_));
 sky130_fd_sc_hd__mux2i_4 _14714_ (.A0(_04157_),
    .A1(_04162_),
    .S(net592),
    .Y(_04163_));
 sky130_fd_sc_hd__xnor2_1 _14715_ (.A(_04070_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__xnor2_1 _14716_ (.A(_03679_),
    .B(_04164_),
    .Y(_12136_));
 sky130_fd_sc_hd__xnor2_1 _14717_ (.A(_03284_),
    .B(_03574_),
    .Y(_04165_));
 sky130_fd_sc_hd__xnor2_2 _14718_ (.A(_02995_),
    .B(_04165_),
    .Y(_12135_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1443 ();
 sky130_fd_sc_hd__mux4_1 _14720_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net563),
    .S1(net568),
    .X(_04167_));
 sky130_fd_sc_hd__mux4_1 _14721_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net563),
    .S1(net568),
    .X(_04168_));
 sky130_fd_sc_hd__mux4_1 _14722_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net563),
    .S1(net568),
    .X(_04169_));
 sky130_fd_sc_hd__mux4_1 _14723_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net563),
    .S1(net568),
    .X(_04170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1442 ();
 sky130_fd_sc_hd__mux4_4 _14725_ (.A0(_04167_),
    .A1(_04168_),
    .A2(_04169_),
    .A3(_04170_),
    .S0(net558),
    .S1(net556),
    .X(_04172_));
 sky130_fd_sc_hd__mux4_1 _14726_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net565),
    .S1(net568),
    .X(_04173_));
 sky130_fd_sc_hd__mux4_1 _14727_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net565),
    .S1(net568),
    .X(_04174_));
 sky130_fd_sc_hd__mux4_1 _14728_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net565),
    .S1(net569),
    .X(_04175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1441 ();
 sky130_fd_sc_hd__mux4_1 _14730_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net565),
    .S1(net569),
    .X(_04177_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1440 ();
 sky130_fd_sc_hd__mux4_1 _14732_ (.A0(_04173_),
    .A1(_04174_),
    .A2(_04175_),
    .A3(_04177_),
    .S0(net558),
    .S1(net556),
    .X(_04179_));
 sky130_fd_sc_hd__mux2i_4 _14733_ (.A0(_04172_),
    .A1(_04179_),
    .S(net554),
    .Y(_12134_));
 sky130_fd_sc_hd__mux4_1 _14734_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net636),
    .S1(net646),
    .X(_04180_));
 sky130_fd_sc_hd__mux4_1 _14735_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net636),
    .S1(net646),
    .X(_04181_));
 sky130_fd_sc_hd__mux4_1 _14736_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net636),
    .S1(net646),
    .X(_04182_));
 sky130_fd_sc_hd__mux4_1 _14737_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net636),
    .S1(net646),
    .X(_04183_));
 sky130_fd_sc_hd__mux4_4 _14738_ (.A0(_04180_),
    .A1(_04181_),
    .A2(_04182_),
    .A3(_04183_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04184_));
 sky130_fd_sc_hd__mux4_1 _14739_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net639),
    .S1(net647),
    .X(_04185_));
 sky130_fd_sc_hd__mux4_1 _14740_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net639),
    .S1(net647),
    .X(_04186_));
 sky130_fd_sc_hd__mux4_1 _14741_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net639),
    .S1(net647),
    .X(_04187_));
 sky130_fd_sc_hd__mux4_1 _14742_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net639),
    .S1(net647),
    .X(_04188_));
 sky130_fd_sc_hd__mux4_1 _14743_ (.A0(_04185_),
    .A1(_04186_),
    .A2(_04187_),
    .A3(_04188_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04189_));
 sky130_fd_sc_hd__mux2i_4 _14744_ (.A0(_04184_),
    .A1(_04189_),
    .S(\count16_2[5] ),
    .Y(_12139_));
 sky130_fd_sc_hd__mux4_1 _14745_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net601),
    .S1(net608),
    .X(_04190_));
 sky130_fd_sc_hd__mux4_1 _14746_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net601),
    .S1(net608),
    .X(_04191_));
 sky130_fd_sc_hd__mux4_1 _14747_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net601),
    .S1(net608),
    .X(_04192_));
 sky130_fd_sc_hd__mux4_1 _14748_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net601),
    .S1(net608),
    .X(_04193_));
 sky130_fd_sc_hd__mux4_4 _14749_ (.A0(_04190_),
    .A1(_04191_),
    .A2(_04192_),
    .A3(_04193_),
    .S0(net597),
    .S1(net594),
    .X(_04194_));
 sky130_fd_sc_hd__mux4_1 _14750_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net599),
    .S1(net606),
    .X(_04195_));
 sky130_fd_sc_hd__mux4_1 _14751_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04196_));
 sky130_fd_sc_hd__mux4_1 _14752_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04197_));
 sky130_fd_sc_hd__mux4_1 _14753_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_04198_));
 sky130_fd_sc_hd__mux4_1 _14754_ (.A0(_04195_),
    .A1(_04196_),
    .A2(_04197_),
    .A3(_04198_),
    .S0(net597),
    .S1(net594),
    .X(_04199_));
 sky130_fd_sc_hd__mux2i_4 _14755_ (.A0(_04194_),
    .A1(_04199_),
    .S(net592),
    .Y(_04200_));
 sky130_fd_sc_hd__xnor2_1 _14756_ (.A(_04116_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__xnor2_1 _14757_ (.A(_03739_),
    .B(_04201_),
    .Y(_12144_));
 sky130_fd_sc_hd__xnor2_1 _14758_ (.A(_03353_),
    .B(_03632_),
    .Y(_04202_));
 sky130_fd_sc_hd__xnor2_2 _14759_ (.A(_03147_),
    .B(_04202_),
    .Y(_12143_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1439 ();
 sky130_fd_sc_hd__mux4_1 _14761_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04204_));
 sky130_fd_sc_hd__mux4_1 _14762_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04205_));
 sky130_fd_sc_hd__mux4_1 _14763_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04206_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1438 ();
 sky130_fd_sc_hd__mux4_1 _14765_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1437 ();
 sky130_fd_sc_hd__mux4_2 _14767_ (.A0(_04204_),
    .A1(_04205_),
    .A2(_04206_),
    .A3(_04208_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_04210_));
 sky130_fd_sc_hd__mux4_1 _14768_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04211_));
 sky130_fd_sc_hd__mux4_1 _14769_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04212_));
 sky130_fd_sc_hd__mux4_1 _14770_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04213_));
 sky130_fd_sc_hd__mux4_1 _14771_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04214_));
 sky130_fd_sc_hd__mux4_1 _14772_ (.A0(_04211_),
    .A1(_04212_),
    .A2(_04213_),
    .A3(_04214_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_04215_));
 sky130_fd_sc_hd__mux2i_4 _14773_ (.A0(_04210_),
    .A1(_04215_),
    .S(\count7_2[5] ),
    .Y(_12142_));
 sky130_fd_sc_hd__mux4_1 _14774_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net635),
    .S1(net644),
    .X(_04216_));
 sky130_fd_sc_hd__mux4_1 _14775_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net635),
    .S1(net644),
    .X(_04217_));
 sky130_fd_sc_hd__mux4_1 _14776_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net635),
    .S1(net644),
    .X(_04218_));
 sky130_fd_sc_hd__mux4_1 _14777_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net635),
    .S1(net644),
    .X(_04219_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1436 ();
 sky130_fd_sc_hd__mux4_4 _14779_ (.A0(_04216_),
    .A1(_04217_),
    .A2(_04218_),
    .A3(_04219_),
    .S0(net633),
    .S1(net632),
    .X(_04221_));
 sky130_fd_sc_hd__mux4_1 _14780_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net638),
    .S1(net645),
    .X(_04222_));
 sky130_fd_sc_hd__mux4_1 _14781_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net638),
    .S1(net645),
    .X(_04223_));
 sky130_fd_sc_hd__mux4_1 _14782_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net638),
    .S1(net645),
    .X(_04224_));
 sky130_fd_sc_hd__mux4_1 _14783_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net638),
    .S1(net645),
    .X(_04225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1435 ();
 sky130_fd_sc_hd__mux4_1 _14785_ (.A0(_04222_),
    .A1(_04223_),
    .A2(_04224_),
    .A3(_04225_),
    .S0(net634),
    .S1(net632),
    .X(_04227_));
 sky130_fd_sc_hd__mux2i_4 _14786_ (.A0(_04221_),
    .A1(_04227_),
    .S(net630),
    .Y(_12147_));
 sky130_fd_sc_hd__mux4_1 _14787_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net603),
    .S1(net605),
    .X(_04228_));
 sky130_fd_sc_hd__mux4_1 _14788_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net603),
    .S1(net605),
    .X(_04229_));
 sky130_fd_sc_hd__mux4_1 _14789_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net603),
    .S1(net605),
    .X(_04230_));
 sky130_fd_sc_hd__mux4_1 _14790_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net603),
    .S1(net605),
    .X(_04231_));
 sky130_fd_sc_hd__mux4_4 _14791_ (.A0(_04228_),
    .A1(_04229_),
    .A2(_04230_),
    .A3(_04231_),
    .S0(net596),
    .S1(net595),
    .X(_04232_));
 sky130_fd_sc_hd__mux4_1 _14792_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net600),
    .S1(net607),
    .X(_04233_));
 sky130_fd_sc_hd__mux4_1 _14793_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net600),
    .S1(net607),
    .X(_04234_));
 sky130_fd_sc_hd__mux4_1 _14794_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net600),
    .S1(net607),
    .X(_04235_));
 sky130_fd_sc_hd__mux4_1 _14795_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net600),
    .S1(net607),
    .X(_04236_));
 sky130_fd_sc_hd__mux4_1 _14796_ (.A0(_04233_),
    .A1(_04234_),
    .A2(_04235_),
    .A3(_04236_),
    .S0(net596),
    .S1(net595),
    .X(_04237_));
 sky130_fd_sc_hd__mux2i_4 _14797_ (.A0(_04232_),
    .A1(_04237_),
    .S(net593),
    .Y(_04238_));
 sky130_fd_sc_hd__xnor2_1 _14798_ (.A(_04163_),
    .B(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__xnor2_1 _14799_ (.A(_03805_),
    .B(_04239_),
    .Y(_12152_));
 sky130_fd_sc_hd__xnor2_1 _14800_ (.A(_03436_),
    .B(_03702_),
    .Y(_04240_));
 sky130_fd_sc_hd__xnor2_2 _14801_ (.A(_03271_),
    .B(_04240_),
    .Y(_12151_));
 sky130_fd_sc_hd__mux4_1 _14802_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04241_));
 sky130_fd_sc_hd__mux4_1 _14803_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04242_));
 sky130_fd_sc_hd__mux4_1 _14804_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04243_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1434 ();
 sky130_fd_sc_hd__mux4_1 _14806_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04245_));
 sky130_fd_sc_hd__mux4_2 _14807_ (.A0(_04241_),
    .A1(_04242_),
    .A2(_04243_),
    .A3(_04245_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_04246_));
 sky130_fd_sc_hd__mux4_1 _14808_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net562),
    .S1(net567),
    .X(_04247_));
 sky130_fd_sc_hd__mux4_1 _14809_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net562),
    .S1(net567),
    .X(_04248_));
 sky130_fd_sc_hd__mux4_1 _14810_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net562),
    .S1(net567),
    .X(_04249_));
 sky130_fd_sc_hd__mux4_1 _14811_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net562),
    .S1(net567),
    .X(_04250_));
 sky130_fd_sc_hd__mux4_1 _14812_ (.A0(_04247_),
    .A1(_04248_),
    .A2(_04249_),
    .A3(_04250_),
    .S0(net559),
    .S1(\count7_2[4] ),
    .X(_04251_));
 sky130_fd_sc_hd__mux2i_4 _14813_ (.A0(_04246_),
    .A1(_04251_),
    .S(\count7_2[5] ),
    .Y(_12150_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1433 ();
 sky130_fd_sc_hd__mux4_1 _14815_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net635),
    .S1(net644),
    .X(_04253_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1432 ();
 sky130_fd_sc_hd__mux4_1 _14817_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net635),
    .S1(net644),
    .X(_04255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1431 ();
 sky130_fd_sc_hd__mux4_1 _14819_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net635),
    .S1(net644),
    .X(_04257_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1430 ();
 sky130_fd_sc_hd__mux4_1 _14821_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net635),
    .S1(net644),
    .X(_04259_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1429 ();
 sky130_fd_sc_hd__mux4_4 _14823_ (.A0(_04253_),
    .A1(_04255_),
    .A2(_04257_),
    .A3(_04259_),
    .S0(net634),
    .S1(net632),
    .X(_04261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1428 ();
 sky130_fd_sc_hd__mux4_1 _14825_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04263_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1427 ();
 sky130_fd_sc_hd__mux4_1 _14827_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04265_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1426 ();
 sky130_fd_sc_hd__mux4_1 _14829_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1425 ();
 sky130_fd_sc_hd__mux4_1 _14831_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04269_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1424 ();
 sky130_fd_sc_hd__mux4_1 _14833_ (.A0(_04263_),
    .A1(_04265_),
    .A2(_04267_),
    .A3(_04269_),
    .S0(\count16_2[3] ),
    .S1(\count16_2[4] ),
    .X(_04271_));
 sky130_fd_sc_hd__mux2i_2 _14834_ (.A0(_04261_),
    .A1(_04271_),
    .S(net630),
    .Y(_12155_));
 sky130_fd_sc_hd__mux4_1 _14835_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net601),
    .S1(net608),
    .X(_04272_));
 sky130_fd_sc_hd__mux4_1 _14836_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net601),
    .S1(net608),
    .X(_04273_));
 sky130_fd_sc_hd__mux4_1 _14837_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net601),
    .S1(net608),
    .X(_04274_));
 sky130_fd_sc_hd__mux4_1 _14838_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net601),
    .S1(net608),
    .X(_04275_));
 sky130_fd_sc_hd__mux4_4 _14839_ (.A0(_04272_),
    .A1(_04273_),
    .A2(_04274_),
    .A3(_04275_),
    .S0(net597),
    .S1(net594),
    .X(_04276_));
 sky130_fd_sc_hd__mux4_1 _14840_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net599),
    .S1(net606),
    .X(_04277_));
 sky130_fd_sc_hd__mux4_1 _14841_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net599),
    .S1(net606),
    .X(_04278_));
 sky130_fd_sc_hd__mux4_1 _14842_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net599),
    .S1(net606),
    .X(_04279_));
 sky130_fd_sc_hd__mux4_1 _14843_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net599),
    .S1(net606),
    .X(_04280_));
 sky130_fd_sc_hd__mux4_1 _14844_ (.A0(_04277_),
    .A1(_04278_),
    .A2(_04279_),
    .A3(_04280_),
    .S0(net598),
    .S1(net594),
    .X(_04281_));
 sky130_fd_sc_hd__mux2i_4 _14845_ (.A0(_04276_),
    .A1(_04281_),
    .S(net592),
    .Y(_04282_));
 sky130_fd_sc_hd__xnor2_1 _14846_ (.A(_04200_),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__xnor2_2 _14847_ (.A(_03869_),
    .B(_04283_),
    .Y(_12160_));
 sky130_fd_sc_hd__xnor2_1 _14848_ (.A(_03517_),
    .B(_03751_),
    .Y(_04284_));
 sky130_fd_sc_hd__xnor2_2 _14849_ (.A(_03366_),
    .B(_04284_),
    .Y(_12159_));
 sky130_fd_sc_hd__mux4_1 _14850_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04285_));
 sky130_fd_sc_hd__mux4_1 _14851_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04286_));
 sky130_fd_sc_hd__mux4_1 _14852_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04287_));
 sky130_fd_sc_hd__mux4_1 _14853_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04288_));
 sky130_fd_sc_hd__mux4_4 _14854_ (.A0(_04285_),
    .A1(_04286_),
    .A2(_04287_),
    .A3(_04288_),
    .S0(net558),
    .S1(net556),
    .X(_04289_));
 sky130_fd_sc_hd__mux4_1 _14855_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04290_));
 sky130_fd_sc_hd__mux4_1 _14856_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04291_));
 sky130_fd_sc_hd__mux4_1 _14857_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04292_));
 sky130_fd_sc_hd__mux4_1 _14858_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net563),
    .S1(net568),
    .X(_04293_));
 sky130_fd_sc_hd__mux4_1 _14859_ (.A0(_04290_),
    .A1(_04291_),
    .A2(_04292_),
    .A3(_04293_),
    .S0(net558),
    .S1(net556),
    .X(_04294_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1423 ();
 sky130_fd_sc_hd__mux2i_4 _14861_ (.A0(_04289_),
    .A1(_04294_),
    .S(net554),
    .Y(_12158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1422 ();
 sky130_fd_sc_hd__mux4_1 _14863_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1421 ();
 sky130_fd_sc_hd__mux4_1 _14865_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1420 ();
 sky130_fd_sc_hd__mux4_1 _14867_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1419 ();
 sky130_fd_sc_hd__mux4_1 _14869_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04303_));
 sky130_fd_sc_hd__mux4_2 _14870_ (.A0(_04297_),
    .A1(_04299_),
    .A2(_04301_),
    .A3(_04303_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04304_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1418 ();
 sky130_fd_sc_hd__mux4_1 _14872_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04306_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1417 ();
 sky130_fd_sc_hd__mux4_1 _14874_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04308_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1416 ();
 sky130_fd_sc_hd__mux4_1 _14876_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04310_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1415 ();
 sky130_fd_sc_hd__mux4_1 _14878_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04312_));
 sky130_fd_sc_hd__mux4_1 _14879_ (.A0(_04306_),
    .A1(_04308_),
    .A2(_04310_),
    .A3(_04312_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04313_));
 sky130_fd_sc_hd__mux2i_4 _14880_ (.A0(_04304_),
    .A1(_04313_),
    .S(net630),
    .Y(_12163_));
 sky130_fd_sc_hd__mux4_1 _14881_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net599),
    .S1(net606),
    .X(_04314_));
 sky130_fd_sc_hd__mux4_1 _14882_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net599),
    .S1(net606),
    .X(_04315_));
 sky130_fd_sc_hd__mux4_1 _14883_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net599),
    .S1(net606),
    .X(_04316_));
 sky130_fd_sc_hd__mux4_1 _14884_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net599),
    .S1(net606),
    .X(_04317_));
 sky130_fd_sc_hd__mux4_4 _14885_ (.A0(_04314_),
    .A1(_04315_),
    .A2(_04316_),
    .A3(_04317_),
    .S0(net598),
    .S1(net595),
    .X(_04318_));
 sky130_fd_sc_hd__mux4_1 _14886_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net600),
    .S1(net607),
    .X(_04319_));
 sky130_fd_sc_hd__mux4_1 _14887_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net600),
    .S1(net607),
    .X(_04320_));
 sky130_fd_sc_hd__mux4_1 _14888_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net600),
    .S1(net607),
    .X(_04321_));
 sky130_fd_sc_hd__mux4_1 _14889_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net600),
    .S1(net607),
    .X(_04322_));
 sky130_fd_sc_hd__mux4_1 _14890_ (.A0(_04319_),
    .A1(_04320_),
    .A2(_04321_),
    .A3(_04322_),
    .S0(net598),
    .S1(net594),
    .X(_04323_));
 sky130_fd_sc_hd__mux2i_4 _14891_ (.A0(_04318_),
    .A1(_04323_),
    .S(net592),
    .Y(_04324_));
 sky130_fd_sc_hd__xnor2_1 _14892_ (.A(_04238_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__xnor2_1 _14893_ (.A(_03915_),
    .B(_04325_),
    .Y(_12168_));
 sky130_fd_sc_hd__xnor2_2 _14894_ (.A(_03574_),
    .B(_03828_),
    .Y(_04326_));
 sky130_fd_sc_hd__xnor2_4 _14895_ (.A(_03024_),
    .B(_04326_),
    .Y(_12167_));
 sky130_fd_sc_hd__mux4_1 _14896_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net561),
    .S1(net572),
    .X(_04327_));
 sky130_fd_sc_hd__mux4_1 _14897_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net561),
    .S1(net572),
    .X(_04328_));
 sky130_fd_sc_hd__mux4_1 _14898_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net561),
    .S1(net572),
    .X(_04329_));
 sky130_fd_sc_hd__mux4_1 _14899_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net561),
    .S1(net572),
    .X(_04330_));
 sky130_fd_sc_hd__mux4_4 _14900_ (.A0(_04327_),
    .A1(_04328_),
    .A2(_04329_),
    .A3(_04330_),
    .S0(net559),
    .S1(net555),
    .X(_04331_));
 sky130_fd_sc_hd__mux4_1 _14901_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net566),
    .S1(net571),
    .X(_04332_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1414 ();
 sky130_fd_sc_hd__mux4_1 _14903_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net566),
    .S1(net571),
    .X(_04334_));
 sky130_fd_sc_hd__mux4_1 _14904_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net566),
    .S1(net571),
    .X(_04335_));
 sky130_fd_sc_hd__mux4_1 _14905_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net566),
    .S1(net571),
    .X(_04336_));
 sky130_fd_sc_hd__mux4_1 _14906_ (.A0(_04332_),
    .A1(_04334_),
    .A2(_04335_),
    .A3(_04336_),
    .S0(net557),
    .S1(net555),
    .X(_04337_));
 sky130_fd_sc_hd__mux2i_4 _14907_ (.A0(_04331_),
    .A1(_04337_),
    .S(net553),
    .Y(_12166_));
 sky130_fd_sc_hd__mux4_1 _14908_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net635),
    .S1(net644),
    .X(_04338_));
 sky130_fd_sc_hd__mux4_1 _14909_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net635),
    .S1(net644),
    .X(_04339_));
 sky130_fd_sc_hd__mux4_1 _14910_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net635),
    .S1(net644),
    .X(_04340_));
 sky130_fd_sc_hd__mux4_1 _14911_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net635),
    .S1(net644),
    .X(_04341_));
 sky130_fd_sc_hd__mux4_4 _14912_ (.A0(_04338_),
    .A1(_04339_),
    .A2(_04340_),
    .A3(_04341_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04342_));
 sky130_fd_sc_hd__mux4_1 _14913_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04343_));
 sky130_fd_sc_hd__mux4_1 _14914_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04344_));
 sky130_fd_sc_hd__mux4_1 _14915_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04345_));
 sky130_fd_sc_hd__mux4_1 _14916_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(\count16_2[2] ),
    .S1(net642),
    .X(_04346_));
 sky130_fd_sc_hd__mux4_1 _14917_ (.A0(_04343_),
    .A1(_04344_),
    .A2(_04345_),
    .A3(_04346_),
    .S0(net634),
    .S1(net632),
    .X(_04347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1413 ();
 sky130_fd_sc_hd__mux2i_4 _14919_ (.A0(_04342_),
    .A1(_04347_),
    .S(net630),
    .Y(_12171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1412 ();
 sky130_fd_sc_hd__mux4_1 _14921_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04350_));
 sky130_fd_sc_hd__mux4_1 _14922_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04351_));
 sky130_fd_sc_hd__mux4_1 _14923_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04352_));
 sky130_fd_sc_hd__mux4_1 _14924_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04353_));
 sky130_fd_sc_hd__mux4_4 _14925_ (.A0(_04350_),
    .A1(_04351_),
    .A2(_04352_),
    .A3(_04353_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_04354_));
 sky130_fd_sc_hd__mux4_1 _14926_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04355_));
 sky130_fd_sc_hd__mux4_1 _14927_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04356_));
 sky130_fd_sc_hd__mux4_1 _14928_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04357_));
 sky130_fd_sc_hd__mux4_1 _14929_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net604),
    .S1(net609),
    .X(_04358_));
 sky130_fd_sc_hd__mux4_1 _14930_ (.A0(_04355_),
    .A1(_04356_),
    .A2(_04357_),
    .A3(_04358_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_04359_));
 sky130_fd_sc_hd__mux2i_4 _14931_ (.A0(_04354_),
    .A1(_04359_),
    .S(net593),
    .Y(_04360_));
 sky130_fd_sc_hd__xnor2_1 _14932_ (.A(_04282_),
    .B(_04360_),
    .Y(_12176_));
 sky130_fd_sc_hd__xnor2_1 _14933_ (.A(_03632_),
    .B(_03881_),
    .Y(_04361_));
 sky130_fd_sc_hd__xnor2_2 _14934_ (.A(_03163_),
    .B(_04361_),
    .Y(_12175_));
 sky130_fd_sc_hd__mux4_1 _14935_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net561),
    .S1(net572),
    .X(_04362_));
 sky130_fd_sc_hd__mux4_1 _14936_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net561),
    .S1(net572),
    .X(_04363_));
 sky130_fd_sc_hd__mux4_1 _14937_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net561),
    .S1(net572),
    .X(_04364_));
 sky130_fd_sc_hd__mux4_1 _14938_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net561),
    .S1(net572),
    .X(_04365_));
 sky130_fd_sc_hd__mux4_2 _14939_ (.A0(_04362_),
    .A1(_04363_),
    .A2(_04364_),
    .A3(_04365_),
    .S0(net559),
    .S1(net555),
    .X(_04366_));
 sky130_fd_sc_hd__mux4_1 _14940_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net566),
    .S1(net571),
    .X(_04367_));
 sky130_fd_sc_hd__mux4_1 _14941_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net566),
    .S1(net571),
    .X(_04368_));
 sky130_fd_sc_hd__mux4_1 _14942_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net566),
    .S1(net571),
    .X(_04369_));
 sky130_fd_sc_hd__mux4_1 _14943_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net566),
    .S1(net571),
    .X(_04370_));
 sky130_fd_sc_hd__mux4_1 _14944_ (.A0(_04367_),
    .A1(_04368_),
    .A2(_04369_),
    .A3(_04370_),
    .S0(net559),
    .S1(net555),
    .X(_04371_));
 sky130_fd_sc_hd__mux2i_4 _14945_ (.A0(_04366_),
    .A1(_04371_),
    .S(net553),
    .Y(_12174_));
 sky130_fd_sc_hd__mux4_1 _14946_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04372_));
 sky130_fd_sc_hd__mux4_1 _14947_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04373_));
 sky130_fd_sc_hd__mux4_1 _14948_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04374_));
 sky130_fd_sc_hd__mux4_1 _14949_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04375_));
 sky130_fd_sc_hd__mux4_4 _14950_ (.A0(_04372_),
    .A1(_04373_),
    .A2(_04374_),
    .A3(_04375_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04376_));
 sky130_fd_sc_hd__mux4_1 _14951_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04377_));
 sky130_fd_sc_hd__mux4_1 _14952_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04378_));
 sky130_fd_sc_hd__mux4_1 _14953_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04379_));
 sky130_fd_sc_hd__mux4_1 _14954_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net640),
    .S1(net645),
    .X(_04380_));
 sky130_fd_sc_hd__mux4_1 _14955_ (.A0(_04377_),
    .A1(_04378_),
    .A2(_04379_),
    .A3(_04380_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04381_));
 sky130_fd_sc_hd__mux2i_4 _14956_ (.A0(_04376_),
    .A1(_04381_),
    .S(net630),
    .Y(_12179_));
 sky130_fd_sc_hd__xnor2_1 _14957_ (.A(_02941_),
    .B(_04324_),
    .Y(_12184_));
 sky130_fd_sc_hd__xnor2_2 _14958_ (.A(_03702_),
    .B(_03927_),
    .Y(_04382_));
 sky130_fd_sc_hd__xnor2_4 _14959_ (.A(_03295_),
    .B(_04382_),
    .Y(_12183_));
 sky130_fd_sc_hd__mux4_1 _14960_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04383_));
 sky130_fd_sc_hd__mux4_1 _14961_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04384_));
 sky130_fd_sc_hd__mux4_1 _14962_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04385_));
 sky130_fd_sc_hd__mux4_1 _14963_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_04386_));
 sky130_fd_sc_hd__mux4_4 _14964_ (.A0(_04383_),
    .A1(_04384_),
    .A2(_04385_),
    .A3(_04386_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_04387_));
 sky130_fd_sc_hd__mux4_1 _14965_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net565),
    .S1(net572),
    .X(_04388_));
 sky130_fd_sc_hd__mux4_1 _14966_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net565),
    .S1(net572),
    .X(_04389_));
 sky130_fd_sc_hd__mux4_1 _14967_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net565),
    .S1(net572),
    .X(_04390_));
 sky130_fd_sc_hd__mux4_1 _14968_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net565),
    .S1(net572),
    .X(_04391_));
 sky130_fd_sc_hd__mux4_1 _14969_ (.A0(_04388_),
    .A1(_04389_),
    .A2(_04390_),
    .A3(_04391_),
    .S0(net558),
    .S1(net556),
    .X(_04392_));
 sky130_fd_sc_hd__mux2i_4 _14970_ (.A0(_04387_),
    .A1(_04392_),
    .S(net554),
    .Y(_12182_));
 sky130_fd_sc_hd__mux4_1 _14971_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net638),
    .S1(net643),
    .X(_04393_));
 sky130_fd_sc_hd__mux4_1 _14972_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net637),
    .S1(net643),
    .X(_04394_));
 sky130_fd_sc_hd__mux4_1 _14973_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net638),
    .S1(net643),
    .X(_04395_));
 sky130_fd_sc_hd__mux4_1 _14974_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net638),
    .S1(net643),
    .X(_04396_));
 sky130_fd_sc_hd__mux4_4 _14975_ (.A0(_04393_),
    .A1(_04394_),
    .A2(_04395_),
    .A3(_04396_),
    .S0(net633),
    .S1(net632),
    .X(_04397_));
 sky130_fd_sc_hd__mux4_1 _14976_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net635),
    .S1(net644),
    .X(_04398_));
 sky130_fd_sc_hd__mux4_1 _14977_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net635),
    .S1(net644),
    .X(_04399_));
 sky130_fd_sc_hd__mux4_1 _14978_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net638),
    .S1(net644),
    .X(_04400_));
 sky130_fd_sc_hd__mux4_1 _14979_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net638),
    .S1(net644),
    .X(_04401_));
 sky130_fd_sc_hd__mux4_1 _14980_ (.A0(_04398_),
    .A1(_04399_),
    .A2(_04400_),
    .A3(_04401_),
    .S0(net633),
    .S1(net632),
    .X(_04402_));
 sky130_fd_sc_hd__mux2i_4 _14981_ (.A0(_04397_),
    .A1(_04402_),
    .S(net629),
    .Y(_12187_));
 sky130_fd_sc_hd__xnor2_1 _14982_ (.A(_03109_),
    .B(_04360_),
    .Y(_12192_));
 sky130_fd_sc_hd__xnor2_1 _14983_ (.A(_03751_),
    .B(_03987_),
    .Y(_04403_));
 sky130_fd_sc_hd__xnor2_2 _14984_ (.A(_03377_),
    .B(_04403_),
    .Y(_12191_));
 sky130_fd_sc_hd__mux4_1 _14985_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net564),
    .S1(net568),
    .X(_04404_));
 sky130_fd_sc_hd__mux4_1 _14986_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net564),
    .S1(net568),
    .X(_04405_));
 sky130_fd_sc_hd__mux4_1 _14987_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net564),
    .S1(net568),
    .X(_04406_));
 sky130_fd_sc_hd__mux4_1 _14988_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net564),
    .S1(net568),
    .X(_04407_));
 sky130_fd_sc_hd__mux4_2 _14989_ (.A0(_04404_),
    .A1(_04405_),
    .A2(_04406_),
    .A3(_04407_),
    .S0(net558),
    .S1(net556),
    .X(_04408_));
 sky130_fd_sc_hd__mux4_1 _14990_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net564),
    .S1(net569),
    .X(_04409_));
 sky130_fd_sc_hd__mux4_1 _14991_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net564),
    .S1(net568),
    .X(_04410_));
 sky130_fd_sc_hd__mux4_1 _14992_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net564),
    .S1(net569),
    .X(_04411_));
 sky130_fd_sc_hd__mux4_1 _14993_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net564),
    .S1(net569),
    .X(_04412_));
 sky130_fd_sc_hd__mux4_1 _14994_ (.A0(_04409_),
    .A1(_04410_),
    .A2(_04411_),
    .A3(_04412_),
    .S0(net558),
    .S1(net556),
    .X(_04413_));
 sky130_fd_sc_hd__mux2i_4 _14995_ (.A0(_04408_),
    .A1(_04413_),
    .S(net554),
    .Y(_12190_));
 sky130_fd_sc_hd__mux4_1 _14996_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net636),
    .S1(net646),
    .X(_04414_));
 sky130_fd_sc_hd__mux4_1 _14997_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net636),
    .S1(net646),
    .X(_04415_));
 sky130_fd_sc_hd__mux4_1 _14998_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net636),
    .S1(net646),
    .X(_04416_));
 sky130_fd_sc_hd__mux4_1 _14999_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net636),
    .S1(net646),
    .X(_04417_));
 sky130_fd_sc_hd__mux4_4 _15000_ (.A0(_04414_),
    .A1(_04415_),
    .A2(_04416_),
    .A3(_04417_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_04418_));
 sky130_fd_sc_hd__mux4_1 _15001_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net637),
    .S1(net647),
    .X(_04419_));
 sky130_fd_sc_hd__mux4_1 _15002_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net637),
    .S1(net647),
    .X(_04420_));
 sky130_fd_sc_hd__mux4_1 _15003_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net637),
    .S1(net647),
    .X(_04421_));
 sky130_fd_sc_hd__mux4_1 _15004_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net637),
    .S1(net647),
    .X(_04422_));
 sky130_fd_sc_hd__mux4_1 _15005_ (.A0(_04419_),
    .A1(_04420_),
    .A2(_04421_),
    .A3(_04422_),
    .S0(net633),
    .S1(net631),
    .X(_04423_));
 sky130_fd_sc_hd__mux2i_4 _15006_ (.A0(_04418_),
    .A1(_04423_),
    .S(\count16_2[5] ),
    .Y(_12195_));
 sky130_fd_sc_hd__xnor2_1 _15007_ (.A(_02941_),
    .B(_03248_),
    .Y(_12200_));
 sky130_fd_sc_hd__xnor2_2 _15008_ (.A(_03828_),
    .B(_04036_),
    .Y(_04424_));
 sky130_fd_sc_hd__xnor2_4 _15009_ (.A(_03447_),
    .B(_04424_),
    .Y(_12199_));
 sky130_fd_sc_hd__mux4_1 _15010_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net560),
    .S1(net570),
    .X(_04425_));
 sky130_fd_sc_hd__mux4_1 _15011_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net560),
    .S1(net570),
    .X(_04426_));
 sky130_fd_sc_hd__mux4_1 _15012_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net560),
    .S1(net570),
    .X(_04427_));
 sky130_fd_sc_hd__mux4_1 _15013_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net560),
    .S1(net570),
    .X(_04428_));
 sky130_fd_sc_hd__mux4_4 _15014_ (.A0(_04425_),
    .A1(_04426_),
    .A2(_04427_),
    .A3(_04428_),
    .S0(net557),
    .S1(net555),
    .X(_04429_));
 sky130_fd_sc_hd__mux4_1 _15015_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net565),
    .S1(net571),
    .X(_04430_));
 sky130_fd_sc_hd__mux4_1 _15016_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net565),
    .S1(net571),
    .X(_04431_));
 sky130_fd_sc_hd__mux4_1 _15017_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net565),
    .S1(net571),
    .X(_04432_));
 sky130_fd_sc_hd__mux4_1 _15018_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net565),
    .S1(net571),
    .X(_04433_));
 sky130_fd_sc_hd__mux4_1 _15019_ (.A0(_04430_),
    .A1(_04431_),
    .A2(_04432_),
    .A3(_04433_),
    .S0(net558),
    .S1(net556),
    .X(_04434_));
 sky130_fd_sc_hd__mux2i_4 _15020_ (.A0(_04429_),
    .A1(_04434_),
    .S(net554),
    .Y(_12198_));
 sky130_fd_sc_hd__mux4_1 _15021_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net637),
    .S1(net646),
    .X(_04435_));
 sky130_fd_sc_hd__mux4_1 _15022_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net637),
    .S1(net646),
    .X(_04436_));
 sky130_fd_sc_hd__mux4_1 _15023_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net637),
    .S1(net646),
    .X(_04437_));
 sky130_fd_sc_hd__mux4_1 _15024_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net637),
    .S1(net646),
    .X(_04438_));
 sky130_fd_sc_hd__mux4_4 _15025_ (.A0(_04435_),
    .A1(_04436_),
    .A2(_04437_),
    .A3(_04438_),
    .S0(net633),
    .S1(net631),
    .X(_04439_));
 sky130_fd_sc_hd__mux4_1 _15026_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net637),
    .S1(net643),
    .X(_04440_));
 sky130_fd_sc_hd__mux4_1 _15027_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net637),
    .S1(net643),
    .X(_04441_));
 sky130_fd_sc_hd__mux4_1 _15028_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net637),
    .S1(net643),
    .X(_04442_));
 sky130_fd_sc_hd__mux4_1 _15029_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net637),
    .S1(net643),
    .X(_04443_));
 sky130_fd_sc_hd__mux4_1 _15030_ (.A0(_04440_),
    .A1(_04441_),
    .A2(_04442_),
    .A3(_04443_),
    .S0(net633),
    .S1(net631),
    .X(_04444_));
 sky130_fd_sc_hd__mux2i_4 _15031_ (.A0(_04439_),
    .A1(_04444_),
    .S(net629),
    .Y(_12203_));
 sky130_fd_sc_hd__xnor2_1 _15032_ (.A(_03109_),
    .B(_03329_),
    .Y(_12208_));
 sky130_fd_sc_hd__xnor2_2 _15033_ (.A(_03881_),
    .B(_04082_),
    .Y(_04445_));
 sky130_fd_sc_hd__xnor2_4 _15034_ (.A(_03505_),
    .B(_04445_),
    .Y(_12207_));
 sky130_fd_sc_hd__mux4_1 _15035_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net560),
    .S1(net570),
    .X(_04446_));
 sky130_fd_sc_hd__mux4_1 _15036_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net560),
    .S1(net570),
    .X(_04447_));
 sky130_fd_sc_hd__mux4_1 _15037_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net560),
    .S1(net570),
    .X(_04448_));
 sky130_fd_sc_hd__mux4_1 _15038_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net560),
    .S1(net570),
    .X(_04449_));
 sky130_fd_sc_hd__mux4_4 _15039_ (.A0(_04446_),
    .A1(_04447_),
    .A2(_04448_),
    .A3(_04449_),
    .S0(net557),
    .S1(net555),
    .X(_04450_));
 sky130_fd_sc_hd__mux4_1 _15040_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net565),
    .S1(net571),
    .X(_04451_));
 sky130_fd_sc_hd__mux4_1 _15041_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net565),
    .S1(net571),
    .X(_04452_));
 sky130_fd_sc_hd__mux4_1 _15042_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net565),
    .S1(net571),
    .X(_04453_));
 sky130_fd_sc_hd__mux4_1 _15043_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net565),
    .S1(net571),
    .X(_04454_));
 sky130_fd_sc_hd__mux4_1 _15044_ (.A0(_04451_),
    .A1(_04452_),
    .A2(_04453_),
    .A3(_04454_),
    .S0(net558),
    .S1(net556),
    .X(_04455_));
 sky130_fd_sc_hd__mux2i_4 _15045_ (.A0(_04450_),
    .A1(_04455_),
    .S(net554),
    .Y(_12206_));
 sky130_fd_sc_hd__mux4_1 _15046_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net637),
    .S1(net643),
    .X(_04456_));
 sky130_fd_sc_hd__mux4_1 _15047_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net637),
    .S1(net643),
    .X(_04457_));
 sky130_fd_sc_hd__mux4_1 _15048_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net637),
    .S1(net643),
    .X(_04458_));
 sky130_fd_sc_hd__mux4_1 _15049_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net637),
    .S1(net643),
    .X(_04459_));
 sky130_fd_sc_hd__mux4_4 _15050_ (.A0(_04456_),
    .A1(_04457_),
    .A2(_04458_),
    .A3(_04459_),
    .S0(net633),
    .S1(net632),
    .X(_04460_));
 sky130_fd_sc_hd__mux4_1 _15051_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net638),
    .S1(net643),
    .X(_04461_));
 sky130_fd_sc_hd__mux4_1 _15052_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net638),
    .S1(net643),
    .X(_04462_));
 sky130_fd_sc_hd__mux4_1 _15053_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net638),
    .S1(net643),
    .X(_04463_));
 sky130_fd_sc_hd__mux4_1 _15054_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net638),
    .S1(net643),
    .X(_04464_));
 sky130_fd_sc_hd__mux4_1 _15055_ (.A0(_04461_),
    .A1(_04462_),
    .A2(_04463_),
    .A3(_04464_),
    .S0(net633),
    .S1(net632),
    .X(_04465_));
 sky130_fd_sc_hd__mux2i_4 _15056_ (.A0(_04460_),
    .A1(_04465_),
    .S(net629),
    .Y(_12211_));
 sky130_fd_sc_hd__xnor2_1 _15057_ (.A(_03248_),
    .B(_03422_),
    .Y(_12216_));
 sky130_fd_sc_hd__xnor2_2 _15058_ (.A(_03927_),
    .B(_04128_),
    .Y(_04466_));
 sky130_fd_sc_hd__xnor2_4 _15059_ (.A(_03585_),
    .B(_04466_),
    .Y(_12215_));
 sky130_fd_sc_hd__mux4_1 _15060_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net564),
    .S1(net569),
    .X(_04467_));
 sky130_fd_sc_hd__mux4_1 _15061_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net564),
    .S1(net569),
    .X(_04468_));
 sky130_fd_sc_hd__mux4_1 _15062_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net564),
    .S1(net569),
    .X(_04469_));
 sky130_fd_sc_hd__mux4_1 _15063_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net564),
    .S1(net569),
    .X(_04470_));
 sky130_fd_sc_hd__mux4_4 _15064_ (.A0(_04467_),
    .A1(_04468_),
    .A2(_04469_),
    .A3(_04470_),
    .S0(net558),
    .S1(net556),
    .X(_04471_));
 sky130_fd_sc_hd__mux4_1 _15065_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net564),
    .S1(net571),
    .X(_04472_));
 sky130_fd_sc_hd__mux4_1 _15066_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net564),
    .S1(net571),
    .X(_04473_));
 sky130_fd_sc_hd__mux4_1 _15067_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net564),
    .S1(net571),
    .X(_04474_));
 sky130_fd_sc_hd__mux4_1 _15068_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net564),
    .S1(net571),
    .X(_04475_));
 sky130_fd_sc_hd__mux4_1 _15069_ (.A0(_04472_),
    .A1(_04473_),
    .A2(_04474_),
    .A3(_04475_),
    .S0(net558),
    .S1(net556),
    .X(_04476_));
 sky130_fd_sc_hd__mux2i_4 _15070_ (.A0(_04471_),
    .A1(_04476_),
    .S(net554),
    .Y(_12214_));
 sky130_fd_sc_hd__mux4_1 _15071_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net637),
    .S1(net646),
    .X(_04477_));
 sky130_fd_sc_hd__mux4_1 _15072_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net637),
    .S1(net646),
    .X(_04478_));
 sky130_fd_sc_hd__mux4_1 _15073_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net637),
    .S1(net646),
    .X(_04479_));
 sky130_fd_sc_hd__mux4_1 _15074_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net637),
    .S1(net646),
    .X(_04480_));
 sky130_fd_sc_hd__mux4_4 _15075_ (.A0(_04477_),
    .A1(_04478_),
    .A2(_04479_),
    .A3(_04480_),
    .S0(net633),
    .S1(net632),
    .X(_04481_));
 sky130_fd_sc_hd__mux4_1 _15076_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net638),
    .S1(net643),
    .X(_04482_));
 sky130_fd_sc_hd__mux4_1 _15077_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net638),
    .S1(net643),
    .X(_04483_));
 sky130_fd_sc_hd__mux4_1 _15078_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net638),
    .S1(net643),
    .X(_04484_));
 sky130_fd_sc_hd__mux4_1 _15079_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net638),
    .S1(net643),
    .X(_04485_));
 sky130_fd_sc_hd__mux4_1 _15080_ (.A0(_04482_),
    .A1(_04483_),
    .A2(_04484_),
    .A3(_04485_),
    .S0(net633),
    .S1(net631),
    .X(_04486_));
 sky130_fd_sc_hd__mux2i_4 _15081_ (.A0(_04481_),
    .A1(_04486_),
    .S(net629),
    .Y(_12219_));
 sky130_fd_sc_hd__xnor2_1 _15082_ (.A(_03329_),
    .B(_03481_),
    .Y(_12224_));
 sky130_fd_sc_hd__xnor2_2 _15083_ (.A(_03643_),
    .B(_03987_),
    .Y(_04487_));
 sky130_fd_sc_hd__xnor2_4 _15084_ (.A(_02995_),
    .B(_04487_),
    .Y(_12223_));
 sky130_fd_sc_hd__mux4_1 _15085_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04488_));
 sky130_fd_sc_hd__mux4_1 _15086_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04489_));
 sky130_fd_sc_hd__mux4_1 _15087_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04490_));
 sky130_fd_sc_hd__mux4_1 _15088_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04491_));
 sky130_fd_sc_hd__mux4_4 _15089_ (.A0(_04488_),
    .A1(_04489_),
    .A2(_04490_),
    .A3(_04491_),
    .S0(net558),
    .S1(net556),
    .X(_04492_));
 sky130_fd_sc_hd__mux4_1 _15090_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04493_));
 sky130_fd_sc_hd__mux4_1 _15091_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04494_));
 sky130_fd_sc_hd__mux4_1 _15092_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04495_));
 sky130_fd_sc_hd__mux4_1 _15093_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net564),
    .S1(net569),
    .X(_04496_));
 sky130_fd_sc_hd__mux4_1 _15094_ (.A0(_04493_),
    .A1(_04494_),
    .A2(_04495_),
    .A3(_04496_),
    .S0(net558),
    .S1(net556),
    .X(_04497_));
 sky130_fd_sc_hd__mux2i_4 _15095_ (.A0(_04492_),
    .A1(_04497_),
    .S(net554),
    .Y(_12222_));
 sky130_fd_sc_hd__mux4_1 _15096_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net638),
    .S1(net643),
    .X(_04498_));
 sky130_fd_sc_hd__mux4_1 _15097_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net638),
    .S1(net643),
    .X(_04499_));
 sky130_fd_sc_hd__mux4_1 _15098_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net638),
    .S1(net643),
    .X(_04500_));
 sky130_fd_sc_hd__mux4_1 _15099_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net638),
    .S1(net643),
    .X(_04501_));
 sky130_fd_sc_hd__mux4_4 _15100_ (.A0(_04498_),
    .A1(_04499_),
    .A2(_04500_),
    .A3(_04501_),
    .S0(net633),
    .S1(net632),
    .X(_04502_));
 sky130_fd_sc_hd__mux4_1 _15101_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net635),
    .S1(net644),
    .X(_04503_));
 sky130_fd_sc_hd__mux4_1 _15102_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net635),
    .S1(net644),
    .X(_04504_));
 sky130_fd_sc_hd__mux4_1 _15103_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net635),
    .S1(net644),
    .X(_04505_));
 sky130_fd_sc_hd__mux4_1 _15104_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net635),
    .S1(net644),
    .X(_04506_));
 sky130_fd_sc_hd__mux4_1 _15105_ (.A0(_04503_),
    .A1(_04504_),
    .A2(_04505_),
    .A3(_04506_),
    .S0(net634),
    .S1(net632),
    .X(_04507_));
 sky130_fd_sc_hd__mux2i_4 _15106_ (.A0(_04502_),
    .A1(_04507_),
    .S(net629),
    .Y(_12227_));
 sky130_fd_sc_hd__xnor2_1 _15107_ (.A(_03422_),
    .B(_03551_),
    .Y(_12232_));
 sky130_fd_sc_hd__xnor2_4 _15108_ (.A(_03147_),
    .B(_03691_),
    .Y(_12231_));
 sky130_fd_sc_hd__mux4_1 _15109_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net561),
    .S1(net572),
    .X(_04508_));
 sky130_fd_sc_hd__mux4_1 _15110_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net561),
    .S1(net572),
    .X(_04509_));
 sky130_fd_sc_hd__mux4_1 _15111_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net561),
    .S1(net572),
    .X(_04510_));
 sky130_fd_sc_hd__mux4_1 _15112_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net561),
    .S1(net572),
    .X(_04511_));
 sky130_fd_sc_hd__mux4_4 _15113_ (.A0(_04508_),
    .A1(_04509_),
    .A2(_04510_),
    .A3(_04511_),
    .S0(net559),
    .S1(net555),
    .X(_04512_));
 sky130_fd_sc_hd__mux4_1 _15114_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net566),
    .S1(net571),
    .X(_04513_));
 sky130_fd_sc_hd__mux4_1 _15115_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net566),
    .S1(net571),
    .X(_04514_));
 sky130_fd_sc_hd__mux4_1 _15116_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net566),
    .S1(net571),
    .X(_04515_));
 sky130_fd_sc_hd__mux4_1 _15117_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net566),
    .S1(net571),
    .X(_04516_));
 sky130_fd_sc_hd__mux4_1 _15118_ (.A0(_04513_),
    .A1(_04514_),
    .A2(_04515_),
    .A3(_04516_),
    .S0(net557),
    .S1(net555),
    .X(_04517_));
 sky130_fd_sc_hd__mux2i_4 _15119_ (.A0(_04512_),
    .A1(_04517_),
    .S(net553),
    .Y(_12230_));
 sky130_fd_sc_hd__mux4_1 _15120_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net640),
    .S1(net645),
    .X(_04518_));
 sky130_fd_sc_hd__mux4_1 _15121_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net640),
    .S1(net645),
    .X(_04519_));
 sky130_fd_sc_hd__mux4_1 _15122_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net640),
    .S1(net645),
    .X(_04520_));
 sky130_fd_sc_hd__mux4_1 _15123_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net640),
    .S1(net645),
    .X(_04521_));
 sky130_fd_sc_hd__mux4_4 _15124_ (.A0(_04518_),
    .A1(_04519_),
    .A2(_04520_),
    .A3(_04521_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04522_));
 sky130_fd_sc_hd__mux4_1 _15125_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net640),
    .S1(net645),
    .X(_04523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1411 ();
 sky130_fd_sc_hd__mux4_1 _15127_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net635),
    .S1(net644),
    .X(_04525_));
 sky130_fd_sc_hd__mux4_1 _15128_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net635),
    .S1(net644),
    .X(_04526_));
 sky130_fd_sc_hd__mux4_1 _15129_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net635),
    .S1(net644),
    .X(_04527_));
 sky130_fd_sc_hd__mux4_1 _15130_ (.A0(_04523_),
    .A1(_04525_),
    .A2(_04526_),
    .A3(_04527_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_04528_));
 sky130_fd_sc_hd__mux2i_4 _15131_ (.A0(_04522_),
    .A1(_04528_),
    .S(net630),
    .Y(_12235_));
 sky130_fd_sc_hd__xnor2_1 _15132_ (.A(_02959_),
    .B(_03481_),
    .Y(_12240_));
 sky130_fd_sc_hd__xnor2_2 _15133_ (.A(_03271_),
    .B(_03762_),
    .Y(_12239_));
 sky130_fd_sc_hd__mux4_1 _15134_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04529_));
 sky130_fd_sc_hd__mux4_1 _15135_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04530_));
 sky130_fd_sc_hd__mux4_1 _15136_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04531_));
 sky130_fd_sc_hd__mux4_1 _15137_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_04532_));
 sky130_fd_sc_hd__mux4_4 _15138_ (.A0(_04529_),
    .A1(_04530_),
    .A2(_04531_),
    .A3(_04532_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_04533_));
 sky130_fd_sc_hd__mux4_1 _15139_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net562),
    .S1(net567),
    .X(_04534_));
 sky130_fd_sc_hd__mux4_1 _15140_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net562),
    .S1(net567),
    .X(_04535_));
 sky130_fd_sc_hd__mux4_1 _15141_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net562),
    .S1(net567),
    .X(_04536_));
 sky130_fd_sc_hd__mux4_1 _15142_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net562),
    .S1(net567),
    .X(_04537_));
 sky130_fd_sc_hd__mux4_1 _15143_ (.A0(_04534_),
    .A1(_04535_),
    .A2(_04536_),
    .A3(_04537_),
    .S0(net559),
    .S1(\count7_2[4] ),
    .X(_04538_));
 sky130_fd_sc_hd__mux2i_4 _15144_ (.A0(_04533_),
    .A1(_04538_),
    .S(net553),
    .Y(_12238_));
 sky130_fd_sc_hd__mux4_1 _15145_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04539_));
 sky130_fd_sc_hd__mux4_1 _15146_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04540_));
 sky130_fd_sc_hd__mux4_1 _15147_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04541_));
 sky130_fd_sc_hd__mux4_1 _15148_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04542_));
 sky130_fd_sc_hd__mux4_2 _15149_ (.A0(_04539_),
    .A1(_04540_),
    .A2(_04541_),
    .A3(_04542_),
    .S0(net634),
    .S1(net632),
    .X(_04543_));
 sky130_fd_sc_hd__mux4_1 _15150_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04544_));
 sky130_fd_sc_hd__mux4_1 _15151_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04545_));
 sky130_fd_sc_hd__mux4_1 _15152_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04546_));
 sky130_fd_sc_hd__mux4_1 _15153_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net635),
    .S1(net644),
    .X(_04547_));
 sky130_fd_sc_hd__mux4_1 _15154_ (.A0(_04544_),
    .A1(_04545_),
    .A2(_04546_),
    .A3(_04547_),
    .S0(net634),
    .S1(net632),
    .X(_04548_));
 sky130_fd_sc_hd__mux2i_4 _15155_ (.A0(_04543_),
    .A1(_04548_),
    .S(net630),
    .Y(_12243_));
 sky130_fd_sc_hd__a21o_1 _15156_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_13090_),
    .B1(\hash.CA2.b_dash[0] ),
    .X(_04549_));
 sky130_fd_sc_hd__o21ai_0 _15157_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_13090_),
    .B1(_04549_),
    .Y(_12248_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1408 ();
 sky130_fd_sc_hd__xnor2_4 _15161_ (.A(\hash.CA2.S1.X[6] ),
    .B(net1106),
    .Y(_04553_));
 sky130_fd_sc_hd__xnor2_2 _15162_ (.A(\hash.CA2.S1.X[11] ),
    .B(_04553_),
    .Y(_13398_));
 sky130_fd_sc_hd__o21a_1 _15163_ (.A1(_13130_),
    .A2(_13129_),
    .B1(_13128_),
    .X(_04554_));
 sky130_fd_sc_hd__nor2_1 _15164_ (.A(_13127_),
    .B(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1406 ();
 sky130_fd_sc_hd__inv_1 _15167_ (.A(_13122_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21oi_1 _15168_ (.A1(_13118_),
    .A2(_13119_),
    .B1(_13117_),
    .Y(_04559_));
 sky130_fd_sc_hd__o21bai_1 _15169_ (.A1(_04558_),
    .A2(_04559_),
    .B1_N(_13121_),
    .Y(_04560_));
 sky130_fd_sc_hd__a21o_1 _15170_ (.A1(_13124_),
    .A2(_04560_),
    .B1(_13123_),
    .X(_04561_));
 sky130_fd_sc_hd__a21o_1 _15171_ (.A1(_13126_),
    .A2(_04561_),
    .B1(_13125_),
    .X(_04562_));
 sky130_fd_sc_hd__a2111oi_4 _15172_ (.A1(_13132_),
    .A2(_04562_),
    .B1(_13131_),
    .C1(_13129_),
    .D1(_13127_),
    .Y(_04563_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1405 ();
 sky130_fd_sc_hd__and2_2 _15174_ (.A(_13106_),
    .B(_13110_),
    .X(_04565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1404 ();
 sky130_fd_sc_hd__a22oi_4 _15176_ (.A1(_13110_),
    .A2(_13105_),
    .B1(_13107_),
    .B2(_04565_),
    .Y(_04567_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1402 ();
 sky130_fd_sc_hd__o21ai_0 _15179_ (.A1(_13098_),
    .A2(_13097_),
    .B1(_13096_),
    .Y(_04570_));
 sky130_fd_sc_hd__nand2b_2 _15180_ (.A_N(_13095_),
    .B(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21o_1 _15181_ (.A1(_12252_),
    .A2(_13092_),
    .B1(_13091_),
    .X(_04572_));
 sky130_fd_sc_hd__a21oi_4 _15182_ (.A1(_13104_),
    .A2(_04572_),
    .B1(_13103_),
    .Y(_04573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1401 ();
 sky130_fd_sc_hd__nand2_1 _15184_ (.A(_13100_),
    .B(_13102_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21oi_2 _15185_ (.A1(_13100_),
    .A2(_13101_),
    .B1(_13099_),
    .Y(_04576_));
 sky130_fd_sc_hd__nor2_1 _15186_ (.A(_13095_),
    .B(_13097_),
    .Y(_04577_));
 sky130_fd_sc_hd__o211ai_4 _15187_ (.A1(_04575_),
    .A2(_04573_),
    .B1(_04576_),
    .C1(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand4_4 _15188_ (.A(_04571_),
    .B(_04578_),
    .C(_13108_),
    .D(_04565_),
    .Y(_04579_));
 sky130_fd_sc_hd__nor3_1 _15189_ (.A(_13109_),
    .B(_13111_),
    .C(_13115_),
    .Y(_04580_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1400 ();
 sky130_fd_sc_hd__nor2_1 _15191_ (.A(_13112_),
    .B(_13111_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2b_2 _15192_ (.A(_04582_),
    .B_N(_13116_),
    .Y(_04583_));
 sky130_fd_sc_hd__o21ai_4 _15193_ (.A1(_13115_),
    .A2(_04583_),
    .B1(_13114_),
    .Y(_04584_));
 sky130_fd_sc_hd__a31oi_4 _15194_ (.A1(_04567_),
    .A2(_04579_),
    .A3(_04580_),
    .B1(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__nand4_1 _15195_ (.A(_13126_),
    .B(_13128_),
    .C(_13130_),
    .D(_13132_),
    .Y(_04586_));
 sky130_fd_sc_hd__nand4_4 _15196_ (.A(_13118_),
    .B(_13120_),
    .C(_13122_),
    .D(_13124_),
    .Y(_04587_));
 sky130_fd_sc_hd__nor2_2 _15197_ (.A(_04586_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__o21ai_2 _15198_ (.A1(_13113_),
    .A2(_04585_),
    .B1(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__o21ai_4 _15199_ (.A1(_04555_),
    .A2(_04563_),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__xor2_4 _15200_ (.A(_04590_),
    .B(_13134_),
    .X(_04591_));
 sky130_fd_sc_hd__xor2_4 _15201_ (.A(_13092_),
    .B(_12252_),
    .X(_04592_));
 sky130_fd_sc_hd__a21oi_2 _15202_ (.A1(_13098_),
    .A2(_13099_),
    .B1(_13097_),
    .Y(_04593_));
 sky130_fd_sc_hd__nand2_1 _15203_ (.A(_13096_),
    .B(_13108_),
    .Y(_04594_));
 sky130_fd_sc_hd__a21oi_1 _15204_ (.A1(_13108_),
    .A2(_13095_),
    .B1(_13107_),
    .Y(_04595_));
 sky130_fd_sc_hd__o21ai_2 _15205_ (.A1(_04593_),
    .A2(_04594_),
    .B1(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__a21o_1 _15206_ (.A1(_13110_),
    .A2(_13105_),
    .B1(_13109_),
    .X(_04597_));
 sky130_fd_sc_hd__a211o_1 _15207_ (.A1(_13116_),
    .A2(_13111_),
    .B1(_13115_),
    .C1(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__a21oi_2 _15208_ (.A1(_04565_),
    .A2(_04596_),
    .B1(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__a211oi_2 _15209_ (.A1(_12251_),
    .A2(_13094_),
    .B1(_13091_),
    .C1(_13093_),
    .Y(_04600_));
 sky130_fd_sc_hd__o21ai_1 _15210_ (.A1(_13092_),
    .A2(_13091_),
    .B1(_13104_),
    .Y(_04601_));
 sky130_fd_sc_hd__o21bai_4 _15211_ (.A1(_04600_),
    .A2(_04601_),
    .B1_N(_13103_),
    .Y(_04602_));
 sky130_fd_sc_hd__nand2_1 _15212_ (.A(_13106_),
    .B(_13110_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand3_1 _15213_ (.A(_13100_),
    .B(_13102_),
    .C(_13098_),
    .Y(_04604_));
 sky130_fd_sc_hd__nor3_1 _15214_ (.A(_04603_),
    .B(_04594_),
    .C(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__nand3_1 _15215_ (.A(_13100_),
    .B(_13098_),
    .C(_13101_),
    .Y(_04606_));
 sky130_fd_sc_hd__nor3_1 _15216_ (.A(_04603_),
    .B(_04594_),
    .C(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__a21oi_4 _15217_ (.A1(_04602_),
    .A2(_04605_),
    .B1(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__nand2_2 _15218_ (.A(_04599_),
    .B(_04608_),
    .Y(_04609_));
 sky130_fd_sc_hd__o21a_2 _15219_ (.A1(_13115_),
    .A2(_04583_),
    .B1(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__xnor2_4 _15220_ (.A(_13114_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__xnor2_2 _15221_ (.A(_04592_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__xnor2_4 _15222_ (.A(net1120),
    .B(_04612_),
    .Y(_12246_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1398 ();
 sky130_fd_sc_hd__nor2_1 _15225_ (.A(net520),
    .B(_13403_),
    .Y(_00658_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1397 ();
 sky130_fd_sc_hd__a21o_1 _15227_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_12253_),
    .B1(\hash.CA2.b_dash[1] ),
    .X(_04616_));
 sky130_fd_sc_hd__o21ai_1 _15228_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_12253_),
    .B1(_04616_),
    .Y(_12261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1394 ();
 sky130_fd_sc_hd__xnor2_4 _15232_ (.A(\hash.CA2.S1.X[12] ),
    .B(\hash.CA2.S1.X[26] ),
    .Y(_04620_));
 sky130_fd_sc_hd__xnor2_2 _15233_ (.A(\hash.CA2.S1.X[7] ),
    .B(_04620_),
    .Y(_13405_));
 sky130_fd_sc_hd__inv_1 _15234_ (.A(_13405_),
    .Y(_12256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1393 ();
 sky130_fd_sc_hd__mux2_1 _15236_ (.A0(\hash.CA2.f_dash[1] ),
    .A1(\hash.CA2.e_dash[1] ),
    .S(\hash.CA2.S1.X[1] ),
    .X(_13404_));
 sky130_fd_sc_hd__inv_1 _15237_ (.A(_13404_),
    .Y(_12255_));
 sky130_fd_sc_hd__nor4_2 _15238_ (.A(_13109_),
    .B(_13111_),
    .C(_13113_),
    .D(_13115_),
    .Y(_04622_));
 sky130_fd_sc_hd__o21a_2 _15239_ (.A1(_13115_),
    .A2(_04583_),
    .B1(_13114_),
    .X(_04623_));
 sky130_fd_sc_hd__o21ai_1 _15240_ (.A1(_13113_),
    .A2(_04623_),
    .B1(_13120_),
    .Y(_04624_));
 sky130_fd_sc_hd__a31oi_4 _15241_ (.A1(_04567_),
    .A2(_04579_),
    .A3(_04622_),
    .B1(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__nor3_2 _15242_ (.A(_13120_),
    .B(_13113_),
    .C(_04585_),
    .Y(_04626_));
 sky130_fd_sc_hd__nor2_8 _15243_ (.A(_04625_),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1392 ();
 sky130_fd_sc_hd__a21oi_4 _15245_ (.A1(_04599_),
    .A2(_04608_),
    .B1(_04584_),
    .Y(_04629_));
 sky130_fd_sc_hd__inv_1 _15246_ (.A(_13118_),
    .Y(_04630_));
 sky130_fd_sc_hd__a21oi_1 _15247_ (.A1(_13120_),
    .A2(_13113_),
    .B1(_13119_),
    .Y(_04631_));
 sky130_fd_sc_hd__inv_1 _15248_ (.A(_13117_),
    .Y(_04632_));
 sky130_fd_sc_hd__o21ai_1 _15249_ (.A1(_04630_),
    .A2(_04631_),
    .B1(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__a21o_1 _15250_ (.A1(_13124_),
    .A2(_13121_),
    .B1(_13123_),
    .X(_04634_));
 sky130_fd_sc_hd__a31oi_4 _15251_ (.A1(_13122_),
    .A2(_13124_),
    .A3(_04633_),
    .B1(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__inv_1 _15252_ (.A(_13130_),
    .Y(_04636_));
 sky130_fd_sc_hd__a21oi_1 _15253_ (.A1(_13132_),
    .A2(_13125_),
    .B1(_13131_),
    .Y(_04637_));
 sky130_fd_sc_hd__o21bai_1 _15254_ (.A1(_04636_),
    .A2(_04637_),
    .B1_N(_13129_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand2_1 _15255_ (.A(_13128_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__o21ai_2 _15256_ (.A1(_04586_),
    .A2(_04635_),
    .B1(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__a211o_1 _15257_ (.A1(_04588_),
    .A2(_04629_),
    .B1(_04640_),
    .C1(_13127_),
    .X(_04641_));
 sky130_fd_sc_hd__a21o_1 _15258_ (.A1(_13134_),
    .A2(_04641_),
    .B1(_13133_),
    .X(_04642_));
 sky130_fd_sc_hd__xor2_4 _15259_ (.A(_13138_),
    .B(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__a21o_1 _15260_ (.A1(_12251_),
    .A2(_13094_),
    .B1(_13093_),
    .X(_04644_));
 sky130_fd_sc_hd__a21oi_2 _15261_ (.A1(_13092_),
    .A2(_04644_),
    .B1(_13091_),
    .Y(_04645_));
 sky130_fd_sc_hd__xor2_4 _15262_ (.A(_13104_),
    .B(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__xnor2_2 _15263_ (.A(_04643_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__xnor2_4 _15264_ (.A(_04627_),
    .B(_04647_),
    .Y(_12259_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1391 ();
 sky130_fd_sc_hd__or2_0 _15266_ (.A(net520),
    .B(_13409_),
    .X(\hash.CA1.S0.X[1] ));
 sky130_fd_sc_hd__inv_1 _15267_ (.A(\hash.CA1.S0.X[1] ),
    .Y(_13711_));
 sky130_fd_sc_hd__maj3_1 _15268_ (.A(\hash.CA2.b_dash[2] ),
    .B(\hash.CA2.a_dash[2] ),
    .C(_04592_),
    .X(_04649_));
 sky130_fd_sc_hd__inv_1 _15269_ (.A(_04649_),
    .Y(_12270_));
 sky130_fd_sc_hd__xnor2_1 _15270_ (.A(_12257_),
    .B(_13413_),
    .Y(_13414_));
 sky130_fd_sc_hd__inv_1 _15271_ (.A(_13414_),
    .Y(_12269_));
 sky130_fd_sc_hd__a21o_1 _15272_ (.A1(_13138_),
    .A2(_13133_),
    .B1(_13137_),
    .X(_04650_));
 sky130_fd_sc_hd__a31oi_4 _15273_ (.A1(_13134_),
    .A2(_13138_),
    .A3(_04590_),
    .B1(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__xnor2_4 _15274_ (.A(_04651_),
    .B(_13136_),
    .Y(_04652_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1390 ();
 sky130_fd_sc_hd__xnor2_4 _15276_ (.A(_13102_),
    .B(net1126),
    .Y(_04654_));
 sky130_fd_sc_hd__inv_1 _15277_ (.A(_13119_),
    .Y(_04655_));
 sky130_fd_sc_hd__o21ai_2 _15278_ (.A1(_13113_),
    .A2(_04629_),
    .B1(_13120_),
    .Y(_04656_));
 sky130_fd_sc_hd__a21oi_4 _15279_ (.A1(_04655_),
    .A2(_04656_),
    .B1(_04630_),
    .Y(_04657_));
 sky130_fd_sc_hd__and3_2 _15280_ (.A(_04630_),
    .B(_04655_),
    .C(_04656_),
    .X(_04658_));
 sky130_fd_sc_hd__nor2_8 _15281_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__xor2_2 _15282_ (.A(_04654_),
    .B(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__xnor2_4 _15283_ (.A(net1135),
    .B(_04660_),
    .Y(_12268_));
 sky130_fd_sc_hd__inv_1 _15284_ (.A(\hash.CA2.b_dash[3] ),
    .Y(_04661_));
 sky130_fd_sc_hd__inv_1 _15285_ (.A(\hash.CA2.a_dash[3] ),
    .Y(_04662_));
 sky130_fd_sc_hd__maj3_1 _15286_ (.A(_04661_),
    .B(_04662_),
    .C(_04646_),
    .X(_12284_));
 sky130_fd_sc_hd__a21o_1 _15287_ (.A1(_13399_),
    .A2(_13407_),
    .B1(_13406_),
    .X(_04663_));
 sky130_fd_sc_hd__a21oi_1 _15288_ (.A1(_13413_),
    .A2(_04663_),
    .B1(_13412_),
    .Y(_04664_));
 sky130_fd_sc_hd__xnor2_1 _15289_ (.A(_13420_),
    .B(_04664_),
    .Y(_13421_));
 sky130_fd_sc_hd__inv_1 _15290_ (.A(_13421_),
    .Y(_12283_));
 sky130_fd_sc_hd__a21o_1 _15291_ (.A1(_13138_),
    .A2(_04642_),
    .B1(_13137_),
    .X(_04665_));
 sky130_fd_sc_hd__a21oi_2 _15292_ (.A1(_13136_),
    .A2(_04665_),
    .B1(_13135_),
    .Y(_04666_));
 sky130_fd_sc_hd__xnor2_4 _15293_ (.A(_04666_),
    .B(_13140_),
    .Y(_04667_));
 sky130_fd_sc_hd__nor4_1 _15294_ (.A(_04558_),
    .B(_13117_),
    .C(_13119_),
    .D(_04625_),
    .Y(_04668_));
 sky130_fd_sc_hd__nor3_1 _15295_ (.A(_13118_),
    .B(_04558_),
    .C(_13117_),
    .Y(_04669_));
 sky130_fd_sc_hd__a31oi_1 _15296_ (.A1(_13118_),
    .A2(_04558_),
    .A3(_13119_),
    .B1(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__o21ai_1 _15297_ (.A1(_13122_),
    .A2(_04632_),
    .B1(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__a311oi_4 _15298_ (.A1(_13118_),
    .A2(_04558_),
    .A3(_04625_),
    .B1(_04671_),
    .C1(_04668_),
    .Y(_04672_));
 sky130_fd_sc_hd__a21oi_4 _15299_ (.A1(_13102_),
    .A2(_04602_),
    .B1(_13101_),
    .Y(_04673_));
 sky130_fd_sc_hd__xnor2_4 _15300_ (.A(_13100_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__xnor2_2 _15301_ (.A(_04672_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__xnor2_4 _15302_ (.A(net1166),
    .B(_04675_),
    .Y(_12282_));
 sky130_fd_sc_hd__nand2_1 _15303_ (.A(\hash.CA2.a_dash[4] ),
    .B(_04654_),
    .Y(_04676_));
 sky130_fd_sc_hd__o21ai_0 _15304_ (.A1(\hash.CA2.a_dash[4] ),
    .A2(_04654_),
    .B1(\hash.CA2.b_dash[4] ),
    .Y(_04677_));
 sky130_fd_sc_hd__and2_0 _15305_ (.A(_04676_),
    .B(_04677_),
    .X(_12293_));
 sky130_fd_sc_hd__inv_1 _15306_ (.A(_13419_),
    .Y(_04678_));
 sky130_fd_sc_hd__nor2b_2 _15307_ (.A(_12257_),
    .B_N(_13413_),
    .Y(_04679_));
 sky130_fd_sc_hd__o21ai_2 _15308_ (.A1(_13412_),
    .A2(_04679_),
    .B1(_13420_),
    .Y(_04680_));
 sky130_fd_sc_hd__a21boi_2 _15309_ (.A1(_04680_),
    .A2(_04678_),
    .B1_N(_13427_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand2_1 _15310_ (.A(_04678_),
    .B(_04680_),
    .Y(_04682_));
 sky130_fd_sc_hd__nor2_1 _15311_ (.A(_13427_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__nor2_1 _15312_ (.A(net1029),
    .B(_04683_),
    .Y(_13428_));
 sky130_fd_sc_hd__inv_1 _15313_ (.A(_13428_),
    .Y(_12292_));
 sky130_fd_sc_hd__and3_1 _15314_ (.A(_13136_),
    .B(_13138_),
    .C(_13140_),
    .X(_04684_));
 sky130_fd_sc_hd__and3_1 _15315_ (.A(_13134_),
    .B(_13144_),
    .C(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__o211ai_4 _15316_ (.A1(_13113_),
    .A2(_04585_),
    .B1(_04588_),
    .C1(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand3_1 _15317_ (.A(_13134_),
    .B(_13144_),
    .C(_04684_),
    .Y(_04687_));
 sky130_fd_sc_hd__a21o_1 _15318_ (.A1(_13136_),
    .A2(_04650_),
    .B1(_13135_),
    .X(_04688_));
 sky130_fd_sc_hd__a21o_1 _15319_ (.A1(_13140_),
    .A2(_04688_),
    .B1(_13139_),
    .X(_04689_));
 sky130_fd_sc_hd__nand2_1 _15320_ (.A(_13144_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__o31a_2 _15321_ (.A1(_04555_),
    .A2(_04563_),
    .A3(_04687_),
    .B1(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__nand2_2 _15322_ (.A(_04686_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__a311oi_4 _15323_ (.A1(_13134_),
    .A2(_04590_),
    .A3(_04684_),
    .B1(_04689_),
    .C1(_13144_),
    .Y(_04693_));
 sky130_fd_sc_hd__nor2_8 _15324_ (.A(_04693_),
    .B(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__nor3_1 _15325_ (.A(_13117_),
    .B(_13119_),
    .C(_13121_),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_1 _15326_ (.A(_04630_),
    .B(_04632_),
    .Y(_04696_));
 sky130_fd_sc_hd__a21oi_1 _15327_ (.A1(_13122_),
    .A2(_04696_),
    .B1(_13121_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21oi_2 _15328_ (.A1(_04656_),
    .A2(_04695_),
    .B1(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__xor2_4 _15329_ (.A(_13124_),
    .B(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__o21ai_2 _15330_ (.A1(net1158),
    .A2(_04575_),
    .B1(_04576_),
    .Y(_04700_));
 sky130_fd_sc_hd__xor2_4 _15331_ (.A(_13098_),
    .B(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__xor2_2 _15332_ (.A(_04699_),
    .B(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__xnor2_4 _15333_ (.A(_04694_),
    .B(_04702_),
    .Y(_12291_));
 sky130_fd_sc_hd__maj3_1 _15334_ (.A(\hash.CA2.b_dash[5] ),
    .B(\hash.CA2.a_dash[5] ),
    .C(_04674_),
    .X(_04703_));
 sky130_fd_sc_hd__inv_1 _15335_ (.A(_04703_),
    .Y(_12302_));
 sky130_fd_sc_hd__a211oi_1 _15336_ (.A1(net1024),
    .A2(_13407_),
    .B1(_13406_),
    .C1(_13412_),
    .Y(_04704_));
 sky130_fd_sc_hd__o21ai_0 _15337_ (.A1(_13413_),
    .A2(_13412_),
    .B1(_13420_),
    .Y(_04705_));
 sky130_fd_sc_hd__o21ai_0 _15338_ (.A1(_04704_),
    .A2(_04705_),
    .B1(_04678_),
    .Y(_04706_));
 sky130_fd_sc_hd__a21oi_1 _15339_ (.A1(_13427_),
    .A2(_04706_),
    .B1(_13426_),
    .Y(_04707_));
 sky130_fd_sc_hd__xnor2_1 _15340_ (.A(_13434_),
    .B(_04707_),
    .Y(_13435_));
 sky130_fd_sc_hd__inv_1 _15341_ (.A(_13435_),
    .Y(_12301_));
 sky130_fd_sc_hd__a31oi_4 _15342_ (.A1(_04623_),
    .A2(_04588_),
    .A3(_04609_),
    .B1(_04640_),
    .Y(_04708_));
 sky130_fd_sc_hd__a21o_1 _15343_ (.A1(_13136_),
    .A2(_13137_),
    .B1(_13135_),
    .X(_04709_));
 sky130_fd_sc_hd__a21oi_2 _15344_ (.A1(_13140_),
    .A2(_04709_),
    .B1(_13139_),
    .Y(_04710_));
 sky130_fd_sc_hd__nor2_1 _15345_ (.A(_13127_),
    .B(_13133_),
    .Y(_04711_));
 sky130_fd_sc_hd__or2_0 _15346_ (.A(_13134_),
    .B(_13133_),
    .X(_04712_));
 sky130_fd_sc_hd__a21boi_2 _15347_ (.A1(_04684_),
    .A2(_04712_),
    .B1_N(_04710_),
    .Y(_04713_));
 sky130_fd_sc_hd__a31oi_1 _15348_ (.A1(_04708_),
    .A2(_04710_),
    .A3(_04711_),
    .B1(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__a21oi_2 _15349_ (.A1(_13144_),
    .A2(_04714_),
    .B1(_13143_),
    .Y(_04715_));
 sky130_fd_sc_hd__xnor2_4 _15350_ (.A(_13142_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand3_2 _15351_ (.A(_04567_),
    .B(_04579_),
    .C(_04622_),
    .Y(_04717_));
 sky130_fd_sc_hd__nor2_1 _15352_ (.A(_13113_),
    .B(_04623_),
    .Y(_04718_));
 sky130_fd_sc_hd__nor2_1 _15353_ (.A(_04587_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__a21oi_2 _15354_ (.A1(_04717_),
    .A2(_04719_),
    .B1(_04561_),
    .Y(_04720_));
 sky130_fd_sc_hd__xnor2_4 _15355_ (.A(_13126_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _15356_ (.A(_13100_),
    .B(_13098_),
    .Y(_04722_));
 sky130_fd_sc_hd__o21ai_2 _15357_ (.A1(_04722_),
    .A2(_04673_),
    .B1(_04593_),
    .Y(_04723_));
 sky130_fd_sc_hd__xor2_4 _15358_ (.A(_13096_),
    .B(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__xnor2_2 _15359_ (.A(_04721_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__xor2_4 _15360_ (.A(_04716_),
    .B(_04725_),
    .X(_12300_));
 sky130_fd_sc_hd__maj3_1 _15361_ (.A(\hash.CA2.b_dash[6] ),
    .B(\hash.CA2.a_dash[6] ),
    .C(_04701_),
    .X(_04726_));
 sky130_fd_sc_hd__inv_1 _15362_ (.A(_04726_),
    .Y(_12311_));
 sky130_fd_sc_hd__inv_1 _15363_ (.A(_13441_),
    .Y(_04727_));
 sky130_fd_sc_hd__inv_1 _15364_ (.A(_13433_),
    .Y(_04728_));
 sky130_fd_sc_hd__o21ai_2 _15365_ (.A1(_04681_),
    .A2(_13426_),
    .B1(_13434_),
    .Y(_04729_));
 sky130_fd_sc_hd__nand2_1 _15366_ (.A(_04728_),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__xnor2_1 _15367_ (.A(_04727_),
    .B(_04730_),
    .Y(_13442_));
 sky130_fd_sc_hd__inv_1 _15368_ (.A(_13442_),
    .Y(_12310_));
 sky130_fd_sc_hd__nor2_1 _15369_ (.A(_13141_),
    .B(_13143_),
    .Y(_04731_));
 sky130_fd_sc_hd__o21ai_1 _15370_ (.A1(_13142_),
    .A2(_13141_),
    .B1(_13146_),
    .Y(_04732_));
 sky130_fd_sc_hd__a31oi_4 _15371_ (.A1(_04691_),
    .A2(_04686_),
    .A3(_04731_),
    .B1(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__nand3b_1 _15372_ (.A_N(_13143_),
    .B(_04686_),
    .C(_04691_),
    .Y(_04734_));
 sky130_fd_sc_hd__a211oi_4 _15373_ (.A1(_13142_),
    .A2(_04734_),
    .B1(_13141_),
    .C1(_13146_),
    .Y(_04735_));
 sky130_fd_sc_hd__nor2_8 _15374_ (.A(net1137),
    .B(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__inv_1 _15375_ (.A(_04587_),
    .Y(_04737_));
 sky130_fd_sc_hd__a21bo_1 _15376_ (.A1(_04737_),
    .A2(_04629_),
    .B1_N(_04635_),
    .X(_04738_));
 sky130_fd_sc_hd__a21o_2 _15377_ (.A1(_13126_),
    .A2(_04738_),
    .B1(_13125_),
    .X(_04739_));
 sky130_fd_sc_hd__xnor2_4 _15378_ (.A(_13132_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand2_1 _15379_ (.A(_04571_),
    .B(_04578_),
    .Y(_04741_));
 sky130_fd_sc_hd__xnor2_4 _15380_ (.A(_13108_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__xnor2_2 _15381_ (.A(_04740_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__xnor2_4 _15382_ (.A(_04736_),
    .B(_04743_),
    .Y(_12309_));
 sky130_fd_sc_hd__maj3_1 _15383_ (.A(\hash.CA2.b_dash[7] ),
    .B(\hash.CA2.a_dash[7] ),
    .C(_04724_),
    .X(_04744_));
 sky130_fd_sc_hd__inv_1 _15384_ (.A(_04744_),
    .Y(_12320_));
 sky130_fd_sc_hd__o21ai_1 _15385_ (.A1(_13427_),
    .A2(_13426_),
    .B1(_13434_),
    .Y(_04745_));
 sky130_fd_sc_hd__nor3_1 _15386_ (.A(_13419_),
    .B(_13426_),
    .C(_13433_),
    .Y(_04746_));
 sky130_fd_sc_hd__o21a_1 _15387_ (.A1(_04704_),
    .A2(_04705_),
    .B1(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__a21oi_1 _15388_ (.A1(_04728_),
    .A2(_04745_),
    .B1(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__a21oi_1 _15389_ (.A1(_13441_),
    .A2(_04748_),
    .B1(_13440_),
    .Y(_04749_));
 sky130_fd_sc_hd__xnor2_1 _15390_ (.A(_13448_),
    .B(_04749_),
    .Y(_13449_));
 sky130_fd_sc_hd__inv_1 _15391_ (.A(_13449_),
    .Y(_12319_));
 sky130_fd_sc_hd__nand3_1 _15392_ (.A(_13142_),
    .B(_13144_),
    .C(_13146_),
    .Y(_04750_));
 sky130_fd_sc_hd__a311oi_4 _15393_ (.A1(_04708_),
    .A2(_04710_),
    .A3(_04711_),
    .B1(_04713_),
    .C1(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand3_1 _15394_ (.A(_13142_),
    .B(_13146_),
    .C(_13143_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _15395_ (.A(_13146_),
    .B(_13141_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand2_1 _15396_ (.A(_04752_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__nor3_2 _15397_ (.A(_13145_),
    .B(_04751_),
    .C(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__xnor2_4 _15398_ (.A(_13148_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__a31o_1 _15399_ (.A1(_13126_),
    .A2(_04717_),
    .A3(_04719_),
    .B1(_04562_),
    .X(_04757_));
 sky130_fd_sc_hd__nand2b_1 _15400_ (.A_N(_13131_),
    .B(_13130_),
    .Y(_04758_));
 sky130_fd_sc_hd__a311oi_2 _15401_ (.A1(_13126_),
    .A2(_04717_),
    .A3(_04719_),
    .B1(_04758_),
    .C1(_04562_),
    .Y(_04759_));
 sky130_fd_sc_hd__nor3_1 _15402_ (.A(_04636_),
    .B(_13132_),
    .C(_13131_),
    .Y(_04760_));
 sky130_fd_sc_hd__a21o_1 _15403_ (.A1(_04636_),
    .A2(_13131_),
    .B1(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__a311oi_4 _15404_ (.A1(_04757_),
    .A2(_13132_),
    .A3(_04636_),
    .B1(_04759_),
    .C1(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__nand3_2 _15405_ (.A(_13100_),
    .B(_13096_),
    .C(_13098_),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2b_1 _15406_ (.A(_04593_),
    .B_N(_13096_),
    .Y(_04764_));
 sky130_fd_sc_hd__nor2_2 _15407_ (.A(_13095_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__o21a_2 _15408_ (.A1(_04673_),
    .A2(_04763_),
    .B1(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__inv_1 _15409_ (.A(_13106_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _15410_ (.A(_04767_),
    .B(_13108_),
    .Y(_04768_));
 sky130_fd_sc_hd__inv_1 _15411_ (.A(_13107_),
    .Y(_04769_));
 sky130_fd_sc_hd__o2111ai_4 _15412_ (.A1(_04673_),
    .A2(_04763_),
    .B1(_13106_),
    .C1(_04769_),
    .D1(_04765_),
    .Y(_04770_));
 sky130_fd_sc_hd__nor3_1 _15413_ (.A(_04767_),
    .B(_13108_),
    .C(_13107_),
    .Y(_04771_));
 sky130_fd_sc_hd__a21oi_2 _15414_ (.A1(_04767_),
    .A2(_13107_),
    .B1(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__o211ai_4 _15415_ (.A1(_04766_),
    .A2(_04768_),
    .B1(_04770_),
    .C1(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__xnor2_2 _15416_ (.A(_04762_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__xnor2_4 _15417_ (.A(_04756_),
    .B(_04774_),
    .Y(_12318_));
 sky130_fd_sc_hd__maj3_1 _15418_ (.A(\hash.CA2.b_dash[8] ),
    .B(\hash.CA2.a_dash[8] ),
    .C(_04742_),
    .X(_04775_));
 sky130_fd_sc_hd__inv_1 _15419_ (.A(_04775_),
    .Y(_12329_));
 sky130_fd_sc_hd__nor3_1 _15420_ (.A(_13433_),
    .B(_13440_),
    .C(_13447_),
    .Y(_04776_));
 sky130_fd_sc_hd__or2_0 _15421_ (.A(_13441_),
    .B(_13440_),
    .X(_04777_));
 sky130_fd_sc_hd__a21oi_1 _15422_ (.A1(_13448_),
    .A2(_04777_),
    .B1(_13447_),
    .Y(_04778_));
 sky130_fd_sc_hd__a21oi_4 _15423_ (.A1(_04729_),
    .A2(_04776_),
    .B1(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__xor2_1 _15424_ (.A(_13455_),
    .B(_04779_),
    .X(_13456_));
 sky130_fd_sc_hd__inv_1 _15425_ (.A(_13456_),
    .Y(_12328_));
 sky130_fd_sc_hd__o21ai_2 _15426_ (.A1(_13145_),
    .A2(_04733_),
    .B1(_13148_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2b_2 _15427_ (.A_N(_13147_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__xnor2_4 _15428_ (.A(_04781_),
    .B(_13150_),
    .Y(_04782_));
 sky130_fd_sc_hd__nand3_1 _15429_ (.A(_13126_),
    .B(_13130_),
    .C(_13132_),
    .Y(_04783_));
 sky130_fd_sc_hd__nor2_1 _15430_ (.A(_04783_),
    .B(_04635_),
    .Y(_04784_));
 sky130_fd_sc_hd__nor4b_1 _15431_ (.A(_04783_),
    .B(_04584_),
    .C(_04587_),
    .D_N(_04609_),
    .Y(_04785_));
 sky130_fd_sc_hd__o41a_4 _15432_ (.A1(_13128_),
    .A2(_04638_),
    .A3(_04784_),
    .A4(_04785_),
    .B1(_04708_),
    .X(_04786_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1389 ();
 sky130_fd_sc_hd__nand2_4 _15434_ (.A(_04567_),
    .B(_04579_),
    .Y(_04788_));
 sky130_fd_sc_hd__a31o_1 _15435_ (.A1(_13108_),
    .A2(_04571_),
    .A3(_04578_),
    .B1(_13107_),
    .X(_04789_));
 sky130_fd_sc_hd__a211oi_4 _15436_ (.A1(_13106_),
    .A2(_04789_),
    .B1(_13105_),
    .C1(_13110_),
    .Y(_04790_));
 sky130_fd_sc_hd__nor2_8 _15437_ (.A(_04788_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__xnor2_2 _15438_ (.A(_04786_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__xnor2_4 _15439_ (.A(net1119),
    .B(_04792_),
    .Y(_12327_));
 sky130_fd_sc_hd__a21o_1 _15440_ (.A1(\hash.CA2.a_dash[9] ),
    .A2(_04773_),
    .B1(\hash.CA2.b_dash[9] ),
    .X(_04793_));
 sky130_fd_sc_hd__o21ai_1 _15441_ (.A1(\hash.CA2.a_dash[9] ),
    .A2(_04773_),
    .B1(_04793_),
    .Y(_12338_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(_13448_),
    .B(_13455_),
    .Y(_04794_));
 sky130_fd_sc_hd__a211o_1 _15443_ (.A1(_04728_),
    .A2(_04745_),
    .B1(_04794_),
    .C1(_04727_),
    .X(_04795_));
 sky130_fd_sc_hd__a21o_1 _15444_ (.A1(_13448_),
    .A2(_13440_),
    .B1(_13447_),
    .X(_04796_));
 sky130_fd_sc_hd__a21oi_1 _15445_ (.A1(_13455_),
    .A2(_04796_),
    .B1(_13454_),
    .Y(_04797_));
 sky130_fd_sc_hd__o21ai_1 _15446_ (.A1(_04747_),
    .A2(_04795_),
    .B1(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__xor2_1 _15447_ (.A(_13462_),
    .B(_04798_),
    .X(_13463_));
 sky130_fd_sc_hd__inv_1 _15448_ (.A(_13463_),
    .Y(_12337_));
 sky130_fd_sc_hd__xor2_2 _15449_ (.A(\hash.CA2.p1[31] ),
    .B(\hash.CA2.p3[31] ),
    .X(_04799_));
 sky130_fd_sc_hd__or3_1 _15450_ (.A(_13145_),
    .B(_13147_),
    .C(_13149_),
    .X(_04800_));
 sky130_fd_sc_hd__nor3_1 _15451_ (.A(_13148_),
    .B(_13147_),
    .C(_13149_),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _15452_ (.A(_13150_),
    .B(_13149_),
    .Y(_04802_));
 sky130_fd_sc_hd__nor2_1 _15453_ (.A(_04801_),
    .B(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__o31ai_4 _15454_ (.A1(_04751_),
    .A2(_04754_),
    .A3(_04800_),
    .B1(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__xnor2_4 _15455_ (.A(_04799_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__nand3_1 _15456_ (.A(_13108_),
    .B(_13112_),
    .C(_04565_),
    .Y(_04806_));
 sky130_fd_sc_hd__nor3_1 _15457_ (.A(_13112_),
    .B(_04565_),
    .C(_04597_),
    .Y(_04807_));
 sky130_fd_sc_hd__nand3_1 _15458_ (.A(_13112_),
    .B(_13107_),
    .C(_04565_),
    .Y(_04808_));
 sky130_fd_sc_hd__o41ai_1 _15459_ (.A1(_13108_),
    .A2(_13112_),
    .A3(_13107_),
    .A4(_04597_),
    .B1(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__a211oi_2 _15460_ (.A1(_13112_),
    .A2(_04597_),
    .B1(_04807_),
    .C1(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__nor3_1 _15461_ (.A(_13112_),
    .B(_13107_),
    .C(_04597_),
    .Y(_04811_));
 sky130_fd_sc_hd__o211ai_2 _15462_ (.A1(_04673_),
    .A2(_04763_),
    .B1(_04811_),
    .C1(_04765_),
    .Y(_04812_));
 sky130_fd_sc_hd__o211ai_4 _15463_ (.A1(_04766_),
    .A2(_04806_),
    .B1(_04810_),
    .C1(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__xnor2_1 _15464_ (.A(_04591_),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__xnor2_2 _15465_ (.A(_04805_),
    .B(_04814_),
    .Y(_12336_));
 sky130_fd_sc_hd__maj3_1 _15466_ (.A(\hash.CA2.b_dash[10] ),
    .B(\hash.CA2.a_dash[10] ),
    .C(_04791_),
    .X(_04815_));
 sky130_fd_sc_hd__inv_1 _15467_ (.A(_04815_),
    .Y(_12347_));
 sky130_fd_sc_hd__a21o_1 _15468_ (.A1(_13455_),
    .A2(_04779_),
    .B1(_13454_),
    .X(_04816_));
 sky130_fd_sc_hd__a21o_1 _15469_ (.A1(_13462_),
    .A2(_04816_),
    .B1(_13461_),
    .X(_04817_));
 sky130_fd_sc_hd__xor2_1 _15470_ (.A(_13469_),
    .B(_04817_),
    .X(_13470_));
 sky130_fd_sc_hd__inv_1 _15471_ (.A(_13470_),
    .Y(_12346_));
 sky130_fd_sc_hd__nor2b_1 _15472_ (.A(_13116_),
    .B_N(_13112_),
    .Y(_04818_));
 sky130_fd_sc_hd__a21oi_1 _15473_ (.A1(_13112_),
    .A2(_13109_),
    .B1(_13111_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _15474_ (.A(_13116_),
    .B(_04582_),
    .Y(_04820_));
 sky130_fd_sc_hd__o21ai_1 _15475_ (.A1(_13116_),
    .A2(_04819_),
    .B1(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__nor2_1 _15476_ (.A(_13109_),
    .B(_13111_),
    .Y(_04822_));
 sky130_fd_sc_hd__and4_1 _15477_ (.A(_13116_),
    .B(_04567_),
    .C(_04579_),
    .D(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__a211oi_4 _15478_ (.A1(_04818_),
    .A2(_04788_),
    .B1(_04821_),
    .C1(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__xnor2_1 _15479_ (.A(_13090_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__xnor2_1 _15480_ (.A(_04643_),
    .B(_04825_),
    .Y(_12345_));
 sky130_fd_sc_hd__clkinvlp_4 _15481_ (.A(\hash.CA2.b_dash[11] ),
    .Y(_04826_));
 sky130_fd_sc_hd__inv_1 _15482_ (.A(\hash.CA2.a_dash[11] ),
    .Y(_04827_));
 sky130_fd_sc_hd__maj3_1 _15483_ (.A(_04826_),
    .B(_04827_),
    .C(_04813_),
    .X(_12356_));
 sky130_fd_sc_hd__o21ai_0 _15484_ (.A1(_13462_),
    .A2(_13461_),
    .B1(_13469_),
    .Y(_04828_));
 sky130_fd_sc_hd__nand2b_1 _15485_ (.A_N(_13468_),
    .B(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__o31a_2 _15486_ (.A1(_13461_),
    .A2(_13468_),
    .A3(_04798_),
    .B1(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__xor2_1 _15487_ (.A(_13476_),
    .B(_04830_),
    .X(_13477_));
 sky130_fd_sc_hd__inv_1 _15488_ (.A(_13477_),
    .Y(_12355_));
 sky130_fd_sc_hd__xnor2_1 _15489_ (.A(_12253_),
    .B(_04611_),
    .Y(_04831_));
 sky130_fd_sc_hd__xnor2_1 _15490_ (.A(net1135),
    .B(_04831_),
    .Y(_12354_));
 sky130_fd_sc_hd__inv_1 _15491_ (.A(\hash.CA2.b_dash[12] ),
    .Y(_04832_));
 sky130_fd_sc_hd__inv_1 _15492_ (.A(\hash.CA2.a_dash[12] ),
    .Y(_04833_));
 sky130_fd_sc_hd__maj3_1 _15493_ (.A(_04832_),
    .B(_04833_),
    .C(net1161),
    .X(_12365_));
 sky130_fd_sc_hd__and4_1 _15494_ (.A(_13455_),
    .B(_13462_),
    .C(_13469_),
    .D(_13476_),
    .X(_04834_));
 sky130_fd_sc_hd__a21o_1 _15495_ (.A1(_13469_),
    .A2(_13461_),
    .B1(_13468_),
    .X(_04835_));
 sky130_fd_sc_hd__a21oi_1 _15496_ (.A1(_13476_),
    .A2(_04835_),
    .B1(_13475_),
    .Y(_04836_));
 sky130_fd_sc_hd__nand4_1 _15497_ (.A(_13462_),
    .B(_13469_),
    .C(_13476_),
    .D(_13454_),
    .Y(_04837_));
 sky130_fd_sc_hd__nand2_1 _15498_ (.A(_04836_),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21oi_4 _15499_ (.A1(_04834_),
    .A2(_04779_),
    .B1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__xnor2_1 _15500_ (.A(_13483_),
    .B(_04839_),
    .Y(_13484_));
 sky130_fd_sc_hd__inv_1 _15501_ (.A(_13484_),
    .Y(_12364_));
 sky130_fd_sc_hd__xnor2_4 _15502_ (.A(_13092_),
    .B(net1136),
    .Y(_04840_));
 sky130_fd_sc_hd__xnor2_1 _15503_ (.A(_04840_),
    .B(_04627_),
    .Y(_04841_));
 sky130_fd_sc_hd__xnor2_1 _15504_ (.A(net1166),
    .B(_04841_),
    .Y(_12363_));
 sky130_fd_sc_hd__xor2_4 _15505_ (.A(_13114_),
    .B(_04610_),
    .X(_04842_));
 sky130_fd_sc_hd__nor2_1 _15506_ (.A(\hash.CA2.a_dash[13] ),
    .B(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__a21oi_1 _15507_ (.A1(\hash.CA2.a_dash[13] ),
    .A2(_04842_),
    .B1(\hash.CA2.b_dash[13] ),
    .Y(_04844_));
 sky130_fd_sc_hd__nor2_1 _15508_ (.A(_04843_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__inv_1 _15509_ (.A(_04845_),
    .Y(_12374_));
 sky130_fd_sc_hd__inv_1 _15510_ (.A(_13483_),
    .Y(_04846_));
 sky130_fd_sc_hd__a21oi_1 _15511_ (.A1(_13476_),
    .A2(_04830_),
    .B1(_13475_),
    .Y(_04847_));
 sky130_fd_sc_hd__o21bai_1 _15512_ (.A1(_04846_),
    .A2(_04847_),
    .B1_N(_13482_),
    .Y(_04848_));
 sky130_fd_sc_hd__xor2_1 _15513_ (.A(_13490_),
    .B(_04848_),
    .X(_13491_));
 sky130_fd_sc_hd__inv_1 _15514_ (.A(_13491_),
    .Y(_12373_));
 sky130_fd_sc_hd__xnor2_1 _15515_ (.A(_04646_),
    .B(_04659_),
    .Y(_04849_));
 sky130_fd_sc_hd__xnor2_2 _15516_ (.A(_04849_),
    .B(_04694_),
    .Y(_12372_));
 sky130_fd_sc_hd__nor2_1 _15517_ (.A(\hash.CA2.a_dash[14] ),
    .B(_04627_),
    .Y(_04850_));
 sky130_fd_sc_hd__a21oi_1 _15518_ (.A1(\hash.CA2.a_dash[14] ),
    .A2(_04627_),
    .B1(\hash.CA2.b_dash[14] ),
    .Y(_04851_));
 sky130_fd_sc_hd__or2_0 _15519_ (.A(_04850_),
    .B(_04851_),
    .X(_12383_));
 sky130_fd_sc_hd__o21bai_1 _15520_ (.A1(_04846_),
    .A2(_04839_),
    .B1_N(_13482_),
    .Y(_04852_));
 sky130_fd_sc_hd__a21oi_1 _15521_ (.A1(_13490_),
    .A2(_04852_),
    .B1(_13489_),
    .Y(_04853_));
 sky130_fd_sc_hd__xnor2_1 _15522_ (.A(net1114),
    .B(_04853_),
    .Y(_13498_));
 sky130_fd_sc_hd__inv_1 _15523_ (.A(_13498_),
    .Y(_12382_));
 sky130_fd_sc_hd__xnor2_1 _15524_ (.A(_04654_),
    .B(_04672_),
    .Y(_04854_));
 sky130_fd_sc_hd__xnor2_1 _15525_ (.A(_04716_),
    .B(_04854_),
    .Y(_12381_));
 sky130_fd_sc_hd__maj3_1 _15526_ (.A(\hash.CA2.b_dash[15] ),
    .B(\hash.CA2.a_dash[15] ),
    .C(_04659_),
    .X(_04855_));
 sky130_fd_sc_hd__inv_1 _15527_ (.A(_04855_),
    .Y(_12392_));
 sky130_fd_sc_hd__and3_1 _15528_ (.A(_13483_),
    .B(_13490_),
    .C(_13497_),
    .X(_04856_));
 sky130_fd_sc_hd__inv_2 _15529_ (.A(_13497_),
    .Y(_04857_));
 sky130_fd_sc_hd__a21o_1 _15530_ (.A1(_13483_),
    .A2(_13475_),
    .B1(_13482_),
    .X(_04858_));
 sky130_fd_sc_hd__a21oi_1 _15531_ (.A1(_13490_),
    .A2(_04858_),
    .B1(_13489_),
    .Y(_04859_));
 sky130_fd_sc_hd__o21bai_1 _15532_ (.A1(_04857_),
    .A2(_04859_),
    .B1_N(_13496_),
    .Y(_04860_));
 sky130_fd_sc_hd__a31oi_4 _15533_ (.A1(_13476_),
    .A2(_04856_),
    .A3(_04830_),
    .B1(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__xnor2_1 _15534_ (.A(_13504_),
    .B(net1105),
    .Y(_13505_));
 sky130_fd_sc_hd__inv_1 _15535_ (.A(_13505_),
    .Y(_12391_));
 sky130_fd_sc_hd__xor2_1 _15536_ (.A(_04674_),
    .B(_04699_),
    .X(_04862_));
 sky130_fd_sc_hd__xnor2_1 _15537_ (.A(_04736_),
    .B(_04862_),
    .Y(_12390_));
 sky130_fd_sc_hd__inv_1 _15538_ (.A(\hash.CA2.b_dash[16] ),
    .Y(_04863_));
 sky130_fd_sc_hd__inv_1 _15539_ (.A(\hash.CA2.a_dash[16] ),
    .Y(_04864_));
 sky130_fd_sc_hd__maj3_1 _15540_ (.A(_04863_),
    .B(_04864_),
    .C(net1130),
    .X(_12401_));
 sky130_fd_sc_hd__nand3_2 _15541_ (.A(_13483_),
    .B(_13490_),
    .C(_13497_),
    .Y(_04865_));
 sky130_fd_sc_hd__a21oi_1 _15542_ (.A1(_13490_),
    .A2(_13482_),
    .B1(_13489_),
    .Y(_04866_));
 sky130_fd_sc_hd__o22ai_4 _15543_ (.A1(_04865_),
    .A2(_04839_),
    .B1(_04866_),
    .B2(_04857_),
    .Y(_04867_));
 sky130_fd_sc_hd__o21ai_0 _15544_ (.A1(_13496_),
    .A2(_04867_),
    .B1(_13504_),
    .Y(_04868_));
 sky130_fd_sc_hd__nor2b_1 _15545_ (.A(_13503_),
    .B_N(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__xnor2_2 _15546_ (.A(_13511_),
    .B(_04869_),
    .Y(_13512_));
 sky130_fd_sc_hd__inv_1 _15547_ (.A(_13512_),
    .Y(_12400_));
 sky130_fd_sc_hd__xor2_1 _15548_ (.A(_04701_),
    .B(_04721_),
    .X(_04870_));
 sky130_fd_sc_hd__xnor2_1 _15549_ (.A(_04756_),
    .B(_04870_),
    .Y(_12399_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1388 ();
 sky130_fd_sc_hd__nor2_1 _15551_ (.A(\hash.CA2.a_dash[17] ),
    .B(_04699_),
    .Y(_04872_));
 sky130_fd_sc_hd__a21oi_1 _15552_ (.A1(\hash.CA2.a_dash[17] ),
    .A2(_04699_),
    .B1(\hash.CA2.b_dash[17] ),
    .Y(_04873_));
 sky130_fd_sc_hd__nor2_1 _15553_ (.A(_04872_),
    .B(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__inv_1 _15554_ (.A(_04874_),
    .Y(_12410_));
 sky130_fd_sc_hd__nor2b_1 _15555_ (.A(_04861_),
    .B_N(_13504_),
    .Y(_04875_));
 sky130_fd_sc_hd__o21ai_0 _15556_ (.A1(_13503_),
    .A2(_04875_),
    .B1(_13511_),
    .Y(_04876_));
 sky130_fd_sc_hd__nand2b_1 _15557_ (.A_N(_13510_),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__xor2_2 _15558_ (.A(_13518_),
    .B(_04877_),
    .X(_13519_));
 sky130_fd_sc_hd__inv_1 _15559_ (.A(_13519_),
    .Y(_12409_));
 sky130_fd_sc_hd__xor2_2 _15560_ (.A(_13132_),
    .B(_04739_),
    .X(_04878_));
 sky130_fd_sc_hd__xnor2_1 _15561_ (.A(_04724_),
    .B(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__xnor2_1 _15562_ (.A(net1119),
    .B(_04879_),
    .Y(_12408_));
 sky130_fd_sc_hd__nor2_1 _15563_ (.A(\hash.CA2.a_dash[18] ),
    .B(_04721_),
    .Y(_04880_));
 sky130_fd_sc_hd__a21oi_1 _15564_ (.A1(\hash.CA2.a_dash[18] ),
    .A2(_04721_),
    .B1(\hash.CA2.b_dash[18] ),
    .Y(_04881_));
 sky130_fd_sc_hd__nor2_1 _15565_ (.A(_04880_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__inv_1 _15566_ (.A(_04882_),
    .Y(_12419_));
 sky130_fd_sc_hd__inv_1 _15567_ (.A(_13525_),
    .Y(_04883_));
 sky130_fd_sc_hd__a21o_1 _15568_ (.A1(_13504_),
    .A2(_13496_),
    .B1(_13503_),
    .X(_04884_));
 sky130_fd_sc_hd__a21o_1 _15569_ (.A1(_13511_),
    .A2(_04884_),
    .B1(_13510_),
    .X(_04885_));
 sky130_fd_sc_hd__a31o_1 _15570_ (.A1(_04867_),
    .A2(_13511_),
    .A3(_13504_),
    .B1(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__a21o_1 _15571_ (.A1(_04886_),
    .A2(_13518_),
    .B1(_13517_),
    .X(_04887_));
 sky130_fd_sc_hd__xnor2_1 _15572_ (.A(_04883_),
    .B(_04887_),
    .Y(_13526_));
 sky130_fd_sc_hd__inv_1 _15573_ (.A(_13526_),
    .Y(_12418_));
 sky130_fd_sc_hd__xnor2_1 _15574_ (.A(_04742_),
    .B(net1138),
    .Y(_04888_));
 sky130_fd_sc_hd__xnor2_1 _15575_ (.A(_04805_),
    .B(_04888_),
    .Y(_12417_));
 sky130_fd_sc_hd__maj3_1 _15576_ (.A(\hash.CA2.b_dash[19] ),
    .B(\hash.CA2.a_dash[19] ),
    .C(_04878_),
    .X(_04889_));
 sky130_fd_sc_hd__inv_1 _15577_ (.A(_04889_),
    .Y(_12428_));
 sky130_fd_sc_hd__nand3_1 _15578_ (.A(_13504_),
    .B(_13511_),
    .C(_13518_),
    .Y(_04890_));
 sky130_fd_sc_hd__a21o_1 _15579_ (.A1(_13511_),
    .A2(_13503_),
    .B1(_13510_),
    .X(_04891_));
 sky130_fd_sc_hd__a21oi_1 _15580_ (.A1(_13518_),
    .A2(_04891_),
    .B1(_13517_),
    .Y(_04892_));
 sky130_fd_sc_hd__o21ai_0 _15581_ (.A1(_04861_),
    .A2(_04890_),
    .B1(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__a21oi_2 _15582_ (.A1(_04893_),
    .A2(_13525_),
    .B1(_13524_),
    .Y(_04894_));
 sky130_fd_sc_hd__xnor2_1 _15583_ (.A(_13532_),
    .B(_04894_),
    .Y(_13533_));
 sky130_fd_sc_hd__inv_1 _15584_ (.A(_13533_),
    .Y(_12427_));
 sky130_fd_sc_hd__o211a_4 _15585_ (.A1(_04766_),
    .A2(_04768_),
    .B1(_04770_),
    .C1(_04772_),
    .X(_04895_));
 sky130_fd_sc_hd__xnor2_2 _15586_ (.A(_13090_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__xnor2_1 _15587_ (.A(_04786_),
    .B(_04896_),
    .Y(_12426_));
 sky130_fd_sc_hd__inv_1 _15588_ (.A(\hash.CA2.b_dash[20] ),
    .Y(_04897_));
 sky130_fd_sc_hd__inv_1 _15589_ (.A(\hash.CA2.a_dash[20] ),
    .Y(_04898_));
 sky130_fd_sc_hd__maj3_1 _15590_ (.A(_04897_),
    .B(_04898_),
    .C(net1139),
    .X(_12437_));
 sky130_fd_sc_hd__inv_1 _15591_ (.A(_13539_),
    .Y(_04899_));
 sky130_fd_sc_hd__inv_1 _15592_ (.A(_13532_),
    .Y(_04900_));
 sky130_fd_sc_hd__a21oi_2 _15593_ (.A1(_04887_),
    .A2(_13525_),
    .B1(_13524_),
    .Y(_04901_));
 sky130_fd_sc_hd__o21bai_1 _15594_ (.A1(_04900_),
    .A2(net1115),
    .B1_N(_13531_),
    .Y(_04902_));
 sky130_fd_sc_hd__xnor2_2 _15595_ (.A(_04902_),
    .B(_04899_),
    .Y(_13540_));
 sky130_fd_sc_hd__inv_1 _15596_ (.A(_13540_),
    .Y(_12436_));
 sky130_fd_sc_hd__xnor2_1 _15597_ (.A(_12253_),
    .B(_04791_),
    .Y(_04903_));
 sky130_fd_sc_hd__xor2_1 _15598_ (.A(_04591_),
    .B(_04903_),
    .X(_12435_));
 sky130_fd_sc_hd__maj3_1 _15599_ (.A(\hash.CA2.b_dash[21] ),
    .B(\hash.CA2.a_dash[21] ),
    .C(_04786_),
    .X(_04904_));
 sky130_fd_sc_hd__inv_1 _15600_ (.A(_04904_),
    .Y(_12446_));
 sky130_fd_sc_hd__inv_1 _15601_ (.A(_13538_),
    .Y(_04905_));
 sky130_fd_sc_hd__nor2_1 _15602_ (.A(_04900_),
    .B(_04894_),
    .Y(_04906_));
 sky130_fd_sc_hd__o21ai_0 _15603_ (.A1(_13531_),
    .A2(_04906_),
    .B1(_13539_),
    .Y(_04907_));
 sky130_fd_sc_hd__nand2_1 _15604_ (.A(_04905_),
    .B(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__xor2_2 _15605_ (.A(_13546_),
    .B(_04908_),
    .X(_13547_));
 sky130_fd_sc_hd__inv_1 _15606_ (.A(_13547_),
    .Y(_12445_));
 sky130_fd_sc_hd__xnor2_2 _15607_ (.A(_04592_),
    .B(_04813_),
    .Y(_04909_));
 sky130_fd_sc_hd__xnor2_4 _15608_ (.A(net1170),
    .B(_04909_),
    .Y(_12444_));
 sky130_fd_sc_hd__nor2_1 _15609_ (.A(\hash.CA2.a_dash[22] ),
    .B(net1121),
    .Y(_04910_));
 sky130_fd_sc_hd__a21oi_1 _15610_ (.A1(\hash.CA2.a_dash[22] ),
    .A2(net1121),
    .B1(\hash.CA2.b_dash[22] ),
    .Y(_04911_));
 sky130_fd_sc_hd__nor2_1 _15611_ (.A(_04910_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__inv_1 _15612_ (.A(_04912_),
    .Y(_12455_));
 sky130_fd_sc_hd__nand2_1 _15613_ (.A(_13532_),
    .B(_13539_),
    .Y(_04913_));
 sky130_fd_sc_hd__nand2_1 _15614_ (.A(_13539_),
    .B(_13531_),
    .Y(_04914_));
 sky130_fd_sc_hd__o211ai_2 _15615_ (.A1(_04913_),
    .A2(_04901_),
    .B1(_04914_),
    .C1(_04905_),
    .Y(_04915_));
 sky130_fd_sc_hd__a21oi_4 _15616_ (.A1(_13546_),
    .A2(_04915_),
    .B1(_13545_),
    .Y(_04916_));
 sky130_fd_sc_hd__xor2_2 _15617_ (.A(_13553_),
    .B(_04916_),
    .X(_12454_));
 sky130_fd_sc_hd__xor2_1 _15618_ (.A(_04646_),
    .B(net1159),
    .X(_04917_));
 sky130_fd_sc_hd__xnor2_1 _15619_ (.A(net1135),
    .B(_04917_),
    .Y(_12453_));
 sky130_fd_sc_hd__maj3_1 _15620_ (.A(\hash.CA2.b_dash[23] ),
    .B(\hash.CA2.a_dash[23] ),
    .C(net1167),
    .X(_04918_));
 sky130_fd_sc_hd__inv_1 _15621_ (.A(_04918_),
    .Y(_12464_));
 sky130_fd_sc_hd__nand2_1 _15622_ (.A(_13546_),
    .B(_13553_),
    .Y(_04919_));
 sky130_fd_sc_hd__or3_1 _15623_ (.A(_04883_),
    .B(_04913_),
    .C(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__nor2_1 _15624_ (.A(_04890_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__inv_1 _15625_ (.A(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__nor2_1 _15626_ (.A(_13524_),
    .B(_13531_),
    .Y(_04923_));
 sky130_fd_sc_hd__o21ai_0 _15627_ (.A1(_04883_),
    .A2(_04892_),
    .B1(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__o211ai_1 _15628_ (.A1(_13532_),
    .A2(_13531_),
    .B1(_04924_),
    .C1(_13539_),
    .Y(_04925_));
 sky130_fd_sc_hd__nor3_1 _15629_ (.A(_13538_),
    .B(_13545_),
    .C(_13552_),
    .Y(_04926_));
 sky130_fd_sc_hd__or2_0 _15630_ (.A(_13546_),
    .B(_13545_),
    .X(_04927_));
 sky130_fd_sc_hd__a21oi_1 _15631_ (.A1(_13553_),
    .A2(_04927_),
    .B1(_13552_),
    .Y(_04928_));
 sky130_fd_sc_hd__a21oi_1 _15632_ (.A1(_04925_),
    .A2(_04926_),
    .B1(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__o21bai_4 _15633_ (.A1(net1104),
    .A2(_04922_),
    .B1_N(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__xor2_1 _15634_ (.A(_13560_),
    .B(_04930_),
    .X(_13561_));
 sky130_fd_sc_hd__inv_1 _15635_ (.A(_13561_),
    .Y(_12463_));
 sky130_fd_sc_hd__xnor2_2 _15636_ (.A(_04611_),
    .B(_04654_),
    .Y(_04931_));
 sky130_fd_sc_hd__xnor2_1 _15637_ (.A(net1166),
    .B(_04931_),
    .Y(_12462_));
 sky130_fd_sc_hd__nand2_1 _15638_ (.A(\hash.CA2.a_dash[24] ),
    .B(_04652_),
    .Y(_04932_));
 sky130_fd_sc_hd__o21ai_0 _15639_ (.A1(\hash.CA2.a_dash[24] ),
    .A2(_04652_),
    .B1(\hash.CA2.b_dash[24] ),
    .Y(_04933_));
 sky130_fd_sc_hd__nand2_1 _15640_ (.A(_04932_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__inv_1 _15641_ (.A(_04934_),
    .Y(_12473_));
 sky130_fd_sc_hd__a21oi_1 _15642_ (.A1(_13518_),
    .A2(_04885_),
    .B1(_13517_),
    .Y(_04935_));
 sky130_fd_sc_hd__a21oi_1 _15643_ (.A1(_13532_),
    .A2(_13524_),
    .B1(_13531_),
    .Y(_04936_));
 sky130_fd_sc_hd__o21ai_0 _15644_ (.A1(_04899_),
    .A2(_04936_),
    .B1(_04905_),
    .Y(_04937_));
 sky130_fd_sc_hd__a21o_1 _15645_ (.A1(_13546_),
    .A2(_04937_),
    .B1(_13545_),
    .X(_04938_));
 sky130_fd_sc_hd__a21oi_1 _15646_ (.A1(_13553_),
    .A2(_04938_),
    .B1(_13552_),
    .Y(_04939_));
 sky130_fd_sc_hd__o21ai_0 _15647_ (.A1(_04920_),
    .A2(_04935_),
    .B1(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__a21o_1 _15648_ (.A1(_04867_),
    .A2(_04921_),
    .B1(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__a21oi_1 _15649_ (.A1(_13560_),
    .A2(_04941_),
    .B1(_13559_),
    .Y(_04942_));
 sky130_fd_sc_hd__xnor2_1 _15650_ (.A(_13567_),
    .B(_04942_),
    .Y(_13568_));
 sky130_fd_sc_hd__inv_1 _15651_ (.A(_13568_),
    .Y(_12472_));
 sky130_fd_sc_hd__xor2_4 _15652_ (.A(_04627_),
    .B(_04674_),
    .X(_04943_));
 sky130_fd_sc_hd__xnor2_1 _15653_ (.A(_04694_),
    .B(_04943_),
    .Y(_12471_));
 sky130_fd_sc_hd__maj3_1 _15654_ (.A(\hash.CA2.b_dash[25] ),
    .B(\hash.CA2.a_dash[25] ),
    .C(_04667_),
    .X(_04944_));
 sky130_fd_sc_hd__inv_1 _15655_ (.A(_04944_),
    .Y(_12482_));
 sky130_fd_sc_hd__a21o_1 _15656_ (.A1(_13560_),
    .A2(_04930_),
    .B1(_13559_),
    .X(_04945_));
 sky130_fd_sc_hd__a21o_1 _15657_ (.A1(_13567_),
    .A2(_04945_),
    .B1(_13566_),
    .X(_04946_));
 sky130_fd_sc_hd__xor2_2 _15658_ (.A(_13574_),
    .B(_04946_),
    .X(_13575_));
 sky130_fd_sc_hd__inv_1 _15659_ (.A(_13575_),
    .Y(_12481_));
 sky130_fd_sc_hd__xor2_2 _15660_ (.A(_04659_),
    .B(_04701_),
    .X(_04947_));
 sky130_fd_sc_hd__xnor2_1 _15661_ (.A(_04716_),
    .B(_04947_),
    .Y(_12480_));
 sky130_fd_sc_hd__maj3_1 _15662_ (.A(\hash.CA2.b_dash[26] ),
    .B(\hash.CA2.a_dash[26] ),
    .C(_04694_),
    .X(_04948_));
 sky130_fd_sc_hd__inv_1 _15663_ (.A(_04948_),
    .Y(_12491_));
 sky130_fd_sc_hd__and3_1 _15664_ (.A(_13560_),
    .B(_13567_),
    .C(_13574_),
    .X(_04949_));
 sky130_fd_sc_hd__a21o_1 _15665_ (.A1(_13567_),
    .A2(_13559_),
    .B1(_13566_),
    .X(_04950_));
 sky130_fd_sc_hd__a21oi_2 _15666_ (.A1(_13574_),
    .A2(_04950_),
    .B1(_13573_),
    .Y(_04951_));
 sky130_fd_sc_hd__a21boi_2 _15667_ (.A1(_04941_),
    .A2(_04949_),
    .B1_N(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__xnor2_1 _15668_ (.A(_13581_),
    .B(_04952_),
    .Y(_13582_));
 sky130_fd_sc_hd__inv_1 _15669_ (.A(_13582_),
    .Y(_12490_));
 sky130_fd_sc_hd__xnor2_2 _15670_ (.A(net1131),
    .B(_04724_),
    .Y(_04953_));
 sky130_fd_sc_hd__xnor2_1 _15671_ (.A(_04736_),
    .B(_04953_),
    .Y(_12489_));
 sky130_fd_sc_hd__nand2_1 _15672_ (.A(\hash.CA2.a_dash[27] ),
    .B(_04716_),
    .Y(_04954_));
 sky130_fd_sc_hd__o21ai_0 _15673_ (.A1(\hash.CA2.a_dash[27] ),
    .A2(_04716_),
    .B1(\hash.CA2.b_dash[27] ),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _15674_ (.A(_04954_),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__inv_1 _15675_ (.A(_04956_),
    .Y(_12500_));
 sky130_fd_sc_hd__a21bo_1 _15676_ (.A1(_04930_),
    .A2(_04949_),
    .B1_N(_04951_),
    .X(_04957_));
 sky130_fd_sc_hd__a21oi_1 _15677_ (.A1(_13581_),
    .A2(_04957_),
    .B1(_13580_),
    .Y(_04958_));
 sky130_fd_sc_hd__xnor2_1 _15678_ (.A(_13588_),
    .B(_04958_),
    .Y(_13589_));
 sky130_fd_sc_hd__inv_1 _15679_ (.A(_13589_),
    .Y(_12499_));
 sky130_fd_sc_hd__xor2_2 _15680_ (.A(_04699_),
    .B(_04742_),
    .X(_04959_));
 sky130_fd_sc_hd__xnor2_1 _15681_ (.A(_04756_),
    .B(_04959_),
    .Y(_12498_));
 sky130_fd_sc_hd__nor2_1 _15682_ (.A(\hash.CA2.a_dash[28] ),
    .B(_04736_),
    .Y(_04960_));
 sky130_fd_sc_hd__a21oi_1 _15683_ (.A1(\hash.CA2.a_dash[28] ),
    .A2(_04736_),
    .B1(\hash.CA2.b_dash[28] ),
    .Y(_04961_));
 sky130_fd_sc_hd__nor2_1 _15684_ (.A(_04960_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__inv_1 _15685_ (.A(_04962_),
    .Y(_12509_));
 sky130_fd_sc_hd__nand2_1 _15686_ (.A(_13581_),
    .B(_13588_),
    .Y(_04963_));
 sky130_fd_sc_hd__nand2_1 _15687_ (.A(_13588_),
    .B(_13580_),
    .Y(_04964_));
 sky130_fd_sc_hd__inv_1 _15688_ (.A(_13587_),
    .Y(_04965_));
 sky130_fd_sc_hd__o211ai_1 _15689_ (.A1(_04952_),
    .A2(_04963_),
    .B1(_04964_),
    .C1(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__xor2_1 _15690_ (.A(_13595_),
    .B(_04966_),
    .X(_13596_));
 sky130_fd_sc_hd__inv_1 _15691_ (.A(_13596_),
    .Y(_12508_));
 sky130_fd_sc_hd__xnor2_2 _15692_ (.A(_04721_),
    .B(_04773_),
    .Y(_04967_));
 sky130_fd_sc_hd__xnor2_1 _15693_ (.A(net1119),
    .B(_04967_),
    .Y(_12507_));
 sky130_fd_sc_hd__maj3_1 _15694_ (.A(\hash.CA2.b_dash[29] ),
    .B(\hash.CA2.a_dash[29] ),
    .C(_04756_),
    .X(_04968_));
 sky130_fd_sc_hd__inv_1 _15695_ (.A(_04968_),
    .Y(_12518_));
 sky130_fd_sc_hd__nand3_1 _15696_ (.A(_13560_),
    .B(_13567_),
    .C(_13574_),
    .Y(_04969_));
 sky130_fd_sc_hd__nor2_1 _15697_ (.A(_04969_),
    .B(_04963_),
    .Y(_04970_));
 sky130_fd_sc_hd__o21ai_1 _15698_ (.A1(_04951_),
    .A2(_04963_),
    .B1(_04964_),
    .Y(_04971_));
 sky130_fd_sc_hd__a21oi_2 _15699_ (.A1(_04930_),
    .A2(_04970_),
    .B1(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_1 _15700_ (.A(_04965_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__a21o_1 _15701_ (.A1(_13595_),
    .A2(_04973_),
    .B1(_13594_),
    .X(_04974_));
 sky130_fd_sc_hd__xor2_1 _15702_ (.A(_13602_),
    .B(_04974_),
    .X(_13603_));
 sky130_fd_sc_hd__inv_1 _15703_ (.A(_13603_),
    .Y(_12517_));
 sky130_fd_sc_hd__xnor2_2 _15704_ (.A(_04740_),
    .B(_04791_),
    .Y(_04975_));
 sky130_fd_sc_hd__xnor2_1 _15705_ (.A(_04805_),
    .B(_04975_),
    .Y(_12516_));
 sky130_fd_sc_hd__inv_1 _15706_ (.A(\hash.CA2.a_dash[30] ),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2_1 _15707_ (.A(_04976_),
    .B(net1119),
    .Y(_04977_));
 sky130_fd_sc_hd__nor2_1 _15708_ (.A(_04976_),
    .B(net1119),
    .Y(_04978_));
 sky130_fd_sc_hd__a21oi_1 _15709_ (.A1(\hash.CA2.b_dash[30] ),
    .A2(_04977_),
    .B1(_04978_),
    .Y(_12527_));
 sky130_fd_sc_hd__a21o_1 _15710_ (.A1(_13595_),
    .A2(_04966_),
    .B1(_13594_),
    .X(_04979_));
 sky130_fd_sc_hd__a21o_1 _15711_ (.A1(_13602_),
    .A2(_04979_),
    .B1(_13601_),
    .X(_04980_));
 sky130_fd_sc_hd__xnor2_2 _15712_ (.A(_13609_),
    .B(_04980_),
    .Y(_12526_));
 sky130_fd_sc_hd__xor2_4 _15713_ (.A(_13090_),
    .B(_04813_),
    .X(_04981_));
 sky130_fd_sc_hd__xnor2_2 _15714_ (.A(net1139),
    .B(_04981_),
    .Y(_12525_));
 sky130_fd_sc_hd__nor2_8 _15715_ (.A(\hash.reset ),
    .B(_13613_),
    .Y(_00781_));
 sky130_fd_sc_hd__nor2b_4 _15716_ (.A(net762),
    .B_N(_13696_),
    .Y(_04982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1387 ();
 sky130_fd_sc_hd__nand2_8 _15718_ (.A(_09897_),
    .B(_04982_),
    .Y(_04984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1384 ();
 sky130_fd_sc_hd__mux2i_4 _15722_ (.A0(_13154_),
    .A1(\w[62][0] ),
    .S(net530),
    .Y(_04988_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1382 ();
 sky130_fd_sc_hd__nand2_1 _15725_ (.A(net245),
    .B(_04984_),
    .Y(_04991_));
 sky130_fd_sc_hd__o21ai_0 _15726_ (.A1(_04984_),
    .A2(_04988_),
    .B1(_04991_),
    .Y(_00129_));
 sky130_fd_sc_hd__mux2i_4 _15727_ (.A0(_13157_),
    .A1(\w[62][1] ),
    .S(net529),
    .Y(_04992_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1381 ();
 sky130_fd_sc_hd__nand2_1 _15729_ (.A(net234),
    .B(_04984_),
    .Y(_04994_));
 sky130_fd_sc_hd__o21ai_0 _15730_ (.A1(_04984_),
    .A2(_04992_),
    .B1(_04994_),
    .Y(_00140_));
 sky130_fd_sc_hd__mux2i_4 _15731_ (.A0(_11773_),
    .A1(\w[62][2] ),
    .S(net527),
    .Y(_04995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1380 ();
 sky130_fd_sc_hd__nand2_1 _15733_ (.A(net222),
    .B(_04984_),
    .Y(_04997_));
 sky130_fd_sc_hd__o21ai_0 _15734_ (.A1(_04984_),
    .A2(_04995_),
    .B1(_04997_),
    .Y(_00151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1378 ();
 sky130_fd_sc_hd__nor2b_1 _15737_ (.A(_13165_),
    .B_N(_11772_),
    .Y(_05000_));
 sky130_fd_sc_hd__nor2b_1 _15738_ (.A(_11772_),
    .B_N(_13165_),
    .Y(_05001_));
 sky130_fd_sc_hd__nor3_2 _15739_ (.A(net530),
    .B(_05000_),
    .C(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__a21oi_4 _15740_ (.A1(\w[62][3] ),
    .A2(net530),
    .B1(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1377 ();
 sky130_fd_sc_hd__nand2_1 _15742_ (.A(net211),
    .B(_04984_),
    .Y(_05005_));
 sky130_fd_sc_hd__o21ai_0 _15743_ (.A1(_04984_),
    .A2(_05003_),
    .B1(_05005_),
    .Y(_00154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1376 ();
 sky130_fd_sc_hd__inv_1 _15745_ (.A(_13169_),
    .Y(_05007_));
 sky130_fd_sc_hd__a21o_1 _15746_ (.A1(_13156_),
    .A2(_13161_),
    .B1(_13160_),
    .X(_05008_));
 sky130_fd_sc_hd__a21oi_2 _15747_ (.A1(_13165_),
    .A2(_05008_),
    .B1(_13164_),
    .Y(_05009_));
 sky130_fd_sc_hd__xnor2_1 _15748_ (.A(_05007_),
    .B(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__nor2_2 _15749_ (.A(net530),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__a21oi_4 _15750_ (.A1(\w[62][4] ),
    .A2(net531),
    .B1(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1375 ();
 sky130_fd_sc_hd__nand2_1 _15752_ (.A(net200),
    .B(_04984_),
    .Y(_05014_));
 sky130_fd_sc_hd__o21ai_0 _15753_ (.A1(_04984_),
    .A2(_05012_),
    .B1(_05014_),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_1 _15754_ (.A(_13168_),
    .Y(_05015_));
 sky130_fd_sc_hd__o21ai_2 _15755_ (.A1(_13164_),
    .A2(_05001_),
    .B1(_13169_),
    .Y(_05016_));
 sky130_fd_sc_hd__a21boi_4 _15756_ (.A1(_05015_),
    .A2(_05016_),
    .B1_N(_13173_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _15757_ (.A(_05015_),
    .B(_05016_),
    .Y(_05018_));
 sky130_fd_sc_hd__nor2_1 _15758_ (.A(_13173_),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__nand2_1 _15759_ (.A(\w[62][5] ),
    .B(net531),
    .Y(_05020_));
 sky130_fd_sc_hd__o31a_4 _15760_ (.A1(net531),
    .A2(_05017_),
    .A3(_05019_),
    .B1(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1374 ();
 sky130_fd_sc_hd__nand2_1 _15762_ (.A(net189),
    .B(_04984_),
    .Y(_05023_));
 sky130_fd_sc_hd__o21ai_0 _15763_ (.A1(_04984_),
    .A2(_05021_),
    .B1(_05023_),
    .Y(_00156_));
 sky130_fd_sc_hd__o21ai_0 _15764_ (.A1(_05007_),
    .A2(_05009_),
    .B1(_05015_),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_1 _15765_ (.A(_13173_),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__nor2_1 _15766_ (.A(_13177_),
    .B(_13172_),
    .Y(_05026_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_13168_),
    .B(_13172_),
    .Y(_05027_));
 sky130_fd_sc_hd__o21ai_2 _15768_ (.A1(_05007_),
    .A2(_05009_),
    .B1(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__o21a_1 _15769_ (.A1(_13173_),
    .A2(_13172_),
    .B1(_13177_),
    .X(_05029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1373 ();
 sky130_fd_sc_hd__a221oi_4 _15771_ (.A1(_05025_),
    .A2(_05026_),
    .B1(_05028_),
    .B2(_05029_),
    .C1(net530),
    .Y(_05031_));
 sky130_fd_sc_hd__a21oi_4 _15772_ (.A1(\w[62][6] ),
    .A2(net531),
    .B1(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1372 ();
 sky130_fd_sc_hd__nand2_1 _15774_ (.A(net178),
    .B(_04984_),
    .Y(_05034_));
 sky130_fd_sc_hd__o21ai_0 _15775_ (.A1(_04984_),
    .A2(_05032_),
    .B1(_05034_),
    .Y(_00157_));
 sky130_fd_sc_hd__o21ai_2 _15776_ (.A1(_13172_),
    .A2(_05017_),
    .B1(_13177_),
    .Y(_05035_));
 sky130_fd_sc_hd__nand2b_2 _15777_ (.A_N(_13176_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__xnor2_4 _15778_ (.A(_13181_),
    .B(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nor2_1 _15779_ (.A(net527),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__a21oi_4 _15780_ (.A1(\w[62][7] ),
    .A2(net527),
    .B1(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1371 ();
 sky130_fd_sc_hd__nand2_1 _15782_ (.A(net167),
    .B(_04984_),
    .Y(_05041_));
 sky130_fd_sc_hd__o21ai_0 _15783_ (.A1(_04984_),
    .A2(_05039_),
    .B1(_05041_),
    .Y(_00158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1370 ();
 sky130_fd_sc_hd__clkinvlp_4 _15785_ (.A(_13185_),
    .Y(_05043_));
 sky130_fd_sc_hd__a21o_2 _15786_ (.A1(_05028_),
    .A2(_05029_),
    .B1(_13176_),
    .X(_05044_));
 sky130_fd_sc_hd__a21oi_4 _15787_ (.A1(_13181_),
    .A2(_05044_),
    .B1(_13180_),
    .Y(_05045_));
 sky130_fd_sc_hd__xnor2_4 _15788_ (.A(_05043_),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__nor2_1 _15789_ (.A(net527),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__a21oi_4 _15790_ (.A1(\w[62][8] ),
    .A2(net527),
    .B1(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1369 ();
 sky130_fd_sc_hd__nand2_1 _15792_ (.A(net156),
    .B(_04984_),
    .Y(_05050_));
 sky130_fd_sc_hd__o21ai_0 _15793_ (.A1(_04984_),
    .A2(_05048_),
    .B1(_05050_),
    .Y(_00159_));
 sky130_fd_sc_hd__a21oi_1 _15794_ (.A1(_13181_),
    .A2(_05036_),
    .B1(_13180_),
    .Y(_05051_));
 sky130_fd_sc_hd__o21bai_2 _15795_ (.A1(_05043_),
    .A2(_05051_),
    .B1_N(_13184_),
    .Y(_05052_));
 sky130_fd_sc_hd__xnor2_4 _15796_ (.A(_13189_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__nor2_1 _15797_ (.A(net538),
    .B(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__a21oi_4 _15798_ (.A1(\w[62][9] ),
    .A2(net538),
    .B1(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1368 ();
 sky130_fd_sc_hd__nand2_1 _15800_ (.A(net145),
    .B(_04984_),
    .Y(_05057_));
 sky130_fd_sc_hd__o21ai_0 _15801_ (.A1(_04984_),
    .A2(_05055_),
    .B1(_05057_),
    .Y(_00160_));
 sky130_fd_sc_hd__o21bai_1 _15802_ (.A1(_05043_),
    .A2(_05045_),
    .B1_N(_13184_),
    .Y(_05058_));
 sky130_fd_sc_hd__a21oi_1 _15803_ (.A1(_13189_),
    .A2(_05058_),
    .B1(_13188_),
    .Y(_05059_));
 sky130_fd_sc_hd__xor2_2 _15804_ (.A(_13193_),
    .B(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__nor2_1 _15805_ (.A(net528),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__a21oi_4 _15806_ (.A1(\w[62][10] ),
    .A2(net528),
    .B1(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1366 ();
 sky130_fd_sc_hd__nand2_1 _15809_ (.A(net134),
    .B(_04984_),
    .Y(_05065_));
 sky130_fd_sc_hd__o21ai_0 _15810_ (.A1(_04984_),
    .A2(_05062_),
    .B1(_05065_),
    .Y(_00130_));
 sky130_fd_sc_hd__a21o_1 _15811_ (.A1(_13189_),
    .A2(_13184_),
    .B1(_13188_),
    .X(_05066_));
 sky130_fd_sc_hd__a21oi_1 _15812_ (.A1(_13193_),
    .A2(_05066_),
    .B1(_13192_),
    .Y(_05067_));
 sky130_fd_sc_hd__nor2b_2 _15813_ (.A(_05067_),
    .B_N(_13197_),
    .Y(_05068_));
 sky130_fd_sc_hd__and4_1 _15814_ (.A(_13185_),
    .B(_13189_),
    .C(_13193_),
    .D(_13197_),
    .X(_05069_));
 sky130_fd_sc_hd__o21a_1 _15815_ (.A1(_13181_),
    .A2(_13180_),
    .B1(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__nor2_1 _15816_ (.A(_05068_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__nor3_2 _15817_ (.A(_13180_),
    .B(_05036_),
    .C(_05068_),
    .Y(_05072_));
 sky130_fd_sc_hd__nor2_2 _15818_ (.A(_05071_),
    .B(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__a21o_1 _15819_ (.A1(_13189_),
    .A2(_05052_),
    .B1(_13188_),
    .X(_05074_));
 sky130_fd_sc_hd__a211oi_4 _15820_ (.A1(_13193_),
    .A2(_05074_),
    .B1(_13192_),
    .C1(_13197_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand2_1 _15821_ (.A(\w[62][11] ),
    .B(net528),
    .Y(_05076_));
 sky130_fd_sc_hd__o31a_4 _15822_ (.A1(net528),
    .A2(_05073_),
    .A3(_05075_),
    .B1(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1365 ();
 sky130_fd_sc_hd__nand2_1 _15824_ (.A(net123),
    .B(_04984_),
    .Y(_05079_));
 sky130_fd_sc_hd__o21ai_0 _15825_ (.A1(_04984_),
    .A2(_05077_),
    .B1(_05079_),
    .Y(_00131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1363 ();
 sky130_fd_sc_hd__inv_1 _15828_ (.A(_13201_),
    .Y(_05082_));
 sky130_fd_sc_hd__a211o_1 _15829_ (.A1(_13180_),
    .A2(_05069_),
    .B1(_05068_),
    .C1(_13196_),
    .X(_05083_));
 sky130_fd_sc_hd__a31oi_4 _15830_ (.A1(_13181_),
    .A2(_05044_),
    .A3(_05069_),
    .B1(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__xnor2_1 _15831_ (.A(_05082_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__nor2_1 _15832_ (.A(net530),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__a21oi_4 _15833_ (.A1(\w[62][12] ),
    .A2(net530),
    .B1(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1362 ();
 sky130_fd_sc_hd__nand2_1 _15835_ (.A(net111),
    .B(_04984_),
    .Y(_05089_));
 sky130_fd_sc_hd__o21ai_0 _15836_ (.A1(_04984_),
    .A2(_05087_),
    .B1(_05089_),
    .Y(_00132_));
 sky130_fd_sc_hd__clkinvlp_4 _15837_ (.A(_13205_),
    .Y(_05090_));
 sky130_fd_sc_hd__o21a_1 _15838_ (.A1(_13196_),
    .A2(_05073_),
    .B1(_13201_),
    .X(_05091_));
 sky130_fd_sc_hd__nor2_1 _15839_ (.A(_13200_),
    .B(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__xnor2_4 _15840_ (.A(_05090_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__nor2_1 _15841_ (.A(net527),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__a21oi_4 _15842_ (.A1(\w[62][13] ),
    .A2(net527),
    .B1(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1361 ();
 sky130_fd_sc_hd__nand2_1 _15844_ (.A(net100),
    .B(_04984_),
    .Y(_05097_));
 sky130_fd_sc_hd__o21ai_0 _15845_ (.A1(_04984_),
    .A2(_05095_),
    .B1(_05097_),
    .Y(_00133_));
 sky130_fd_sc_hd__o21bai_1 _15846_ (.A1(_05082_),
    .A2(_05084_),
    .B1_N(_13200_),
    .Y(_05098_));
 sky130_fd_sc_hd__a21oi_1 _15847_ (.A1(_13205_),
    .A2(_05098_),
    .B1(_13204_),
    .Y(_05099_));
 sky130_fd_sc_hd__xor2_1 _15848_ (.A(_13209_),
    .B(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__nor2_2 _15849_ (.A(net538),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__a21oi_4 _15850_ (.A1(\w[62][14] ),
    .A2(net538),
    .B1(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1360 ();
 sky130_fd_sc_hd__nand2_1 _15852_ (.A(net89),
    .B(_04984_),
    .Y(_05104_));
 sky130_fd_sc_hd__o21ai_0 _15853_ (.A1(_04984_),
    .A2(_05102_),
    .B1(_05104_),
    .Y(_00134_));
 sky130_fd_sc_hd__nand3_2 _15854_ (.A(_13201_),
    .B(_13205_),
    .C(_13209_),
    .Y(_05105_));
 sky130_fd_sc_hd__a21oi_1 _15855_ (.A1(_13201_),
    .A2(_13196_),
    .B1(_13200_),
    .Y(_05106_));
 sky130_fd_sc_hd__o21bai_1 _15856_ (.A1(_05090_),
    .A2(_05106_),
    .B1_N(_13204_),
    .Y(_05107_));
 sky130_fd_sc_hd__a21oi_2 _15857_ (.A1(_13209_),
    .A2(_05107_),
    .B1(_13208_),
    .Y(_05108_));
 sky130_fd_sc_hd__o31ai_4 _15858_ (.A1(_05071_),
    .A2(_05072_),
    .A3(_05105_),
    .B1(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__xnor2_2 _15859_ (.A(_13213_),
    .B(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__nor2_2 _15860_ (.A(net538),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__a21oi_4 _15861_ (.A1(\w[62][15] ),
    .A2(net531),
    .B1(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1359 ();
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(net78),
    .B(_04984_),
    .Y(_05114_));
 sky130_fd_sc_hd__o21ai_0 _15864_ (.A1(_04984_),
    .A2(_05112_),
    .B1(_05114_),
    .Y(_00135_));
 sky130_fd_sc_hd__a21o_1 _15865_ (.A1(_13205_),
    .A2(_13200_),
    .B1(_13204_),
    .X(_05115_));
 sky130_fd_sc_hd__a21oi_1 _15866_ (.A1(_13209_),
    .A2(_05115_),
    .B1(_13208_),
    .Y(_05116_));
 sky130_fd_sc_hd__o21ai_0 _15867_ (.A1(_05084_),
    .A2(_05105_),
    .B1(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__a21oi_2 _15868_ (.A1(_13213_),
    .A2(_05117_),
    .B1(_13212_),
    .Y(_05118_));
 sky130_fd_sc_hd__xor2_4 _15869_ (.A(_13217_),
    .B(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__nor2_1 _15870_ (.A(net529),
    .B(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__a21oi_4 _15871_ (.A1(\w[62][16] ),
    .A2(net529),
    .B1(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1358 ();
 sky130_fd_sc_hd__nand2_1 _15873_ (.A(net67),
    .B(_04984_),
    .Y(_05123_));
 sky130_fd_sc_hd__o21ai_0 _15874_ (.A1(_04984_),
    .A2(_05121_),
    .B1(_05123_),
    .Y(_00136_));
 sky130_fd_sc_hd__a21o_1 _15875_ (.A1(_13213_),
    .A2(_05109_),
    .B1(_13212_),
    .X(_05124_));
 sky130_fd_sc_hd__a21oi_2 _15876_ (.A1(_13217_),
    .A2(_05124_),
    .B1(_13216_),
    .Y(_05125_));
 sky130_fd_sc_hd__xor2_4 _15877_ (.A(_13221_),
    .B(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__nor2_1 _15878_ (.A(net528),
    .B(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__a21oi_4 _15879_ (.A1(\w[62][17] ),
    .A2(net528),
    .B1(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1357 ();
 sky130_fd_sc_hd__nand2_1 _15881_ (.A(net56),
    .B(_04984_),
    .Y(_05130_));
 sky130_fd_sc_hd__o21ai_0 _15882_ (.A1(_04984_),
    .A2(_05128_),
    .B1(_05130_),
    .Y(_00137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1356 ();
 sky130_fd_sc_hd__nand2_1 _15884_ (.A(_13217_),
    .B(_13221_),
    .Y(_05132_));
 sky130_fd_sc_hd__a21oi_1 _15885_ (.A1(_13221_),
    .A2(_13216_),
    .B1(_13220_),
    .Y(_05133_));
 sky130_fd_sc_hd__o21ai_0 _15886_ (.A1(_05118_),
    .A2(_05132_),
    .B1(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__xnor2_1 _15887_ (.A(_13225_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__nor2_2 _15888_ (.A(net530),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__a21oi_4 _15889_ (.A1(\w[62][18] ),
    .A2(net538),
    .B1(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1355 ();
 sky130_fd_sc_hd__nand2_1 _15891_ (.A(net45),
    .B(_04984_),
    .Y(_05139_));
 sky130_fd_sc_hd__o21ai_0 _15892_ (.A1(_04984_),
    .A2(_05137_),
    .B1(_05139_),
    .Y(_00138_));
 sky130_fd_sc_hd__nor3_1 _15893_ (.A(_13176_),
    .B(_13180_),
    .C(_05068_),
    .Y(_05140_));
 sky130_fd_sc_hd__nand2_1 _15894_ (.A(_13213_),
    .B(_13225_),
    .Y(_05141_));
 sky130_fd_sc_hd__nor3_1 _15895_ (.A(_05105_),
    .B(_05132_),
    .C(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21ai_0 _15896_ (.A1(_05068_),
    .A2(_05070_),
    .B1(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__a21oi_2 _15897_ (.A1(_05035_),
    .A2(_05140_),
    .B1(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__nand2_1 _15898_ (.A(_13213_),
    .B(_13217_),
    .Y(_05145_));
 sky130_fd_sc_hd__a21oi_1 _15899_ (.A1(_13217_),
    .A2(_13212_),
    .B1(_13216_),
    .Y(_05146_));
 sky130_fd_sc_hd__o21a_1 _15900_ (.A1(_05108_),
    .A2(_05145_),
    .B1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__nand2_1 _15901_ (.A(_13221_),
    .B(_13225_),
    .Y(_05148_));
 sky130_fd_sc_hd__a21oi_1 _15902_ (.A1(_13225_),
    .A2(_13220_),
    .B1(_13224_),
    .Y(_05149_));
 sky130_fd_sc_hd__o21ai_2 _15903_ (.A1(_05147_),
    .A2(_05148_),
    .B1(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__or2_0 _15904_ (.A(_05144_),
    .B(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__xnor2_2 _15905_ (.A(_13229_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__nor2_4 _15906_ (.A(net530),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21oi_4 _15907_ (.A1(\w[62][19] ),
    .A2(net531),
    .B1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1354 ();
 sky130_fd_sc_hd__nand2_1 _15909_ (.A(net34),
    .B(_04984_),
    .Y(_05156_));
 sky130_fd_sc_hd__o21ai_0 _15910_ (.A1(_04984_),
    .A2(_05154_),
    .B1(_05156_),
    .Y(_00139_));
 sky130_fd_sc_hd__nor4b_1 _15911_ (.A(_13212_),
    .B(_13224_),
    .C(_13228_),
    .D_N(_05133_),
    .Y(_05157_));
 sky130_fd_sc_hd__and2_0 _15912_ (.A(_05116_),
    .B(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__nand2_1 _15913_ (.A(_05105_),
    .B(_05116_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2_1 _15914_ (.A(_13213_),
    .B(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_1 _15915_ (.A(_05133_),
    .B(_05132_),
    .Y(_05161_));
 sky130_fd_sc_hd__a21o_1 _15916_ (.A1(_13225_),
    .A2(_05161_),
    .B1(_13224_),
    .X(_05162_));
 sky130_fd_sc_hd__a21oi_1 _15917_ (.A1(_13229_),
    .A2(_05162_),
    .B1(_13228_),
    .Y(_05163_));
 sky130_fd_sc_hd__a21o_1 _15918_ (.A1(_05157_),
    .A2(_05160_),
    .B1(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__a21oi_2 _15919_ (.A1(_05084_),
    .A2(_05158_),
    .B1(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__xor2_4 _15920_ (.A(_13233_),
    .B(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__mux2i_4 _15921_ (.A0(_05166_),
    .A1(\w[62][20] ),
    .S(net527),
    .Y(_05167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1352 ();
 sky130_fd_sc_hd__nand2_1 _15924_ (.A(net23),
    .B(_04984_),
    .Y(_05170_));
 sky130_fd_sc_hd__o21ai_0 _15925_ (.A1(_04984_),
    .A2(_05167_),
    .B1(_05170_),
    .Y(_00141_));
 sky130_fd_sc_hd__a21o_1 _15926_ (.A1(_13233_),
    .A2(_13228_),
    .B1(_13232_),
    .X(_05171_));
 sky130_fd_sc_hd__a31oi_1 _15927_ (.A1(_13229_),
    .A2(_13233_),
    .A3(_05151_),
    .B1(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__xor2_1 _15928_ (.A(_13237_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__nor2_1 _15929_ (.A(net530),
    .B(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__a21oi_4 _15930_ (.A1(\w[62][21] ),
    .A2(net530),
    .B1(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1351 ();
 sky130_fd_sc_hd__nand2_1 _15932_ (.A(net12),
    .B(_04984_),
    .Y(_05177_));
 sky130_fd_sc_hd__o21ai_0 _15933_ (.A1(_04984_),
    .A2(_05175_),
    .B1(_05177_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _15934_ (.A(_13233_),
    .B(_13237_),
    .Y(_05178_));
 sky130_fd_sc_hd__a211oi_2 _15935_ (.A1(_05084_),
    .A2(_05158_),
    .B1(_05164_),
    .C1(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__a21o_1 _15936_ (.A1(_13237_),
    .A2(_13232_),
    .B1(_13236_),
    .X(_05180_));
 sky130_fd_sc_hd__nor2_1 _15937_ (.A(_05179_),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__xor2_2 _15938_ (.A(_13241_),
    .B(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__nor2_1 _15939_ (.A(net530),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21oi_4 _15940_ (.A1(\w[62][22] ),
    .A2(net530),
    .B1(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1350 ();
 sky130_fd_sc_hd__nand2_1 _15942_ (.A(net761),
    .B(_04984_),
    .Y(_05186_));
 sky130_fd_sc_hd__o21ai_0 _15943_ (.A1(_04984_),
    .A2(_05184_),
    .B1(_05186_),
    .Y(_00143_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1348 ();
 sky130_fd_sc_hd__and2_0 _15946_ (.A(_13237_),
    .B(_13241_),
    .X(_05189_));
 sky130_fd_sc_hd__o2111ai_4 _15947_ (.A1(_05144_),
    .A2(_05150_),
    .B1(_05189_),
    .C1(_13233_),
    .D1(_13229_),
    .Y(_05190_));
 sky130_fd_sc_hd__a21o_1 _15948_ (.A1(_13237_),
    .A2(_05171_),
    .B1(_13236_),
    .X(_05191_));
 sky130_fd_sc_hd__a21oi_1 _15949_ (.A1(_13241_),
    .A2(_05191_),
    .B1(_13240_),
    .Y(_05192_));
 sky130_fd_sc_hd__nand2_1 _15950_ (.A(_05190_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__xnor2_1 _15951_ (.A(_13245_),
    .B(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__nor2_2 _15952_ (.A(net529),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__a21oi_4 _15953_ (.A1(\w[62][23] ),
    .A2(net538),
    .B1(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1347 ();
 sky130_fd_sc_hd__nand2_1 _15955_ (.A(net750),
    .B(_04984_),
    .Y(_05198_));
 sky130_fd_sc_hd__o21ai_0 _15956_ (.A1(_04984_),
    .A2(_05196_),
    .B1(_05198_),
    .Y(_00144_));
 sky130_fd_sc_hd__clkinvlp_4 _15957_ (.A(_13249_),
    .Y(_05199_));
 sky130_fd_sc_hd__nor3_1 _15958_ (.A(_13241_),
    .B(_13240_),
    .C(_13244_),
    .Y(_05200_));
 sky130_fd_sc_hd__nor2_1 _15959_ (.A(_13245_),
    .B(_13244_),
    .Y(_05201_));
 sky130_fd_sc_hd__nor2_1 _15960_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__o41ai_4 _15961_ (.A1(_13240_),
    .A2(_13244_),
    .A3(_05179_),
    .A4(_05180_),
    .B1(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__xnor2_4 _15962_ (.A(_05199_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__nor2_1 _15963_ (.A(net527),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__a21oi_4 _15964_ (.A1(\w[62][24] ),
    .A2(net527),
    .B1(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1346 ();
 sky130_fd_sc_hd__nand2_1 _15966_ (.A(net739),
    .B(_04984_),
    .Y(_05208_));
 sky130_fd_sc_hd__o21ai_0 _15967_ (.A1(_04984_),
    .A2(_05206_),
    .B1(_05208_),
    .Y(_00145_));
 sky130_fd_sc_hd__nor3b_1 _15968_ (.A(_13244_),
    .B(_13248_),
    .C_N(_05192_),
    .Y(_05209_));
 sky130_fd_sc_hd__o21ba_1 _15969_ (.A1(_05199_),
    .A2(_05201_),
    .B1_N(_13248_),
    .X(_05210_));
 sky130_fd_sc_hd__a21oi_1 _15970_ (.A1(_05190_),
    .A2(_05209_),
    .B1(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__xnor2_1 _15971_ (.A(_13253_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nor2_1 _15972_ (.A(net528),
    .B(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__a21oi_4 _15973_ (.A1(\w[62][25] ),
    .A2(net528),
    .B1(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1345 ();
 sky130_fd_sc_hd__nand2_1 _15975_ (.A(net728),
    .B(_04984_),
    .Y(_05216_));
 sky130_fd_sc_hd__o21ai_0 _15976_ (.A1(_04984_),
    .A2(_05214_),
    .B1(_05216_),
    .Y(_00146_));
 sky130_fd_sc_hd__o21bai_1 _15977_ (.A1(_05199_),
    .A2(_05203_),
    .B1_N(_13248_),
    .Y(_05217_));
 sky130_fd_sc_hd__a211o_1 _15978_ (.A1(_13253_),
    .A2(_05217_),
    .B1(_13252_),
    .C1(_13257_),
    .X(_05218_));
 sky130_fd_sc_hd__nand3_1 _15979_ (.A(_13249_),
    .B(_13253_),
    .C(_13257_),
    .Y(_05219_));
 sky130_fd_sc_hd__and3_1 _15980_ (.A(_13253_),
    .B(_13257_),
    .C(_13248_),
    .X(_05220_));
 sky130_fd_sc_hd__a21oi_1 _15981_ (.A1(_13257_),
    .A2(_13252_),
    .B1(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__o21ai_1 _15982_ (.A1(_05203_),
    .A2(_05219_),
    .B1(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__nor2_1 _15983_ (.A(net529),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__a22oi_4 _15984_ (.A1(\w[62][26] ),
    .A2(net529),
    .B1(_05218_),
    .B2(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1344 ();
 sky130_fd_sc_hd__nand2_1 _15986_ (.A(net717),
    .B(_04984_),
    .Y(_05226_));
 sky130_fd_sc_hd__o21ai_0 _15987_ (.A1(_04984_),
    .A2(_05224_),
    .B1(_05226_),
    .Y(_00147_));
 sky130_fd_sc_hd__and2_0 _15988_ (.A(_13253_),
    .B(_05211_),
    .X(_05227_));
 sky130_fd_sc_hd__o21ai_1 _15989_ (.A1(_13252_),
    .A2(_05227_),
    .B1(_13257_),
    .Y(_05228_));
 sky130_fd_sc_hd__nor2_1 _15990_ (.A(_13261_),
    .B(_13256_),
    .Y(_05229_));
 sky130_fd_sc_hd__nand3_1 _15991_ (.A(_13253_),
    .B(_13257_),
    .C(_13261_),
    .Y(_05230_));
 sky130_fd_sc_hd__a211oi_4 _15992_ (.A1(_05190_),
    .A2(_05209_),
    .B1(_05210_),
    .C1(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand2_1 _15993_ (.A(_13261_),
    .B(_13256_),
    .Y(_05232_));
 sky130_fd_sc_hd__nand3_1 _15994_ (.A(_13257_),
    .B(_13261_),
    .C(_13252_),
    .Y(_05233_));
 sky130_fd_sc_hd__nand2_1 _15995_ (.A(_05232_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__a2111oi_4 _15996_ (.A1(_05228_),
    .A2(_05229_),
    .B1(_05231_),
    .C1(_05234_),
    .D1(net529),
    .Y(_05235_));
 sky130_fd_sc_hd__a21oi_4 _15997_ (.A1(\w[62][27] ),
    .A2(net528),
    .B1(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1343 ();
 sky130_fd_sc_hd__nand2_1 _15999_ (.A(net445),
    .B(_04984_),
    .Y(_05238_));
 sky130_fd_sc_hd__o21ai_0 _16000_ (.A1(_04984_),
    .A2(_05236_),
    .B1(_05238_),
    .Y(_00148_));
 sky130_fd_sc_hd__o21a_1 _16001_ (.A1(_13256_),
    .A2(_05222_),
    .B1(_13261_),
    .X(_05239_));
 sky130_fd_sc_hd__nor2_1 _16002_ (.A(_13260_),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__xnor2_4 _16003_ (.A(_13265_),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1342 ();
 sky130_fd_sc_hd__mux2i_4 _16005_ (.A0(_05241_),
    .A1(\w[62][28] ),
    .S(net527),
    .Y(_05243_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1341 ();
 sky130_fd_sc_hd__nand2_1 _16007_ (.A(net334),
    .B(_04984_),
    .Y(_05245_));
 sky130_fd_sc_hd__o21ai_0 _16008_ (.A1(_04984_),
    .A2(_05243_),
    .B1(_05245_),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_1 _16009_ (.A(_13269_),
    .Y(_05246_));
 sky130_fd_sc_hd__or3_1 _16010_ (.A(_13260_),
    .B(_05231_),
    .C(_05234_),
    .X(_05247_));
 sky130_fd_sc_hd__a21oi_1 _16011_ (.A1(_13265_),
    .A2(_05247_),
    .B1(_13264_),
    .Y(_05248_));
 sky130_fd_sc_hd__xnor2_1 _16012_ (.A(_05246_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__nor2_1 _16013_ (.A(net529),
    .B(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__a21oi_4 _16014_ (.A1(\w[62][29] ),
    .A2(net529),
    .B1(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1340 ();
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(net223),
    .B(_04984_),
    .Y(_05253_));
 sky130_fd_sc_hd__o21ai_0 _16017_ (.A1(_04984_),
    .A2(_05251_),
    .B1(_05253_),
    .Y(_00150_));
 sky130_fd_sc_hd__or4_1 _16018_ (.A(_13256_),
    .B(_13260_),
    .C(_13264_),
    .D(_05222_),
    .X(_05254_));
 sky130_fd_sc_hd__nor3_1 _16019_ (.A(_13261_),
    .B(_13260_),
    .C(_13264_),
    .Y(_05255_));
 sky130_fd_sc_hd__nor2_1 _16020_ (.A(_13265_),
    .B(_13264_),
    .Y(_05256_));
 sky130_fd_sc_hd__nor2_1 _16021_ (.A(_05255_),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__a31oi_4 _16022_ (.A1(_13269_),
    .A2(_05254_),
    .A3(_05257_),
    .B1(_13268_),
    .Y(_05258_));
 sky130_fd_sc_hd__xnor2_4 _16023_ (.A(_13273_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__mux2i_4 _16024_ (.A0(_05259_),
    .A1(\w[62][30] ),
    .S(net531),
    .Y(_05260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1339 ();
 sky130_fd_sc_hd__nand2_1 _16026_ (.A(net112),
    .B(_04984_),
    .Y(_05262_));
 sky130_fd_sc_hd__o21ai_0 _16027_ (.A1(_04984_),
    .A2(_05260_),
    .B1(_05262_),
    .Y(_00152_));
 sky130_fd_sc_hd__xor2_1 _16028_ (.A(_11993_),
    .B(_11996_),
    .X(_05263_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1335 ();
 sky130_fd_sc_hd__mux4_1 _16033_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net585),
    .S1(net589),
    .X(_05268_));
 sky130_fd_sc_hd__mux4_1 _16034_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net585),
    .S1(net589),
    .X(_05269_));
 sky130_fd_sc_hd__mux4_1 _16035_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net585),
    .S1(net589),
    .X(_05270_));
 sky130_fd_sc_hd__mux4_1 _16036_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net585),
    .S1(net589),
    .X(_05271_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1334 ();
 sky130_fd_sc_hd__mux4_4 _16038_ (.A0(_05268_),
    .A1(_05269_),
    .A2(_05270_),
    .A3(_05271_),
    .S0(net578),
    .S1(net576),
    .X(_05273_));
 sky130_fd_sc_hd__mux4_1 _16039_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net585),
    .S1(net587),
    .X(_05274_));
 sky130_fd_sc_hd__mux4_1 _16040_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net585),
    .S1(net587),
    .X(_05275_));
 sky130_fd_sc_hd__mux4_1 _16041_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net585),
    .S1(net587),
    .X(_05276_));
 sky130_fd_sc_hd__mux4_1 _16042_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net585),
    .S1(net587),
    .X(_05277_));
 sky130_fd_sc_hd__mux4_1 _16043_ (.A0(_05274_),
    .A1(_05275_),
    .A2(_05276_),
    .A3(_05277_),
    .S0(net578),
    .S1(net576),
    .X(_05278_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1333 ();
 sky130_fd_sc_hd__mux2i_4 _16045_ (.A0(_05273_),
    .A1(_05278_),
    .S(net574),
    .Y(_05280_));
 sky130_fd_sc_hd__xnor2_1 _16046_ (.A(_05263_),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1329 ();
 sky130_fd_sc_hd__mux4_1 _16051_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05286_));
 sky130_fd_sc_hd__mux4_1 _16052_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05287_));
 sky130_fd_sc_hd__mux4_1 _16053_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05288_));
 sky130_fd_sc_hd__mux4_1 _16054_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05289_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1328 ();
 sky130_fd_sc_hd__mux4_4 _16056_ (.A0(_05286_),
    .A1(_05287_),
    .A2(_05288_),
    .A3(_05289_),
    .S0(net653),
    .S1(net651),
    .X(_05291_));
 sky130_fd_sc_hd__mux4_1 _16057_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05292_));
 sky130_fd_sc_hd__mux4_1 _16058_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05293_));
 sky130_fd_sc_hd__mux4_1 _16059_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05294_));
 sky130_fd_sc_hd__mux4_1 _16060_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net654),
    .S1(net661),
    .X(_05295_));
 sky130_fd_sc_hd__mux4_1 _16061_ (.A0(_05292_),
    .A1(_05293_),
    .A2(_05294_),
    .A3(_05295_),
    .S0(net653),
    .S1(net651),
    .X(_05296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1327 ();
 sky130_fd_sc_hd__mux2i_4 _16063_ (.A0(_05291_),
    .A1(_05296_),
    .S(net648),
    .Y(_05298_));
 sky130_fd_sc_hd__xor2_1 _16064_ (.A(_02595_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__xnor2_1 _16065_ (.A(_05281_),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__xor2_1 _16066_ (.A(_11457_),
    .B(_11632_),
    .X(_05301_));
 sky130_fd_sc_hd__xnor2_1 _16067_ (.A(_11349_),
    .B(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__xnor2_2 _16068_ (.A(_05300_),
    .B(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__nor2_1 _16069_ (.A(_05231_),
    .B(_05234_),
    .Y(_05304_));
 sky130_fd_sc_hd__nor3_1 _16070_ (.A(_13260_),
    .B(_13264_),
    .C(_13268_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(_05304_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__o21bai_1 _16072_ (.A1(_05246_),
    .A2(_05256_),
    .B1_N(_13268_),
    .Y(_05307_));
 sky130_fd_sc_hd__a31oi_4 _16073_ (.A1(_13273_),
    .A2(_05306_),
    .A3(_05307_),
    .B1(_13272_),
    .Y(_05308_));
 sky130_fd_sc_hd__xnor2_4 _16074_ (.A(_05303_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__mux2i_4 _16075_ (.A0(_05309_),
    .A1(\w[62][31] ),
    .S(net528),
    .Y(_05310_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1326 ();
 sky130_fd_sc_hd__nand2_1 _16077_ (.A(net1),
    .B(_04984_),
    .Y(_05312_));
 sky130_fd_sc_hd__o21ai_0 _16078_ (.A1(_04984_),
    .A2(_05310_),
    .B1(_05312_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2b_4 _16079_ (.A(net762),
    .B_N(_13704_),
    .Y(_05313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1325 ();
 sky130_fd_sc_hd__nand2_8 _16081_ (.A(_09959_),
    .B(_05313_),
    .Y(_05315_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1324 ();
 sky130_fd_sc_hd__mux2i_4 _16083_ (.A0(_13277_),
    .A1(\w[63][0] ),
    .S(done),
    .Y(_05317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1322 ();
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(net721),
    .B(_05315_),
    .Y(_05320_));
 sky130_fd_sc_hd__o21ai_0 _16087_ (.A1(_05315_),
    .A2(_05317_),
    .B1(_05320_),
    .Y(_00353_));
 sky130_fd_sc_hd__mux2i_4 _16088_ (.A0(_13280_),
    .A1(\w[63][1] ),
    .S(done),
    .Y(_05321_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1321 ();
 sky130_fd_sc_hd__nand2_1 _16090_ (.A(net720),
    .B(_05315_),
    .Y(_05323_));
 sky130_fd_sc_hd__o21ai_0 _16091_ (.A1(_05315_),
    .A2(_05321_),
    .B1(_05323_),
    .Y(_00364_));
 sky130_fd_sc_hd__mux2i_4 _16092_ (.A0(_12021_),
    .A1(\w[63][2] ),
    .S(net537),
    .Y(_05324_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1320 ();
 sky130_fd_sc_hd__nand2_1 _16094_ (.A(net719),
    .B(_05315_),
    .Y(_05326_));
 sky130_fd_sc_hd__o21ai_0 _16095_ (.A1(_05315_),
    .A2(_05324_),
    .B1(_05326_),
    .Y(_00375_));
 sky130_fd_sc_hd__nor2b_1 _16096_ (.A(_13288_),
    .B_N(_12020_),
    .Y(_05327_));
 sky130_fd_sc_hd__nor2b_1 _16097_ (.A(_12020_),
    .B_N(_13288_),
    .Y(_05328_));
 sky130_fd_sc_hd__nor3_1 _16098_ (.A(net537),
    .B(_05327_),
    .C(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__a21oi_4 _16099_ (.A1(\w[63][3] ),
    .A2(net537),
    .B1(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1319 ();
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(net718),
    .B(_05315_),
    .Y(_05332_));
 sky130_fd_sc_hd__o21ai_0 _16102_ (.A1(_05315_),
    .A2(_05330_),
    .B1(_05332_),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_1 _16103_ (.A(_13292_),
    .Y(_05333_));
 sky130_fd_sc_hd__a21o_1 _16104_ (.A1(_13279_),
    .A2(_13284_),
    .B1(_13283_),
    .X(_05334_));
 sky130_fd_sc_hd__a21oi_1 _16105_ (.A1(_13288_),
    .A2(_05334_),
    .B1(_13287_),
    .Y(_05335_));
 sky130_fd_sc_hd__xnor2_1 _16106_ (.A(_05333_),
    .B(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__nor2_2 _16107_ (.A(net537),
    .B(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__a21oi_4 _16108_ (.A1(\w[63][4] ),
    .A2(done),
    .B1(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1318 ();
 sky130_fd_sc_hd__nand2_1 _16110_ (.A(net716),
    .B(_05315_),
    .Y(_05340_));
 sky130_fd_sc_hd__o21ai_0 _16111_ (.A1(_05315_),
    .A2(_05338_),
    .B1(_05340_),
    .Y(_00379_));
 sky130_fd_sc_hd__inv_1 _16112_ (.A(_13291_),
    .Y(_05341_));
 sky130_fd_sc_hd__o21ai_0 _16113_ (.A1(_13287_),
    .A2(_05328_),
    .B1(_13292_),
    .Y(_05342_));
 sky130_fd_sc_hd__a21boi_1 _16114_ (.A1(_05341_),
    .A2(_05342_),
    .B1_N(_13296_),
    .Y(_05343_));
 sky130_fd_sc_hd__nand2_1 _16115_ (.A(_05341_),
    .B(_05342_),
    .Y(_05344_));
 sky130_fd_sc_hd__nor2_1 _16116_ (.A(_13296_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__nor3_2 _16117_ (.A(net537),
    .B(_05343_),
    .C(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__a21oi_4 _16118_ (.A1(\w[63][5] ),
    .A2(done),
    .B1(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1317 ();
 sky130_fd_sc_hd__nand2_1 _16120_ (.A(net715),
    .B(_05315_),
    .Y(_05349_));
 sky130_fd_sc_hd__o21ai_0 _16121_ (.A1(_05315_),
    .A2(_05347_),
    .B1(_05349_),
    .Y(_00380_));
 sky130_fd_sc_hd__nand2b_1 _16122_ (.A_N(_05335_),
    .B(_13292_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2_1 _16123_ (.A(_05341_),
    .B(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__a21oi_1 _16124_ (.A1(_13296_),
    .A2(_05351_),
    .B1(_13295_),
    .Y(_05352_));
 sky130_fd_sc_hd__xnor2_2 _16125_ (.A(_13300_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__mux2i_4 _16126_ (.A0(_05353_),
    .A1(\w[63][6] ),
    .S(net534),
    .Y(_05354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1316 ();
 sky130_fd_sc_hd__nand2_1 _16128_ (.A(net714),
    .B(_05315_),
    .Y(_05356_));
 sky130_fd_sc_hd__o21ai_0 _16129_ (.A1(_05315_),
    .A2(_05354_),
    .B1(_05356_),
    .Y(_00381_));
 sky130_fd_sc_hd__o21a_1 _16130_ (.A1(_13295_),
    .A2(_05343_),
    .B1(_13300_),
    .X(_05357_));
 sky130_fd_sc_hd__nor2_1 _16131_ (.A(_13299_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__xnor2_4 _16132_ (.A(_13304_),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__mux2i_4 _16133_ (.A0(_05359_),
    .A1(\w[63][7] ),
    .S(net532),
    .Y(_05360_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1315 ();
 sky130_fd_sc_hd__nand2_1 _16135_ (.A(net713),
    .B(_05315_),
    .Y(_05362_));
 sky130_fd_sc_hd__o21ai_0 _16136_ (.A1(_05315_),
    .A2(_05360_),
    .B1(_05362_),
    .Y(_00382_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1314 ();
 sky130_fd_sc_hd__nor3_1 _16138_ (.A(_13291_),
    .B(_13295_),
    .C(_13299_),
    .Y(_05364_));
 sky130_fd_sc_hd__o21a_1 _16139_ (.A1(_13296_),
    .A2(_13295_),
    .B1(_13300_),
    .X(_05365_));
 sky130_fd_sc_hd__o21ai_1 _16140_ (.A1(_13299_),
    .A2(_05365_),
    .B1(_13304_),
    .Y(_05366_));
 sky130_fd_sc_hd__a21oi_1 _16141_ (.A1(_05350_),
    .A2(_05364_),
    .B1(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__o21ai_0 _16142_ (.A1(_13303_),
    .A2(_05367_),
    .B1(_13308_),
    .Y(_05368_));
 sky130_fd_sc_hd__or3_1 _16143_ (.A(_13308_),
    .B(_13303_),
    .C(_05367_),
    .X(_05369_));
 sky130_fd_sc_hd__and3b_1 _16144_ (.A_N(net536),
    .B(_05368_),
    .C(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__a21oi_4 _16145_ (.A1(\w[63][8] ),
    .A2(net534),
    .B1(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1313 ();
 sky130_fd_sc_hd__nand2_1 _16147_ (.A(net712),
    .B(_05315_),
    .Y(_05373_));
 sky130_fd_sc_hd__o21ai_0 _16148_ (.A1(_05315_),
    .A2(_05371_),
    .B1(_05373_),
    .Y(_00383_));
 sky130_fd_sc_hd__inv_1 _16149_ (.A(_13303_),
    .Y(_05374_));
 sky130_fd_sc_hd__o21ai_2 _16150_ (.A1(_13299_),
    .A2(_05357_),
    .B1(_13304_),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_1 _16151_ (.A(_05374_),
    .B(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__a21oi_1 _16152_ (.A1(_13308_),
    .A2(_05376_),
    .B1(_13307_),
    .Y(_05377_));
 sky130_fd_sc_hd__xor2_1 _16153_ (.A(_13312_),
    .B(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__nor2_1 _16154_ (.A(net535),
    .B(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__a21oi_4 _16155_ (.A1(\w[63][9] ),
    .A2(net536),
    .B1(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1312 ();
 sky130_fd_sc_hd__nand2_1 _16157_ (.A(net711),
    .B(_05315_),
    .Y(_05382_));
 sky130_fd_sc_hd__o21ai_0 _16158_ (.A1(_05315_),
    .A2(_05380_),
    .B1(_05382_),
    .Y(_00384_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1311 ();
 sky130_fd_sc_hd__nand2b_1 _16160_ (.A_N(_13307_),
    .B(_05368_),
    .Y(_05384_));
 sky130_fd_sc_hd__a21oi_1 _16161_ (.A1(_13312_),
    .A2(_05384_),
    .B1(_13311_),
    .Y(_05385_));
 sky130_fd_sc_hd__xor2_2 _16162_ (.A(_13316_),
    .B(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__nor2_2 _16163_ (.A(net534),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__a21oi_4 _16164_ (.A1(\w[63][10] ),
    .A2(net535),
    .B1(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1309 ();
 sky130_fd_sc_hd__nand2_1 _16167_ (.A(net710),
    .B(_05315_),
    .Y(_05391_));
 sky130_fd_sc_hd__o21ai_0 _16168_ (.A1(_05315_),
    .A2(_05388_),
    .B1(_05391_),
    .Y(_00354_));
 sky130_fd_sc_hd__nor2b_1 _16169_ (.A(_05377_),
    .B_N(_13312_),
    .Y(_05392_));
 sky130_fd_sc_hd__o21ai_1 _16170_ (.A1(_13311_),
    .A2(_05392_),
    .B1(_13316_),
    .Y(_05393_));
 sky130_fd_sc_hd__nor2_1 _16171_ (.A(_13320_),
    .B(_13315_),
    .Y(_05394_));
 sky130_fd_sc_hd__a21oi_1 _16172_ (.A1(_13312_),
    .A2(_13307_),
    .B1(_13311_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_1 _16173_ (.A(_13316_),
    .B(_13320_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand2_1 _16174_ (.A(_13320_),
    .B(_13315_),
    .Y(_05397_));
 sky130_fd_sc_hd__o21ai_4 _16175_ (.A1(_05395_),
    .A2(_05396_),
    .B1(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__nand4_2 _16176_ (.A(_13308_),
    .B(_13312_),
    .C(_13316_),
    .D(_13320_),
    .Y(_05399_));
 sky130_fd_sc_hd__a21oi_4 _16177_ (.A1(_05374_),
    .A2(_05375_),
    .B1(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__a2111oi_4 _16178_ (.A1(_05393_),
    .A2(_05394_),
    .B1(net536),
    .C1(_05398_),
    .D1(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__a21oi_4 _16179_ (.A1(\w[63][11] ),
    .A2(net536),
    .B1(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1308 ();
 sky130_fd_sc_hd__nand2_1 _16181_ (.A(net709),
    .B(_05315_),
    .Y(_05404_));
 sky130_fd_sc_hd__o21ai_0 _16182_ (.A1(_05315_),
    .A2(_05402_),
    .B1(_05404_),
    .Y(_00355_));
 sky130_fd_sc_hd__inv_1 _16183_ (.A(_13324_),
    .Y(_05405_));
 sky130_fd_sc_hd__o21ai_2 _16184_ (.A1(_05333_),
    .A2(_05335_),
    .B1(_05364_),
    .Y(_05406_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_05366_),
    .B(_05399_),
    .Y(_05407_));
 sky130_fd_sc_hd__o21bai_1 _16186_ (.A1(_05374_),
    .A2(_05399_),
    .B1_N(_13319_),
    .Y(_05408_));
 sky130_fd_sc_hd__a211oi_4 _16187_ (.A1(_05406_),
    .A2(_05407_),
    .B1(_05408_),
    .C1(_05398_),
    .Y(_05409_));
 sky130_fd_sc_hd__xnor2_1 _16188_ (.A(_05405_),
    .B(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__nor2_1 _16189_ (.A(net537),
    .B(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__a21oi_4 _16190_ (.A1(\w[63][12] ),
    .A2(net537),
    .B1(_05411_),
    .Y(_05412_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1307 ();
 sky130_fd_sc_hd__nand2_1 _16192_ (.A(net708),
    .B(_05315_),
    .Y(_05414_));
 sky130_fd_sc_hd__o21ai_0 _16193_ (.A1(_05315_),
    .A2(_05412_),
    .B1(_05414_),
    .Y(_00356_));
 sky130_fd_sc_hd__or3_1 _16194_ (.A(_13319_),
    .B(_05398_),
    .C(_05400_),
    .X(_05415_));
 sky130_fd_sc_hd__a21oi_1 _16195_ (.A1(_13324_),
    .A2(_05415_),
    .B1(_13323_),
    .Y(_05416_));
 sky130_fd_sc_hd__xor2_2 _16196_ (.A(_13328_),
    .B(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__nor2_1 _16197_ (.A(net535),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__a21oi_4 _16198_ (.A1(\w[63][13] ),
    .A2(net535),
    .B1(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1306 ();
 sky130_fd_sc_hd__nand2_1 _16200_ (.A(net705),
    .B(_05315_),
    .Y(_05421_));
 sky130_fd_sc_hd__o21ai_0 _16201_ (.A1(_05315_),
    .A2(_05419_),
    .B1(_05421_),
    .Y(_00357_));
 sky130_fd_sc_hd__o21bai_1 _16202_ (.A1(_05405_),
    .A2(_05409_),
    .B1_N(_13323_),
    .Y(_05422_));
 sky130_fd_sc_hd__a21oi_1 _16203_ (.A1(_13328_),
    .A2(_05422_),
    .B1(_13327_),
    .Y(_05423_));
 sky130_fd_sc_hd__xor2_2 _16204_ (.A(_13332_),
    .B(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__nor2_2 _16205_ (.A(net534),
    .B(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__a21oi_4 _16206_ (.A1(\w[63][14] ),
    .A2(net532),
    .B1(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1305 ();
 sky130_fd_sc_hd__nand2_1 _16208_ (.A(net444),
    .B(_05315_),
    .Y(_05428_));
 sky130_fd_sc_hd__o21ai_0 _16209_ (.A1(_05315_),
    .A2(_05426_),
    .B1(_05428_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand3_1 _16210_ (.A(_13324_),
    .B(_13328_),
    .C(_13332_),
    .Y(_05429_));
 sky130_fd_sc_hd__inv_1 _16211_ (.A(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__o21ai_0 _16212_ (.A1(_05398_),
    .A2(_05400_),
    .B1(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__a21o_1 _16213_ (.A1(_13324_),
    .A2(_13319_),
    .B1(_13323_),
    .X(_05432_));
 sky130_fd_sc_hd__a21o_1 _16214_ (.A1(_13328_),
    .A2(_05432_),
    .B1(_13327_),
    .X(_05433_));
 sky130_fd_sc_hd__a21oi_1 _16215_ (.A1(_13332_),
    .A2(_05433_),
    .B1(_13331_),
    .Y(_05434_));
 sky130_fd_sc_hd__nand2_1 _16216_ (.A(_05431_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__xnor2_1 _16217_ (.A(_13336_),
    .B(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__nor2_2 _16218_ (.A(net537),
    .B(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__a21oi_4 _16219_ (.A1(\w[63][15] ),
    .A2(net532),
    .B1(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1304 ();
 sky130_fd_sc_hd__nand2_1 _16221_ (.A(net433),
    .B(_05315_),
    .Y(_05440_));
 sky130_fd_sc_hd__o21ai_0 _16222_ (.A1(_05315_),
    .A2(_05438_),
    .B1(_05440_),
    .Y(_00359_));
 sky130_fd_sc_hd__a21o_1 _16223_ (.A1(_13328_),
    .A2(_13323_),
    .B1(_13327_),
    .X(_05441_));
 sky130_fd_sc_hd__a21oi_1 _16224_ (.A1(_13332_),
    .A2(_05441_),
    .B1(_13331_),
    .Y(_05442_));
 sky130_fd_sc_hd__o21ai_0 _16225_ (.A1(_05409_),
    .A2(_05429_),
    .B1(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__a21oi_1 _16226_ (.A1(_13336_),
    .A2(_05443_),
    .B1(_13335_),
    .Y(_05444_));
 sky130_fd_sc_hd__xor2_1 _16227_ (.A(_13340_),
    .B(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__nor2_4 _16228_ (.A(net537),
    .B(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__a21oi_4 _16229_ (.A1(\w[63][16] ),
    .A2(net532),
    .B1(_05446_),
    .Y(_05447_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1303 ();
 sky130_fd_sc_hd__nand2_1 _16231_ (.A(net422),
    .B(_05315_),
    .Y(_05449_));
 sky130_fd_sc_hd__o21ai_0 _16232_ (.A1(_05315_),
    .A2(_05447_),
    .B1(_05449_),
    .Y(_00360_));
 sky130_fd_sc_hd__a21o_1 _16233_ (.A1(_13336_),
    .A2(_05435_),
    .B1(_13335_),
    .X(_05450_));
 sky130_fd_sc_hd__a21oi_2 _16234_ (.A1(_13340_),
    .A2(_05450_),
    .B1(_13339_),
    .Y(_05451_));
 sky130_fd_sc_hd__xnor2_4 _16235_ (.A(_13344_),
    .B(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__mux2i_4 _16236_ (.A0(_05452_),
    .A1(\w[63][17] ),
    .S(net532),
    .Y(_05453_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1302 ();
 sky130_fd_sc_hd__nand2_1 _16238_ (.A(net411),
    .B(_05315_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21ai_0 _16239_ (.A1(_05315_),
    .A2(_05453_),
    .B1(_05455_),
    .Y(_00361_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1301 ();
 sky130_fd_sc_hd__nand2_1 _16241_ (.A(_13336_),
    .B(_13340_),
    .Y(_05457_));
 sky130_fd_sc_hd__inv_1 _16242_ (.A(_13336_),
    .Y(_05458_));
 sky130_fd_sc_hd__o21bai_1 _16243_ (.A1(_05458_),
    .A2(_05442_),
    .B1_N(_13335_),
    .Y(_05459_));
 sky130_fd_sc_hd__a21oi_1 _16244_ (.A1(_13340_),
    .A2(_05459_),
    .B1(_13339_),
    .Y(_05460_));
 sky130_fd_sc_hd__o31ai_1 _16245_ (.A1(_05409_),
    .A2(_05429_),
    .A3(_05457_),
    .B1(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__a21oi_2 _16246_ (.A1(_13344_),
    .A2(_05461_),
    .B1(_13343_),
    .Y(_05462_));
 sky130_fd_sc_hd__xor2_2 _16247_ (.A(_13348_),
    .B(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__nor2_1 _16248_ (.A(net533),
    .B(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__a21oi_4 _16249_ (.A1(\w[63][18] ),
    .A2(net533),
    .B1(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1300 ();
 sky130_fd_sc_hd__nand2_1 _16251_ (.A(net400),
    .B(_05315_),
    .Y(_05467_));
 sky130_fd_sc_hd__o21ai_0 _16252_ (.A1(_05315_),
    .A2(_05465_),
    .B1(_05467_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_1 _16253_ (.A(_13344_),
    .B(_13348_),
    .Y(_05468_));
 sky130_fd_sc_hd__nor2_1 _16254_ (.A(_05457_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__a21o_1 _16255_ (.A1(_13340_),
    .A2(_13335_),
    .B1(_13339_),
    .X(_05470_));
 sky130_fd_sc_hd__a21o_1 _16256_ (.A1(_13344_),
    .A2(_05470_),
    .B1(_13343_),
    .X(_05471_));
 sky130_fd_sc_hd__a21oi_1 _16257_ (.A1(_13348_),
    .A2(_05471_),
    .B1(_13347_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2b_1 _16258_ (.A_N(_13352_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__a21oi_1 _16259_ (.A1(_05435_),
    .A2(_05469_),
    .B1(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__o31ai_1 _16260_ (.A1(_05434_),
    .A2(_05457_),
    .A3(_05468_),
    .B1(_05472_),
    .Y(_05475_));
 sky130_fd_sc_hd__nand2_1 _16261_ (.A(_13352_),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__o2111ai_4 _16262_ (.A1(_05398_),
    .A2(_05400_),
    .B1(_05430_),
    .C1(_05469_),
    .D1(_13352_),
    .Y(_05477_));
 sky130_fd_sc_hd__nand2_1 _16263_ (.A(_05476_),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__nor3_2 _16264_ (.A(net535),
    .B(_05474_),
    .C(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__a21oi_4 _16265_ (.A1(\w[63][19] ),
    .A2(net535),
    .B1(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1299 ();
 sky130_fd_sc_hd__nand2_1 _16267_ (.A(net389),
    .B(_05315_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21ai_0 _16268_ (.A1(_05315_),
    .A2(_05480_),
    .B1(_05482_),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_1 _16269_ (.A(_13348_),
    .B(_13352_),
    .Y(_05483_));
 sky130_fd_sc_hd__a21oi_1 _16270_ (.A1(_13352_),
    .A2(_13347_),
    .B1(_13351_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21ai_2 _16271_ (.A1(_05462_),
    .A2(_05483_),
    .B1(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__xnor2_1 _16272_ (.A(_13356_),
    .B(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__nor2_1 _16273_ (.A(net536),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__a21oi_4 _16274_ (.A1(\w[63][20] ),
    .A2(net536),
    .B1(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1297 ();
 sky130_fd_sc_hd__nand2_1 _16277_ (.A(net378),
    .B(_05315_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_0 _16278_ (.A1(_05315_),
    .A2(_05488_),
    .B1(_05491_),
    .Y(_00365_));
 sky130_fd_sc_hd__o21ai_0 _16279_ (.A1(_13351_),
    .A2(_05478_),
    .B1(_13356_),
    .Y(_05492_));
 sky130_fd_sc_hd__nor2_1 _16280_ (.A(_13360_),
    .B(_13355_),
    .Y(_05493_));
 sky130_fd_sc_hd__nor2_1 _16281_ (.A(_13351_),
    .B(_13355_),
    .Y(_05494_));
 sky130_fd_sc_hd__o21ai_1 _16282_ (.A1(_13356_),
    .A2(_13355_),
    .B1(_13360_),
    .Y(_05495_));
 sky130_fd_sc_hd__a31oi_4 _16283_ (.A1(_05476_),
    .A2(_05477_),
    .A3(_05494_),
    .B1(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__a211oi_2 _16284_ (.A1(_05492_),
    .A2(_05493_),
    .B1(_05496_),
    .C1(net535),
    .Y(_05497_));
 sky130_fd_sc_hd__a21oi_4 _16285_ (.A1(\w[63][21] ),
    .A2(net535),
    .B1(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1296 ();
 sky130_fd_sc_hd__nand2_1 _16287_ (.A(net367),
    .B(_05315_),
    .Y(_05500_));
 sky130_fd_sc_hd__o21ai_0 _16288_ (.A1(_05315_),
    .A2(_05498_),
    .B1(_05500_),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _16289_ (.A(_13364_),
    .B(_13359_),
    .Y(_05501_));
 sky130_fd_sc_hd__nand3_1 _16290_ (.A(_13360_),
    .B(_13364_),
    .C(_13355_),
    .Y(_05502_));
 sky130_fd_sc_hd__nand2_1 _16291_ (.A(_05501_),
    .B(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__a41oi_4 _16292_ (.A1(_13356_),
    .A2(_13360_),
    .A3(_13364_),
    .A4(_05485_),
    .B1(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__a21o_1 _16293_ (.A1(_13356_),
    .A2(_05485_),
    .B1(_13355_),
    .X(_05505_));
 sky130_fd_sc_hd__a211o_1 _16294_ (.A1(_13360_),
    .A2(_05505_),
    .B1(_13359_),
    .C1(_13364_),
    .X(_05506_));
 sky130_fd_sc_hd__nand2_1 _16295_ (.A(_05504_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__nor2_2 _16296_ (.A(net535),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__a21oi_4 _16297_ (.A1(\w[63][22] ),
    .A2(net533),
    .B1(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1295 ();
 sky130_fd_sc_hd__nand2_1 _16299_ (.A(net356),
    .B(_05315_),
    .Y(_05511_));
 sky130_fd_sc_hd__o21ai_0 _16300_ (.A1(_05315_),
    .A2(_05509_),
    .B1(_05511_),
    .Y(_00367_));
 sky130_fd_sc_hd__o21a_1 _16301_ (.A1(_13359_),
    .A2(_05496_),
    .B1(_13364_),
    .X(_05512_));
 sky130_fd_sc_hd__nor2_1 _16302_ (.A(_13363_),
    .B(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hd__xnor2_2 _16303_ (.A(_13368_),
    .B(_05513_),
    .Y(_05514_));
 sky130_fd_sc_hd__mux2i_4 _16304_ (.A0(_05514_),
    .A1(\w[63][23] ),
    .S(net534),
    .Y(_05515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1294 ();
 sky130_fd_sc_hd__nand2_1 _16306_ (.A(net345),
    .B(_05315_),
    .Y(_05517_));
 sky130_fd_sc_hd__o21ai_0 _16307_ (.A1(_05315_),
    .A2(_05515_),
    .B1(_05517_),
    .Y(_00368_));
 sky130_fd_sc_hd__nor2_1 _16308_ (.A(_13363_),
    .B(_13367_),
    .Y(_05518_));
 sky130_fd_sc_hd__nor2_1 _16309_ (.A(_13368_),
    .B(_13367_),
    .Y(_05519_));
 sky130_fd_sc_hd__a21oi_2 _16310_ (.A1(_05504_),
    .A2(_05518_),
    .B1(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__xnor2_4 _16311_ (.A(_13372_),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__nor2_1 _16312_ (.A(net532),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__a21oi_4 _16313_ (.A1(\w[63][24] ),
    .A2(net532),
    .B1(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1293 ();
 sky130_fd_sc_hd__nand2_1 _16315_ (.A(net333),
    .B(_05315_),
    .Y(_05525_));
 sky130_fd_sc_hd__o21ai_0 _16316_ (.A1(_05315_),
    .A2(_05523_),
    .B1(_05525_),
    .Y(_00369_));
 sky130_fd_sc_hd__a21o_1 _16317_ (.A1(_13372_),
    .A2(_13367_),
    .B1(_13371_),
    .X(_05526_));
 sky130_fd_sc_hd__or3_1 _16318_ (.A(_13359_),
    .B(_13363_),
    .C(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__a21oi_1 _16319_ (.A1(_13368_),
    .A2(_13372_),
    .B1(_05526_),
    .Y(_05528_));
 sky130_fd_sc_hd__nor3_1 _16320_ (.A(_13364_),
    .B(_13363_),
    .C(_05526_),
    .Y(_05529_));
 sky130_fd_sc_hd__nor2_1 _16321_ (.A(_05528_),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__o211a_1 _16322_ (.A1(_05496_),
    .A2(_05527_),
    .B1(_05530_),
    .C1(_13376_),
    .X(_05531_));
 sky130_fd_sc_hd__o21a_1 _16323_ (.A1(_05496_),
    .A2(_05527_),
    .B1(_05530_),
    .X(_05532_));
 sky130_fd_sc_hd__nor2_1 _16324_ (.A(_13376_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__nor3_4 _16325_ (.A(net534),
    .B(_05531_),
    .C(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__a21oi_4 _16326_ (.A1(\w[63][25] ),
    .A2(net532),
    .B1(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1292 ();
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(net322),
    .B(_05315_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_0 _16329_ (.A1(_05315_),
    .A2(_05535_),
    .B1(_05537_),
    .Y(_00370_));
 sky130_fd_sc_hd__nor3_1 _16330_ (.A(_13363_),
    .B(_13367_),
    .C(_13371_),
    .Y(_05538_));
 sky130_fd_sc_hd__a21oi_4 _16331_ (.A1(_05504_),
    .A2(_05538_),
    .B1(_05528_),
    .Y(_05539_));
 sky130_fd_sc_hd__a21oi_2 _16332_ (.A1(_13376_),
    .A2(_05539_),
    .B1(_13375_),
    .Y(_05540_));
 sky130_fd_sc_hd__xnor2_4 _16333_ (.A(_13380_),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__mux2i_4 _16334_ (.A0(_05541_),
    .A1(\w[63][26] ),
    .S(net534),
    .Y(_05542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1291 ();
 sky130_fd_sc_hd__nand2_1 _16336_ (.A(net311),
    .B(_05315_),
    .Y(_05544_));
 sky130_fd_sc_hd__o21ai_0 _16337_ (.A1(_05315_),
    .A2(_05542_),
    .B1(_05544_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_1 _16338_ (.A(_13379_),
    .Y(_05545_));
 sky130_fd_sc_hd__o21ai_1 _16339_ (.A1(_13375_),
    .A2(_05531_),
    .B1(_13380_),
    .Y(_05546_));
 sky130_fd_sc_hd__inv_1 _16340_ (.A(_13384_),
    .Y(_05547_));
 sky130_fd_sc_hd__a21oi_2 _16341_ (.A1(_05545_),
    .A2(_05546_),
    .B1(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__and3_1 _16342_ (.A(_05547_),
    .B(_05545_),
    .C(_05546_),
    .X(_05549_));
 sky130_fd_sc_hd__nand2_1 _16343_ (.A(\w[63][27] ),
    .B(net534),
    .Y(_05550_));
 sky130_fd_sc_hd__o31a_4 _16344_ (.A1(net534),
    .A2(_05548_),
    .A3(_05549_),
    .B1(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1290 ();
 sky130_fd_sc_hd__nand2_1 _16346_ (.A(net300),
    .B(_05315_),
    .Y(_05553_));
 sky130_fd_sc_hd__o21ai_0 _16347_ (.A1(_05315_),
    .A2(_05551_),
    .B1(_05553_),
    .Y(_00372_));
 sky130_fd_sc_hd__and3_1 _16348_ (.A(_13376_),
    .B(_13380_),
    .C(_13384_),
    .X(_05554_));
 sky130_fd_sc_hd__a21oi_1 _16349_ (.A1(_13380_),
    .A2(_13375_),
    .B1(_13379_),
    .Y(_05555_));
 sky130_fd_sc_hd__nor2_1 _16350_ (.A(_05547_),
    .B(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__a211oi_2 _16351_ (.A1(_05539_),
    .A2(_05554_),
    .B1(_05556_),
    .C1(_13383_),
    .Y(_05557_));
 sky130_fd_sc_hd__xnor2_2 _16352_ (.A(_13388_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__mux2i_4 _16353_ (.A0(_05558_),
    .A1(\w[63][28] ),
    .S(net533),
    .Y(_05559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1289 ();
 sky130_fd_sc_hd__nand2_1 _16355_ (.A(net289),
    .B(_05315_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21ai_0 _16356_ (.A1(_05315_),
    .A2(_05559_),
    .B1(_05561_),
    .Y(_00373_));
 sky130_fd_sc_hd__and4_1 _16357_ (.A(_13376_),
    .B(_13380_),
    .C(_13384_),
    .D(_13388_),
    .X(_05562_));
 sky130_fd_sc_hd__o21ai_0 _16358_ (.A1(_13383_),
    .A2(_05556_),
    .B1(_13388_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2b_2 _16359_ (.A_N(_13387_),
    .B(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__a21oi_2 _16360_ (.A1(_05532_),
    .A2(_05562_),
    .B1(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__xnor2_4 _16361_ (.A(_13392_),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__mux2i_4 _16362_ (.A0(_05566_),
    .A1(\w[63][29] ),
    .S(net533),
    .Y(_05567_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1288 ();
 sky130_fd_sc_hd__nand2_1 _16364_ (.A(net278),
    .B(_05315_),
    .Y(_05569_));
 sky130_fd_sc_hd__o21ai_0 _16365_ (.A1(_05315_),
    .A2(_05567_),
    .B1(_05569_),
    .Y(_00374_));
 sky130_fd_sc_hd__and2_0 _16366_ (.A(_13392_),
    .B(_05562_),
    .X(_05570_));
 sky130_fd_sc_hd__a221oi_4 _16367_ (.A1(_13392_),
    .A2(_05564_),
    .B1(_05570_),
    .B2(_05539_),
    .C1(_13391_),
    .Y(_05571_));
 sky130_fd_sc_hd__xnor2_4 _16368_ (.A(_13396_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__mux2i_4 _16369_ (.A0(_05572_),
    .A1(\w[63][30] ),
    .S(net533),
    .Y(_05573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1287 ();
 sky130_fd_sc_hd__nand2_1 _16371_ (.A(net267),
    .B(_05315_),
    .Y(_05575_));
 sky130_fd_sc_hd__o21ai_0 _16372_ (.A1(_05315_),
    .A2(_05573_),
    .B1(_05575_),
    .Y(_00376_));
 sky130_fd_sc_hd__o211ai_1 _16373_ (.A1(_05496_),
    .A2(_05527_),
    .B1(_05530_),
    .C1(_05562_),
    .Y(_05576_));
 sky130_fd_sc_hd__nor3_1 _16374_ (.A(_13391_),
    .B(_13395_),
    .C(_05564_),
    .Y(_05577_));
 sky130_fd_sc_hd__or2_0 _16375_ (.A(_13392_),
    .B(_13391_),
    .X(_05578_));
 sky130_fd_sc_hd__a21oi_1 _16376_ (.A1(_13396_),
    .A2(_05578_),
    .B1(_13395_),
    .Y(_05579_));
 sky130_fd_sc_hd__a21oi_2 _16377_ (.A1(_05576_),
    .A2(_05577_),
    .B1(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__xor2_1 _16378_ (.A(_12241_),
    .B(_12244_),
    .X(_05581_));
 sky130_fd_sc_hd__mux4_1 _16379_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net638),
    .S1(net643),
    .X(_05582_));
 sky130_fd_sc_hd__mux4_1 _16380_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net638),
    .S1(net643),
    .X(_05583_));
 sky130_fd_sc_hd__mux4_1 _16381_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net638),
    .S1(net643),
    .X(_05584_));
 sky130_fd_sc_hd__mux4_1 _16382_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net638),
    .S1(net643),
    .X(_05585_));
 sky130_fd_sc_hd__mux4_4 _16383_ (.A0(_05582_),
    .A1(_05583_),
    .A2(_05584_),
    .A3(_05585_),
    .S0(net633),
    .S1(net632),
    .X(_05586_));
 sky130_fd_sc_hd__mux4_1 _16384_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net635),
    .S1(net644),
    .X(_05587_));
 sky130_fd_sc_hd__mux4_1 _16385_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net635),
    .S1(net644),
    .X(_05588_));
 sky130_fd_sc_hd__mux4_1 _16386_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net635),
    .S1(net644),
    .X(_05589_));
 sky130_fd_sc_hd__mux4_1 _16387_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net635),
    .S1(net644),
    .X(_05590_));
 sky130_fd_sc_hd__mux4_1 _16388_ (.A0(_05587_),
    .A1(_05588_),
    .A2(_05589_),
    .A3(_05590_),
    .S0(net634),
    .S1(net632),
    .X(_05591_));
 sky130_fd_sc_hd__mux2i_4 _16389_ (.A0(_05586_),
    .A1(_05591_),
    .S(net629),
    .Y(_05592_));
 sky130_fd_sc_hd__xnor2_1 _16390_ (.A(_05581_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__mux4_1 _16391_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net563),
    .S1(net568),
    .X(_05594_));
 sky130_fd_sc_hd__mux4_1 _16392_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net563),
    .S1(net568),
    .X(_05595_));
 sky130_fd_sc_hd__mux4_1 _16393_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net563),
    .S1(net568),
    .X(_05596_));
 sky130_fd_sc_hd__mux4_1 _16394_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net563),
    .S1(net568),
    .X(_05597_));
 sky130_fd_sc_hd__mux4_4 _16395_ (.A0(_05594_),
    .A1(_05595_),
    .A2(_05596_),
    .A3(_05597_),
    .S0(net558),
    .S1(net556),
    .X(_05598_));
 sky130_fd_sc_hd__mux4_1 _16396_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net564),
    .S1(net568),
    .X(_05599_));
 sky130_fd_sc_hd__mux4_1 _16397_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net563),
    .S1(net569),
    .X(_05600_));
 sky130_fd_sc_hd__mux4_1 _16398_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net563),
    .S1(net569),
    .X(_05601_));
 sky130_fd_sc_hd__mux4_1 _16399_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net563),
    .S1(net569),
    .X(_05602_));
 sky130_fd_sc_hd__mux4_1 _16400_ (.A0(_05599_),
    .A1(_05600_),
    .A2(_05601_),
    .A3(_05602_),
    .S0(net558),
    .S1(net556),
    .X(_05603_));
 sky130_fd_sc_hd__mux2i_4 _16401_ (.A0(_05598_),
    .A1(_05603_),
    .S(net554),
    .Y(_05604_));
 sky130_fd_sc_hd__xnor2_4 _16402_ (.A(_03817_),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__xnor2_2 _16403_ (.A(_05593_),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__xor2_1 _16404_ (.A(_03366_),
    .B(_03551_),
    .X(_05607_));
 sky130_fd_sc_hd__xnor2_2 _16405_ (.A(_03135_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__xnor2_4 _16406_ (.A(_05606_),
    .B(_05608_),
    .Y(_05609_));
 sky130_fd_sc_hd__xnor2_4 _16407_ (.A(_05580_),
    .B(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__mux2i_4 _16408_ (.A0(_05610_),
    .A1(\w[63][31] ),
    .S(net533),
    .Y(_05611_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1286 ();
 sky130_fd_sc_hd__nand2_1 _16410_ (.A(net256),
    .B(_05315_),
    .Y(_05613_));
 sky130_fd_sc_hd__o21ai_0 _16411_ (.A1(_05315_),
    .A2(_05611_),
    .B1(_05613_),
    .Y(_00377_));
 sky130_fd_sc_hd__nor2b_4 _16412_ (.A(net762),
    .B_N(_13699_),
    .Y(_05614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1285 ();
 sky130_fd_sc_hd__nand2_8 _16414_ (.A(_09897_),
    .B(_05614_),
    .Y(_05616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1283 ();
 sky130_fd_sc_hd__nand2_1 _16417_ (.A(net756),
    .B(_05616_),
    .Y(_05619_));
 sky130_fd_sc_hd__o21ai_0 _16418_ (.A1(_04988_),
    .A2(_05616_),
    .B1(_05619_),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _16419_ (.A(net755),
    .B(_05616_),
    .Y(_05620_));
 sky130_fd_sc_hd__o21ai_0 _16420_ (.A1(_04992_),
    .A2(_05616_),
    .B1(_05620_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _16421_ (.A(net754),
    .B(_05616_),
    .Y(_05621_));
 sky130_fd_sc_hd__o21ai_0 _16422_ (.A1(_04995_),
    .A2(_05616_),
    .B1(_05621_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand2_1 _16423_ (.A(net753),
    .B(_05616_),
    .Y(_05622_));
 sky130_fd_sc_hd__o21ai_0 _16424_ (.A1(_05003_),
    .A2(_05616_),
    .B1(_05622_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _16425_ (.A(net752),
    .B(_05616_),
    .Y(_05623_));
 sky130_fd_sc_hd__o21ai_0 _16426_ (.A1(_05012_),
    .A2(_05616_),
    .B1(_05623_),
    .Y(_00411_));
 sky130_fd_sc_hd__nand2_1 _16427_ (.A(net751),
    .B(_05616_),
    .Y(_05624_));
 sky130_fd_sc_hd__o21ai_0 _16428_ (.A1(_05021_),
    .A2(_05616_),
    .B1(_05624_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _16429_ (.A(net749),
    .B(_05616_),
    .Y(_05625_));
 sky130_fd_sc_hd__o21ai_0 _16430_ (.A1(_05032_),
    .A2(_05616_),
    .B1(_05625_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _16431_ (.A(net748),
    .B(_05616_),
    .Y(_05626_));
 sky130_fd_sc_hd__o21ai_0 _16432_ (.A1(_05039_),
    .A2(_05616_),
    .B1(_05626_),
    .Y(_00414_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1282 ();
 sky130_fd_sc_hd__nand2_1 _16434_ (.A(net747),
    .B(_05616_),
    .Y(_05628_));
 sky130_fd_sc_hd__o21ai_0 _16435_ (.A1(_05048_),
    .A2(_05616_),
    .B1(_05628_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _16436_ (.A(net746),
    .B(_05616_),
    .Y(_05629_));
 sky130_fd_sc_hd__o21ai_0 _16437_ (.A1(_05055_),
    .A2(_05616_),
    .B1(_05629_),
    .Y(_00416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1281 ();
 sky130_fd_sc_hd__nand2_1 _16439_ (.A(net745),
    .B(_05616_),
    .Y(_05631_));
 sky130_fd_sc_hd__o21ai_0 _16440_ (.A1(_05062_),
    .A2(_05616_),
    .B1(_05631_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _16441_ (.A(net744),
    .B(_05616_),
    .Y(_05632_));
 sky130_fd_sc_hd__o21ai_0 _16442_ (.A1(_05077_),
    .A2(_05616_),
    .B1(_05632_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(net743),
    .B(_05616_),
    .Y(_05633_));
 sky130_fd_sc_hd__o21ai_0 _16444_ (.A1(_05087_),
    .A2(_05616_),
    .B1(_05633_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _16445_ (.A(net742),
    .B(_05616_),
    .Y(_05634_));
 sky130_fd_sc_hd__o21ai_0 _16446_ (.A1(_05095_),
    .A2(_05616_),
    .B1(_05634_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _16447_ (.A(net741),
    .B(_05616_),
    .Y(_05635_));
 sky130_fd_sc_hd__o21ai_0 _16448_ (.A1(_05102_),
    .A2(_05616_),
    .B1(_05635_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _16449_ (.A(net740),
    .B(_05616_),
    .Y(_05636_));
 sky130_fd_sc_hd__o21ai_0 _16450_ (.A1(_05112_),
    .A2(_05616_),
    .B1(_05636_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_1 _16451_ (.A(net738),
    .B(_05616_),
    .Y(_05637_));
 sky130_fd_sc_hd__o21ai_0 _16452_ (.A1(_05121_),
    .A2(_05616_),
    .B1(_05637_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand2_1 _16453_ (.A(net737),
    .B(_05616_),
    .Y(_05638_));
 sky130_fd_sc_hd__o21ai_0 _16454_ (.A1(_05128_),
    .A2(_05616_),
    .B1(_05638_),
    .Y(_00393_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1280 ();
 sky130_fd_sc_hd__nand2_1 _16456_ (.A(net736),
    .B(_05616_),
    .Y(_05640_));
 sky130_fd_sc_hd__o21ai_0 _16457_ (.A1(_05137_),
    .A2(_05616_),
    .B1(_05640_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _16458_ (.A(net735),
    .B(_05616_),
    .Y(_05641_));
 sky130_fd_sc_hd__o21ai_0 _16459_ (.A1(_05154_),
    .A2(_05616_),
    .B1(_05641_),
    .Y(_00395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1279 ();
 sky130_fd_sc_hd__nand2_1 _16461_ (.A(net734),
    .B(_05616_),
    .Y(_05643_));
 sky130_fd_sc_hd__o21ai_0 _16462_ (.A1(_05167_),
    .A2(_05616_),
    .B1(_05643_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _16463_ (.A(net733),
    .B(_05616_),
    .Y(_05644_));
 sky130_fd_sc_hd__o21ai_0 _16464_ (.A1(_05175_),
    .A2(_05616_),
    .B1(_05644_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _16465_ (.A(net732),
    .B(_05616_),
    .Y(_05645_));
 sky130_fd_sc_hd__o21ai_0 _16466_ (.A1(_05184_),
    .A2(_05616_),
    .B1(_05645_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _16467_ (.A(net731),
    .B(_05616_),
    .Y(_05646_));
 sky130_fd_sc_hd__o21ai_0 _16468_ (.A1(_05196_),
    .A2(_05616_),
    .B1(_05646_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _16469_ (.A(net730),
    .B(_05616_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_0 _16470_ (.A1(_05206_),
    .A2(_05616_),
    .B1(_05647_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _16471_ (.A(net729),
    .B(_05616_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_0 _16472_ (.A1(_05214_),
    .A2(_05616_),
    .B1(_05648_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _16473_ (.A(net727),
    .B(_05616_),
    .Y(_05649_));
 sky130_fd_sc_hd__o21ai_0 _16474_ (.A1(_05224_),
    .A2(_05616_),
    .B1(_05649_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(net726),
    .B(_05616_),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_0 _16476_ (.A1(_05236_),
    .A2(_05616_),
    .B1(_05650_),
    .Y(_00404_));
 sky130_fd_sc_hd__nand2_1 _16477_ (.A(net725),
    .B(_05616_),
    .Y(_05651_));
 sky130_fd_sc_hd__o21ai_0 _16478_ (.A1(_05243_),
    .A2(_05616_),
    .B1(_05651_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _16479_ (.A(net724),
    .B(_05616_),
    .Y(_05652_));
 sky130_fd_sc_hd__o21ai_0 _16480_ (.A1(_05251_),
    .A2(_05616_),
    .B1(_05652_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _16481_ (.A(net723),
    .B(_05616_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21ai_0 _16482_ (.A1(_05260_),
    .A2(_05616_),
    .B1(_05653_),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _16483_ (.A(net722),
    .B(_05616_),
    .Y(_05654_));
 sky130_fd_sc_hd__o21ai_0 _16484_ (.A1(_05310_),
    .A2(_05616_),
    .B1(_05654_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2b_4 _16485_ (.A(net762),
    .B_N(_13707_),
    .Y(_05655_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1278 ();
 sky130_fd_sc_hd__nand2_8 _16487_ (.A(_09959_),
    .B(_05655_),
    .Y(_05657_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1276 ();
 sky130_fd_sc_hd__nand2_1 _16490_ (.A(net31),
    .B(_05657_),
    .Y(_05660_));
 sky130_fd_sc_hd__o21ai_0 _16491_ (.A1(_05317_),
    .A2(_05657_),
    .B1(_05660_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _16492_ (.A(net30),
    .B(_05657_),
    .Y(_05661_));
 sky130_fd_sc_hd__o21ai_0 _16493_ (.A1(_05321_),
    .A2(_05657_),
    .B1(_05661_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _16494_ (.A(net29),
    .B(_05657_),
    .Y(_05662_));
 sky130_fd_sc_hd__o21ai_0 _16495_ (.A1(_05324_),
    .A2(_05657_),
    .B1(_05662_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _16496_ (.A(net28),
    .B(_05657_),
    .Y(_05663_));
 sky130_fd_sc_hd__o21ai_0 _16497_ (.A1(_05330_),
    .A2(_05657_),
    .B1(_05663_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _16498_ (.A(net27),
    .B(_05657_),
    .Y(_05664_));
 sky130_fd_sc_hd__o21ai_0 _16499_ (.A1(_05338_),
    .A2(_05657_),
    .B1(_05664_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _16500_ (.A(net26),
    .B(_05657_),
    .Y(_05665_));
 sky130_fd_sc_hd__o21ai_0 _16501_ (.A1(_05347_),
    .A2(_05657_),
    .B1(_05665_),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _16502_ (.A(net25),
    .B(_05657_),
    .Y(_05666_));
 sky130_fd_sc_hd__o21ai_0 _16503_ (.A1(_05354_),
    .A2(_05657_),
    .B1(_05666_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _16504_ (.A(net24),
    .B(_05657_),
    .Y(_05667_));
 sky130_fd_sc_hd__o21ai_0 _16505_ (.A1(_05360_),
    .A2(_05657_),
    .B1(_05667_),
    .Y(_00446_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1275 ();
 sky130_fd_sc_hd__nand2_1 _16507_ (.A(net22),
    .B(_05657_),
    .Y(_05669_));
 sky130_fd_sc_hd__o21ai_0 _16508_ (.A1(_05371_),
    .A2(_05657_),
    .B1(_05669_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand2_1 _16509_ (.A(net21),
    .B(_05657_),
    .Y(_05670_));
 sky130_fd_sc_hd__o21ai_0 _16510_ (.A1(_05380_),
    .A2(_05657_),
    .B1(_05670_),
    .Y(_00448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1274 ();
 sky130_fd_sc_hd__nand2_1 _16512_ (.A(net20),
    .B(_05657_),
    .Y(_05672_));
 sky130_fd_sc_hd__o21ai_0 _16513_ (.A1(_05388_),
    .A2(_05657_),
    .B1(_05672_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _16514_ (.A(net19),
    .B(_05657_),
    .Y(_05673_));
 sky130_fd_sc_hd__o21ai_0 _16515_ (.A1(_05402_),
    .A2(_05657_),
    .B1(_05673_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _16516_ (.A(net18),
    .B(_05657_),
    .Y(_05674_));
 sky130_fd_sc_hd__o21ai_0 _16517_ (.A1(_05412_),
    .A2(_05657_),
    .B1(_05674_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _16518_ (.A(net17),
    .B(_05657_),
    .Y(_05675_));
 sky130_fd_sc_hd__o21ai_0 _16519_ (.A1(_05419_),
    .A2(_05657_),
    .B1(_05675_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _16520_ (.A(net16),
    .B(_05657_),
    .Y(_05676_));
 sky130_fd_sc_hd__o21ai_0 _16521_ (.A1(_05426_),
    .A2(_05657_),
    .B1(_05676_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _16522_ (.A(net15),
    .B(_05657_),
    .Y(_05677_));
 sky130_fd_sc_hd__o21ai_0 _16523_ (.A1(_05438_),
    .A2(_05657_),
    .B1(_05677_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _16524_ (.A(net14),
    .B(_05657_),
    .Y(_05678_));
 sky130_fd_sc_hd__o21ai_0 _16525_ (.A1(_05447_),
    .A2(_05657_),
    .B1(_05678_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _16526_ (.A(net13),
    .B(_05657_),
    .Y(_05679_));
 sky130_fd_sc_hd__o21ai_0 _16527_ (.A1(_05453_),
    .A2(_05657_),
    .B1(_05679_),
    .Y(_00425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1273 ();
 sky130_fd_sc_hd__nand2_1 _16529_ (.A(net11),
    .B(_05657_),
    .Y(_05681_));
 sky130_fd_sc_hd__o21ai_0 _16530_ (.A1(_05465_),
    .A2(_05657_),
    .B1(_05681_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _16531_ (.A(net10),
    .B(_05657_),
    .Y(_05682_));
 sky130_fd_sc_hd__o21ai_0 _16532_ (.A1(_05480_),
    .A2(_05657_),
    .B1(_05682_),
    .Y(_00427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1272 ();
 sky130_fd_sc_hd__nand2_1 _16534_ (.A(net9),
    .B(_05657_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21ai_0 _16535_ (.A1(_05488_),
    .A2(_05657_),
    .B1(_05684_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _16536_ (.A(net8),
    .B(_05657_),
    .Y(_05685_));
 sky130_fd_sc_hd__o21ai_0 _16537_ (.A1(_05498_),
    .A2(_05657_),
    .B1(_05685_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _16538_ (.A(net7),
    .B(_05657_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21ai_0 _16539_ (.A1(_05509_),
    .A2(_05657_),
    .B1(_05686_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _16540_ (.A(net6),
    .B(_05657_),
    .Y(_05687_));
 sky130_fd_sc_hd__o21ai_0 _16541_ (.A1(_05515_),
    .A2(_05657_),
    .B1(_05687_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _16542_ (.A(net5),
    .B(_05657_),
    .Y(_05688_));
 sky130_fd_sc_hd__o21ai_0 _16543_ (.A1(_05523_),
    .A2(_05657_),
    .B1(_05688_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _16544_ (.A(net4),
    .B(_05657_),
    .Y(_05689_));
 sky130_fd_sc_hd__o21ai_0 _16545_ (.A1(_05535_),
    .A2(_05657_),
    .B1(_05689_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _16546_ (.A(net3),
    .B(_05657_),
    .Y(_05690_));
 sky130_fd_sc_hd__o21ai_0 _16547_ (.A1(_05542_),
    .A2(_05657_),
    .B1(_05690_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _16548_ (.A(net2),
    .B(_05657_),
    .Y(_05691_));
 sky130_fd_sc_hd__o21ai_0 _16549_ (.A1(_05551_),
    .A2(_05657_),
    .B1(_05691_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _16550_ (.A(net760),
    .B(_05657_),
    .Y(_05692_));
 sky130_fd_sc_hd__o21ai_0 _16551_ (.A1(_05559_),
    .A2(_05657_),
    .B1(_05692_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _16552_ (.A(net759),
    .B(_05657_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_0 _16553_ (.A1(_05567_),
    .A2(_05657_),
    .B1(_05693_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _16554_ (.A(net758),
    .B(_05657_),
    .Y(_05694_));
 sky130_fd_sc_hd__o21ai_0 _16555_ (.A1(_05573_),
    .A2(_05657_),
    .B1(_05694_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _16556_ (.A(net757),
    .B(_05657_),
    .Y(_05695_));
 sky130_fd_sc_hd__o21ai_0 _16557_ (.A1(_05611_),
    .A2(_05657_),
    .B1(_05695_),
    .Y(_00441_));
 sky130_fd_sc_hd__nor2b_4 _16558_ (.A(net762),
    .B_N(_13697_),
    .Y(_05696_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1271 ();
 sky130_fd_sc_hd__nand2_8 _16560_ (.A(_09897_),
    .B(_05696_),
    .Y(_05698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1269 ();
 sky130_fd_sc_hd__nand2_1 _16563_ (.A(net66),
    .B(_05698_),
    .Y(_05701_));
 sky130_fd_sc_hd__o21ai_0 _16564_ (.A1(_04988_),
    .A2(_05698_),
    .B1(_05701_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _16565_ (.A(net65),
    .B(_05698_),
    .Y(_05702_));
 sky130_fd_sc_hd__o21ai_0 _16566_ (.A1(_04992_),
    .A2(_05698_),
    .B1(_05702_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _16567_ (.A(net64),
    .B(_05698_),
    .Y(_05703_));
 sky130_fd_sc_hd__o21ai_0 _16568_ (.A1(_04995_),
    .A2(_05698_),
    .B1(_05703_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _16569_ (.A(net63),
    .B(_05698_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21ai_0 _16570_ (.A1(_05003_),
    .A2(_05698_),
    .B1(_05704_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _16571_ (.A(net62),
    .B(_05698_),
    .Y(_05705_));
 sky130_fd_sc_hd__o21ai_0 _16572_ (.A1(_05012_),
    .A2(_05698_),
    .B1(_05705_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _16573_ (.A(net61),
    .B(_05698_),
    .Y(_05706_));
 sky130_fd_sc_hd__o21ai_0 _16574_ (.A1(_05021_),
    .A2(_05698_),
    .B1(_05706_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _16575_ (.A(net60),
    .B(_05698_),
    .Y(_05707_));
 sky130_fd_sc_hd__o21ai_0 _16576_ (.A1(_05032_),
    .A2(_05698_),
    .B1(_05707_),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _16577_ (.A(net59),
    .B(_05698_),
    .Y(_05708_));
 sky130_fd_sc_hd__o21ai_0 _16578_ (.A1(_05039_),
    .A2(_05698_),
    .B1(_05708_),
    .Y(_00478_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1268 ();
 sky130_fd_sc_hd__nand2_1 _16580_ (.A(net58),
    .B(_05698_),
    .Y(_05710_));
 sky130_fd_sc_hd__o21ai_0 _16581_ (.A1(_05048_),
    .A2(_05698_),
    .B1(_05710_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _16582_ (.A(net57),
    .B(_05698_),
    .Y(_05711_));
 sky130_fd_sc_hd__o21ai_0 _16583_ (.A1(_05055_),
    .A2(_05698_),
    .B1(_05711_),
    .Y(_00480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1267 ();
 sky130_fd_sc_hd__nand2_1 _16585_ (.A(net55),
    .B(_05698_),
    .Y(_05713_));
 sky130_fd_sc_hd__o21ai_0 _16586_ (.A1(_05062_),
    .A2(_05698_),
    .B1(_05713_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _16587_ (.A(net54),
    .B(_05698_),
    .Y(_05714_));
 sky130_fd_sc_hd__o21ai_0 _16588_ (.A1(_05077_),
    .A2(_05698_),
    .B1(_05714_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _16589_ (.A(net53),
    .B(_05698_),
    .Y(_05715_));
 sky130_fd_sc_hd__o21ai_0 _16590_ (.A1(_05087_),
    .A2(_05698_),
    .B1(_05715_),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _16591_ (.A(net52),
    .B(_05698_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_0 _16592_ (.A1(_05095_),
    .A2(_05698_),
    .B1(_05716_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _16593_ (.A(net51),
    .B(_05698_),
    .Y(_05717_));
 sky130_fd_sc_hd__o21ai_0 _16594_ (.A1(_05102_),
    .A2(_05698_),
    .B1(_05717_),
    .Y(_00454_));
 sky130_fd_sc_hd__nand2_1 _16595_ (.A(net50),
    .B(_05698_),
    .Y(_05718_));
 sky130_fd_sc_hd__o21ai_0 _16596_ (.A1(_05112_),
    .A2(_05698_),
    .B1(_05718_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _16597_ (.A(net49),
    .B(_05698_),
    .Y(_05719_));
 sky130_fd_sc_hd__o21ai_0 _16598_ (.A1(_05121_),
    .A2(_05698_),
    .B1(_05719_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _16599_ (.A(net48),
    .B(_05698_),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ai_0 _16600_ (.A1(_05128_),
    .A2(_05698_),
    .B1(_05720_),
    .Y(_00457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1266 ();
 sky130_fd_sc_hd__nand2_1 _16602_ (.A(net47),
    .B(_05698_),
    .Y(_05722_));
 sky130_fd_sc_hd__o21ai_0 _16603_ (.A1(_05137_),
    .A2(_05698_),
    .B1(_05722_),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _16604_ (.A(net46),
    .B(_05698_),
    .Y(_05723_));
 sky130_fd_sc_hd__o21ai_0 _16605_ (.A1(_05154_),
    .A2(_05698_),
    .B1(_05723_),
    .Y(_00459_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1265 ();
 sky130_fd_sc_hd__nand2_1 _16607_ (.A(net44),
    .B(_05698_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_0 _16608_ (.A1(_05167_),
    .A2(_05698_),
    .B1(_05725_),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _16609_ (.A(net43),
    .B(_05698_),
    .Y(_05726_));
 sky130_fd_sc_hd__o21ai_0 _16610_ (.A1(_05175_),
    .A2(_05698_),
    .B1(_05726_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _16611_ (.A(net42),
    .B(_05698_),
    .Y(_05727_));
 sky130_fd_sc_hd__o21ai_0 _16612_ (.A1(_05184_),
    .A2(_05698_),
    .B1(_05727_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _16613_ (.A(net41),
    .B(_05698_),
    .Y(_05728_));
 sky130_fd_sc_hd__o21ai_0 _16614_ (.A1(_05196_),
    .A2(_05698_),
    .B1(_05728_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _16615_ (.A(net40),
    .B(_05698_),
    .Y(_05729_));
 sky130_fd_sc_hd__o21ai_0 _16616_ (.A1(_05206_),
    .A2(_05698_),
    .B1(_05729_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _16617_ (.A(net39),
    .B(_05698_),
    .Y(_05730_));
 sky130_fd_sc_hd__o21ai_0 _16618_ (.A1(_05214_),
    .A2(_05698_),
    .B1(_05730_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _16619_ (.A(net38),
    .B(_05698_),
    .Y(_05731_));
 sky130_fd_sc_hd__o21ai_0 _16620_ (.A1(_05224_),
    .A2(_05698_),
    .B1(_05731_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _16621_ (.A(net37),
    .B(_05698_),
    .Y(_05732_));
 sky130_fd_sc_hd__o21ai_0 _16622_ (.A1(_05236_),
    .A2(_05698_),
    .B1(_05732_),
    .Y(_00468_));
 sky130_fd_sc_hd__nand2_1 _16623_ (.A(net36),
    .B(_05698_),
    .Y(_05733_));
 sky130_fd_sc_hd__o21ai_0 _16624_ (.A1(_05243_),
    .A2(_05698_),
    .B1(_05733_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _16625_ (.A(net35),
    .B(_05698_),
    .Y(_05734_));
 sky130_fd_sc_hd__o21ai_0 _16626_ (.A1(_05251_),
    .A2(_05698_),
    .B1(_05734_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _16627_ (.A(net33),
    .B(_05698_),
    .Y(_05735_));
 sky130_fd_sc_hd__o21ai_0 _16628_ (.A1(_05260_),
    .A2(_05698_),
    .B1(_05735_),
    .Y(_00472_));
 sky130_fd_sc_hd__nand2_1 _16629_ (.A(net32),
    .B(_05698_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21ai_0 _16630_ (.A1(_05310_),
    .A2(_05698_),
    .B1(_05736_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2b_4 _16631_ (.A(net762),
    .B_N(_13705_),
    .Y(_05737_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1264 ();
 sky130_fd_sc_hd__nand2_8 _16633_ (.A(_09959_),
    .B(_05737_),
    .Y(_05739_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1262 ();
 sky130_fd_sc_hd__nand2_1 _16636_ (.A(net102),
    .B(_05739_),
    .Y(_05742_));
 sky130_fd_sc_hd__o21ai_0 _16637_ (.A1(_05317_),
    .A2(_05739_),
    .B1(_05742_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _16638_ (.A(net101),
    .B(_05739_),
    .Y(_05743_));
 sky130_fd_sc_hd__o21ai_0 _16639_ (.A1(_05321_),
    .A2(_05739_),
    .B1(_05743_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _16640_ (.A(net99),
    .B(_05739_),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ai_0 _16641_ (.A1(_05324_),
    .A2(_05739_),
    .B1(_05744_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _16642_ (.A(net98),
    .B(_05739_),
    .Y(_05745_));
 sky130_fd_sc_hd__o21ai_0 _16643_ (.A1(_05330_),
    .A2(_05739_),
    .B1(_05745_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _16644_ (.A(net97),
    .B(_05739_),
    .Y(_05746_));
 sky130_fd_sc_hd__o21ai_0 _16645_ (.A1(_05338_),
    .A2(_05739_),
    .B1(_05746_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _16646_ (.A(net96),
    .B(_05739_),
    .Y(_05747_));
 sky130_fd_sc_hd__o21ai_0 _16647_ (.A1(_05347_),
    .A2(_05739_),
    .B1(_05747_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _16648_ (.A(net95),
    .B(_05739_),
    .Y(_05748_));
 sky130_fd_sc_hd__o21ai_0 _16649_ (.A1(_05354_),
    .A2(_05739_),
    .B1(_05748_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _16650_ (.A(net94),
    .B(_05739_),
    .Y(_05749_));
 sky130_fd_sc_hd__o21ai_0 _16651_ (.A1(_05360_),
    .A2(_05739_),
    .B1(_05749_),
    .Y(_00510_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1261 ();
 sky130_fd_sc_hd__nand2_1 _16653_ (.A(net93),
    .B(_05739_),
    .Y(_05751_));
 sky130_fd_sc_hd__o21ai_0 _16654_ (.A1(_05371_),
    .A2(_05739_),
    .B1(_05751_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _16655_ (.A(net92),
    .B(_05739_),
    .Y(_05752_));
 sky130_fd_sc_hd__o21ai_0 _16656_ (.A1(_05380_),
    .A2(_05739_),
    .B1(_05752_),
    .Y(_00512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1260 ();
 sky130_fd_sc_hd__nand2_1 _16658_ (.A(net91),
    .B(_05739_),
    .Y(_05754_));
 sky130_fd_sc_hd__o21ai_0 _16659_ (.A1(_05388_),
    .A2(_05739_),
    .B1(_05754_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _16660_ (.A(net90),
    .B(_05739_),
    .Y(_05755_));
 sky130_fd_sc_hd__o21ai_0 _16661_ (.A1(_05402_),
    .A2(_05739_),
    .B1(_05755_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _16662_ (.A(net88),
    .B(_05739_),
    .Y(_05756_));
 sky130_fd_sc_hd__o21ai_0 _16663_ (.A1(_05412_),
    .A2(_05739_),
    .B1(_05756_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _16664_ (.A(net87),
    .B(_05739_),
    .Y(_05757_));
 sky130_fd_sc_hd__o21ai_0 _16665_ (.A1(_05419_),
    .A2(_05739_),
    .B1(_05757_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _16666_ (.A(net86),
    .B(_05739_),
    .Y(_05758_));
 sky130_fd_sc_hd__o21ai_0 _16667_ (.A1(_05426_),
    .A2(_05739_),
    .B1(_05758_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _16668_ (.A(net85),
    .B(_05739_),
    .Y(_05759_));
 sky130_fd_sc_hd__o21ai_0 _16669_ (.A1(_05438_),
    .A2(_05739_),
    .B1(_05759_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _16670_ (.A(net84),
    .B(_05739_),
    .Y(_05760_));
 sky130_fd_sc_hd__o21ai_0 _16671_ (.A1(_05447_),
    .A2(_05739_),
    .B1(_05760_),
    .Y(_00488_));
 sky130_fd_sc_hd__nand2_1 _16672_ (.A(net83),
    .B(_05739_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_0 _16673_ (.A1(_05453_),
    .A2(_05739_),
    .B1(_05761_),
    .Y(_00489_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1259 ();
 sky130_fd_sc_hd__nand2_1 _16675_ (.A(net82),
    .B(_05739_),
    .Y(_05763_));
 sky130_fd_sc_hd__o21ai_0 _16676_ (.A1(_05465_),
    .A2(_05739_),
    .B1(_05763_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_1 _16677_ (.A(net81),
    .B(_05739_),
    .Y(_05764_));
 sky130_fd_sc_hd__o21ai_0 _16678_ (.A1(_05480_),
    .A2(_05739_),
    .B1(_05764_),
    .Y(_00491_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1258 ();
 sky130_fd_sc_hd__nand2_1 _16680_ (.A(net80),
    .B(_05739_),
    .Y(_05766_));
 sky130_fd_sc_hd__o21ai_0 _16681_ (.A1(_05488_),
    .A2(_05739_),
    .B1(_05766_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _16682_ (.A(net79),
    .B(_05739_),
    .Y(_05767_));
 sky130_fd_sc_hd__o21ai_0 _16683_ (.A1(_05498_),
    .A2(_05739_),
    .B1(_05767_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _16684_ (.A(net77),
    .B(_05739_),
    .Y(_05768_));
 sky130_fd_sc_hd__o21ai_0 _16685_ (.A1(_05509_),
    .A2(_05739_),
    .B1(_05768_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand2_1 _16686_ (.A(net76),
    .B(_05739_),
    .Y(_05769_));
 sky130_fd_sc_hd__o21ai_0 _16687_ (.A1(_05515_),
    .A2(_05739_),
    .B1(_05769_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _16688_ (.A(net75),
    .B(_05739_),
    .Y(_05770_));
 sky130_fd_sc_hd__o21ai_0 _16689_ (.A1(_05523_),
    .A2(_05739_),
    .B1(_05770_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _16690_ (.A(net74),
    .B(_05739_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_0 _16691_ (.A1(_05535_),
    .A2(_05739_),
    .B1(_05771_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _16692_ (.A(net73),
    .B(_05739_),
    .Y(_05772_));
 sky130_fd_sc_hd__o21ai_0 _16693_ (.A1(_05542_),
    .A2(_05739_),
    .B1(_05772_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _16694_ (.A(net72),
    .B(_05739_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21ai_0 _16695_ (.A1(_05551_),
    .A2(_05739_),
    .B1(_05773_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _16696_ (.A(net71),
    .B(_05739_),
    .Y(_05774_));
 sky130_fd_sc_hd__o21ai_0 _16697_ (.A1(_05559_),
    .A2(_05739_),
    .B1(_05774_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _16698_ (.A(net70),
    .B(_05739_),
    .Y(_05775_));
 sky130_fd_sc_hd__o21ai_0 _16699_ (.A1(_05567_),
    .A2(_05739_),
    .B1(_05775_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2_1 _16700_ (.A(net69),
    .B(_05739_),
    .Y(_05776_));
 sky130_fd_sc_hd__o21ai_0 _16701_ (.A1(_05573_),
    .A2(_05739_),
    .B1(_05776_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _16702_ (.A(net68),
    .B(_05739_),
    .Y(_05777_));
 sky130_fd_sc_hd__o21ai_0 _16703_ (.A1(_05611_),
    .A2(_05739_),
    .B1(_05777_),
    .Y(_00505_));
 sky130_fd_sc_hd__nor2b_4 _16704_ (.A(net762),
    .B_N(_13701_),
    .Y(_05778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1257 ();
 sky130_fd_sc_hd__nand2_8 _16706_ (.A(_09897_),
    .B(_05778_),
    .Y(_05780_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1255 ();
 sky130_fd_sc_hd__nand2_1 _16709_ (.A(net138),
    .B(_05780_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21ai_0 _16710_ (.A1(_04988_),
    .A2(_05780_),
    .B1(_05783_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _16711_ (.A(net137),
    .B(_05780_),
    .Y(_05784_));
 sky130_fd_sc_hd__o21ai_0 _16712_ (.A1(_04992_),
    .A2(_05780_),
    .B1(_05784_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _16713_ (.A(net136),
    .B(_05780_),
    .Y(_05785_));
 sky130_fd_sc_hd__o21ai_0 _16714_ (.A1(_04995_),
    .A2(_05780_),
    .B1(_05785_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _16715_ (.A(net135),
    .B(_05780_),
    .Y(_05786_));
 sky130_fd_sc_hd__o21ai_0 _16716_ (.A1(_05003_),
    .A2(_05780_),
    .B1(_05786_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _16717_ (.A(net133),
    .B(_05780_),
    .Y(_05787_));
 sky130_fd_sc_hd__o21ai_0 _16718_ (.A1(_05012_),
    .A2(_05780_),
    .B1(_05787_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand2_1 _16719_ (.A(net132),
    .B(_05780_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21ai_0 _16720_ (.A1(_05021_),
    .A2(_05780_),
    .B1(_05788_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _16721_ (.A(net131),
    .B(_05780_),
    .Y(_05789_));
 sky130_fd_sc_hd__o21ai_0 _16722_ (.A1(_05032_),
    .A2(_05780_),
    .B1(_05789_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _16723_ (.A(net130),
    .B(_05780_),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ai_0 _16724_ (.A1(_05039_),
    .A2(_05780_),
    .B1(_05790_),
    .Y(_00542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1254 ();
 sky130_fd_sc_hd__nand2_1 _16726_ (.A(net129),
    .B(_05780_),
    .Y(_05792_));
 sky130_fd_sc_hd__o21ai_0 _16727_ (.A1(_05048_),
    .A2(_05780_),
    .B1(_05792_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _16728_ (.A(net128),
    .B(_05780_),
    .Y(_05793_));
 sky130_fd_sc_hd__o21ai_0 _16729_ (.A1(_05055_),
    .A2(_05780_),
    .B1(_05793_),
    .Y(_00544_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1253 ();
 sky130_fd_sc_hd__nand2_1 _16731_ (.A(net127),
    .B(_05780_),
    .Y(_05795_));
 sky130_fd_sc_hd__o21ai_0 _16732_ (.A1(_05062_),
    .A2(_05780_),
    .B1(_05795_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _16733_ (.A(net126),
    .B(_05780_),
    .Y(_05796_));
 sky130_fd_sc_hd__o21ai_0 _16734_ (.A1(_05077_),
    .A2(_05780_),
    .B1(_05796_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _16735_ (.A(net125),
    .B(_05780_),
    .Y(_05797_));
 sky130_fd_sc_hd__o21ai_0 _16736_ (.A1(_05087_),
    .A2(_05780_),
    .B1(_05797_),
    .Y(_00516_));
 sky130_fd_sc_hd__nand2_1 _16737_ (.A(net124),
    .B(_05780_),
    .Y(_05798_));
 sky130_fd_sc_hd__o21ai_0 _16738_ (.A1(_05095_),
    .A2(_05780_),
    .B1(_05798_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _16739_ (.A(net122),
    .B(_05780_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ai_0 _16740_ (.A1(_05102_),
    .A2(_05780_),
    .B1(_05799_),
    .Y(_00518_));
 sky130_fd_sc_hd__nand2_1 _16741_ (.A(net121),
    .B(_05780_),
    .Y(_05800_));
 sky130_fd_sc_hd__o21ai_0 _16742_ (.A1(_05112_),
    .A2(_05780_),
    .B1(_05800_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _16743_ (.A(net120),
    .B(_05780_),
    .Y(_05801_));
 sky130_fd_sc_hd__o21ai_0 _16744_ (.A1(_05121_),
    .A2(_05780_),
    .B1(_05801_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _16745_ (.A(net119),
    .B(_05780_),
    .Y(_05802_));
 sky130_fd_sc_hd__o21ai_0 _16746_ (.A1(_05128_),
    .A2(_05780_),
    .B1(_05802_),
    .Y(_00521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1252 ();
 sky130_fd_sc_hd__nand2_1 _16748_ (.A(net118),
    .B(_05780_),
    .Y(_05804_));
 sky130_fd_sc_hd__o21ai_0 _16749_ (.A1(_05137_),
    .A2(_05780_),
    .B1(_05804_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_1 _16750_ (.A(net117),
    .B(_05780_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_0 _16751_ (.A1(_05154_),
    .A2(_05780_),
    .B1(_05805_),
    .Y(_00523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1251 ();
 sky130_fd_sc_hd__nand2_1 _16753_ (.A(net116),
    .B(_05780_),
    .Y(_05807_));
 sky130_fd_sc_hd__o21ai_0 _16754_ (.A1(_05167_),
    .A2(_05780_),
    .B1(_05807_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _16755_ (.A(net115),
    .B(_05780_),
    .Y(_05808_));
 sky130_fd_sc_hd__o21ai_0 _16756_ (.A1(_05175_),
    .A2(_05780_),
    .B1(_05808_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _16757_ (.A(net114),
    .B(_05780_),
    .Y(_05809_));
 sky130_fd_sc_hd__o21ai_0 _16758_ (.A1(_05184_),
    .A2(_05780_),
    .B1(_05809_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _16759_ (.A(net113),
    .B(_05780_),
    .Y(_05810_));
 sky130_fd_sc_hd__o21ai_0 _16760_ (.A1(_05196_),
    .A2(_05780_),
    .B1(_05810_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _16761_ (.A(net110),
    .B(_05780_),
    .Y(_05811_));
 sky130_fd_sc_hd__o21ai_0 _16762_ (.A1(_05206_),
    .A2(_05780_),
    .B1(_05811_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _16763_ (.A(net109),
    .B(_05780_),
    .Y(_05812_));
 sky130_fd_sc_hd__o21ai_0 _16764_ (.A1(_05214_),
    .A2(_05780_),
    .B1(_05812_),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _16765_ (.A(net108),
    .B(_05780_),
    .Y(_05813_));
 sky130_fd_sc_hd__o21ai_0 _16766_ (.A1(_05224_),
    .A2(_05780_),
    .B1(_05813_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _16767_ (.A(net107),
    .B(_05780_),
    .Y(_05814_));
 sky130_fd_sc_hd__o21ai_0 _16768_ (.A1(_05236_),
    .A2(_05780_),
    .B1(_05814_),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _16769_ (.A(net106),
    .B(_05780_),
    .Y(_05815_));
 sky130_fd_sc_hd__o21ai_0 _16770_ (.A1(_05243_),
    .A2(_05780_),
    .B1(_05815_),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2_1 _16771_ (.A(net105),
    .B(_05780_),
    .Y(_05816_));
 sky130_fd_sc_hd__o21ai_0 _16772_ (.A1(_05251_),
    .A2(_05780_),
    .B1(_05816_),
    .Y(_00534_));
 sky130_fd_sc_hd__nand2_1 _16773_ (.A(net104),
    .B(_05780_),
    .Y(_05817_));
 sky130_fd_sc_hd__o21ai_0 _16774_ (.A1(_05260_),
    .A2(_05780_),
    .B1(_05817_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _16775_ (.A(net103),
    .B(_05780_),
    .Y(_05818_));
 sky130_fd_sc_hd__o21ai_0 _16776_ (.A1(_05310_),
    .A2(_05780_),
    .B1(_05818_),
    .Y(_00537_));
 sky130_fd_sc_hd__nor2b_2 _16777_ (.A(\count_2[5] ),
    .B_N(_13709_),
    .Y(_05819_));
 sky130_fd_sc_hd__nor3_4 _16778_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(net762),
    .Y(_05820_));
 sky130_fd_sc_hd__nand2_8 _16779_ (.A(_05819_),
    .B(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1249 ();
 sky130_fd_sc_hd__nand2_1 _16782_ (.A(net173),
    .B(_05821_),
    .Y(_05824_));
 sky130_fd_sc_hd__o21ai_0 _16783_ (.A1(_05317_),
    .A2(_05821_),
    .B1(_05824_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _16784_ (.A(net172),
    .B(_05821_),
    .Y(_05825_));
 sky130_fd_sc_hd__o21ai_0 _16785_ (.A1(_05321_),
    .A2(_05821_),
    .B1(_05825_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand2_1 _16786_ (.A(net171),
    .B(_05821_),
    .Y(_05826_));
 sky130_fd_sc_hd__o21ai_0 _16787_ (.A1(_05324_),
    .A2(_05821_),
    .B1(_05826_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand2_1 _16788_ (.A(net170),
    .B(_05821_),
    .Y(_05827_));
 sky130_fd_sc_hd__o21ai_0 _16789_ (.A1(_05330_),
    .A2(_05821_),
    .B1(_05827_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _16790_ (.A(net169),
    .B(_05821_),
    .Y(_05828_));
 sky130_fd_sc_hd__o21ai_0 _16791_ (.A1(_05338_),
    .A2(_05821_),
    .B1(_05828_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _16792_ (.A(net168),
    .B(_05821_),
    .Y(_05829_));
 sky130_fd_sc_hd__o21ai_0 _16793_ (.A1(_05347_),
    .A2(_05821_),
    .B1(_05829_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _16794_ (.A(net166),
    .B(_05821_),
    .Y(_05830_));
 sky130_fd_sc_hd__o21ai_0 _16795_ (.A1(_05354_),
    .A2(_05821_),
    .B1(_05830_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _16796_ (.A(net165),
    .B(_05821_),
    .Y(_05831_));
 sky130_fd_sc_hd__o21ai_0 _16797_ (.A1(_05360_),
    .A2(_05821_),
    .B1(_05831_),
    .Y(_00574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1248 ();
 sky130_fd_sc_hd__nand2_1 _16799_ (.A(net164),
    .B(_05821_),
    .Y(_05833_));
 sky130_fd_sc_hd__o21ai_0 _16800_ (.A1(_05371_),
    .A2(_05821_),
    .B1(_05833_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _16801_ (.A(net163),
    .B(_05821_),
    .Y(_05834_));
 sky130_fd_sc_hd__o21ai_0 _16802_ (.A1(_05380_),
    .A2(_05821_),
    .B1(_05834_),
    .Y(_00576_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1247 ();
 sky130_fd_sc_hd__nand2_1 _16804_ (.A(net162),
    .B(_05821_),
    .Y(_05836_));
 sky130_fd_sc_hd__o21ai_0 _16805_ (.A1(_05388_),
    .A2(_05821_),
    .B1(_05836_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(net161),
    .B(_05821_),
    .Y(_05837_));
 sky130_fd_sc_hd__o21ai_0 _16807_ (.A1(_05402_),
    .A2(_05821_),
    .B1(_05837_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _16808_ (.A(net160),
    .B(_05821_),
    .Y(_05838_));
 sky130_fd_sc_hd__o21ai_0 _16809_ (.A1(_05412_),
    .A2(_05821_),
    .B1(_05838_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _16810_ (.A(net159),
    .B(_05821_),
    .Y(_05839_));
 sky130_fd_sc_hd__o21ai_0 _16811_ (.A1(_05419_),
    .A2(_05821_),
    .B1(_05839_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _16812_ (.A(net158),
    .B(_05821_),
    .Y(_05840_));
 sky130_fd_sc_hd__o21ai_0 _16813_ (.A1(_05426_),
    .A2(_05821_),
    .B1(_05840_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _16814_ (.A(net157),
    .B(_05821_),
    .Y(_05841_));
 sky130_fd_sc_hd__o21ai_0 _16815_ (.A1(_05438_),
    .A2(_05821_),
    .B1(_05841_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _16816_ (.A(net155),
    .B(_05821_),
    .Y(_05842_));
 sky130_fd_sc_hd__o21ai_0 _16817_ (.A1(_05447_),
    .A2(_05821_),
    .B1(_05842_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _16818_ (.A(net154),
    .B(_05821_),
    .Y(_05843_));
 sky130_fd_sc_hd__o21ai_0 _16819_ (.A1(_05453_),
    .A2(_05821_),
    .B1(_05843_),
    .Y(_00553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1246 ();
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(net153),
    .B(_05821_),
    .Y(_05845_));
 sky130_fd_sc_hd__o21ai_0 _16822_ (.A1(_05465_),
    .A2(_05821_),
    .B1(_05845_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _16823_ (.A(net152),
    .B(_05821_),
    .Y(_05846_));
 sky130_fd_sc_hd__o21ai_0 _16824_ (.A1(_05480_),
    .A2(_05821_),
    .B1(_05846_),
    .Y(_00555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1245 ();
 sky130_fd_sc_hd__nand2_1 _16826_ (.A(net151),
    .B(_05821_),
    .Y(_05848_));
 sky130_fd_sc_hd__o21ai_0 _16827_ (.A1(_05488_),
    .A2(_05821_),
    .B1(_05848_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _16828_ (.A(net150),
    .B(_05821_),
    .Y(_05849_));
 sky130_fd_sc_hd__o21ai_0 _16829_ (.A1(_05498_),
    .A2(_05821_),
    .B1(_05849_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_1 _16830_ (.A(net149),
    .B(_05821_),
    .Y(_05850_));
 sky130_fd_sc_hd__o21ai_0 _16831_ (.A1(_05509_),
    .A2(_05821_),
    .B1(_05850_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _16832_ (.A(net148),
    .B(_05821_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_0 _16833_ (.A1(_05515_),
    .A2(_05821_),
    .B1(_05851_),
    .Y(_00560_));
 sky130_fd_sc_hd__nand2_1 _16834_ (.A(net147),
    .B(_05821_),
    .Y(_05852_));
 sky130_fd_sc_hd__o21ai_0 _16835_ (.A1(_05523_),
    .A2(_05821_),
    .B1(_05852_),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_1 _16836_ (.A(net146),
    .B(_05821_),
    .Y(_05853_));
 sky130_fd_sc_hd__o21ai_0 _16837_ (.A1(_05535_),
    .A2(_05821_),
    .B1(_05853_),
    .Y(_00562_));
 sky130_fd_sc_hd__nand2_1 _16838_ (.A(net144),
    .B(_05821_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_0 _16839_ (.A1(_05542_),
    .A2(_05821_),
    .B1(_05854_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _16840_ (.A(net143),
    .B(_05821_),
    .Y(_05855_));
 sky130_fd_sc_hd__o21ai_0 _16841_ (.A1(_05551_),
    .A2(_05821_),
    .B1(_05855_),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_1 _16842_ (.A(net142),
    .B(_05821_),
    .Y(_05856_));
 sky130_fd_sc_hd__o21ai_0 _16843_ (.A1(_05559_),
    .A2(_05821_),
    .B1(_05856_),
    .Y(_00565_));
 sky130_fd_sc_hd__nand2_1 _16844_ (.A(net141),
    .B(_05821_),
    .Y(_05857_));
 sky130_fd_sc_hd__o21ai_0 _16845_ (.A1(_05567_),
    .A2(_05821_),
    .B1(_05857_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _16846_ (.A(net140),
    .B(_05821_),
    .Y(_05858_));
 sky130_fd_sc_hd__o21ai_0 _16847_ (.A1(_05573_),
    .A2(_05821_),
    .B1(_05858_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _16848_ (.A(net139),
    .B(_05821_),
    .Y(_05859_));
 sky130_fd_sc_hd__o21ai_0 _16849_ (.A1(_05611_),
    .A2(_05821_),
    .B1(_05859_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_8 _16850_ (.A(_09901_),
    .B(_04982_),
    .Y(_05860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1243 ();
 sky130_fd_sc_hd__nand2_1 _16853_ (.A(net208),
    .B(_05860_),
    .Y(_05863_));
 sky130_fd_sc_hd__o21ai_0 _16854_ (.A1(_04988_),
    .A2(_05860_),
    .B1(_05863_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _16855_ (.A(net207),
    .B(_05860_),
    .Y(_05864_));
 sky130_fd_sc_hd__o21ai_0 _16856_ (.A1(_04992_),
    .A2(_05860_),
    .B1(_05864_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(net206),
    .B(_05860_),
    .Y(_05865_));
 sky130_fd_sc_hd__o21ai_0 _16858_ (.A1(_04995_),
    .A2(_05860_),
    .B1(_05865_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _16859_ (.A(net205),
    .B(_05860_),
    .Y(_05866_));
 sky130_fd_sc_hd__o21ai_0 _16860_ (.A1(_05003_),
    .A2(_05860_),
    .B1(_05866_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _16861_ (.A(net204),
    .B(_05860_),
    .Y(_05867_));
 sky130_fd_sc_hd__o21ai_0 _16862_ (.A1(_05012_),
    .A2(_05860_),
    .B1(_05867_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _16863_ (.A(net203),
    .B(_05860_),
    .Y(_05868_));
 sky130_fd_sc_hd__o21ai_0 _16864_ (.A1(_05021_),
    .A2(_05860_),
    .B1(_05868_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _16865_ (.A(net202),
    .B(_05860_),
    .Y(_05869_));
 sky130_fd_sc_hd__o21ai_0 _16866_ (.A1(_05032_),
    .A2(_05860_),
    .B1(_05869_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(net201),
    .B(_05860_),
    .Y(_05870_));
 sky130_fd_sc_hd__o21ai_0 _16868_ (.A1(_05039_),
    .A2(_05860_),
    .B1(_05870_),
    .Y(_00606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1242 ();
 sky130_fd_sc_hd__nand2_1 _16870_ (.A(net199),
    .B(_05860_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21ai_0 _16871_ (.A1(_05048_),
    .A2(_05860_),
    .B1(_05872_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _16872_ (.A(net198),
    .B(_05860_),
    .Y(_05873_));
 sky130_fd_sc_hd__o21ai_0 _16873_ (.A1(_05055_),
    .A2(_05860_),
    .B1(_05873_),
    .Y(_00608_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1241 ();
 sky130_fd_sc_hd__nand2_1 _16875_ (.A(net197),
    .B(_05860_),
    .Y(_05875_));
 sky130_fd_sc_hd__o21ai_0 _16876_ (.A1(_05062_),
    .A2(_05860_),
    .B1(_05875_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _16877_ (.A(net196),
    .B(_05860_),
    .Y(_05876_));
 sky130_fd_sc_hd__o21ai_0 _16878_ (.A1(_05077_),
    .A2(_05860_),
    .B1(_05876_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _16879_ (.A(net195),
    .B(_05860_),
    .Y(_05877_));
 sky130_fd_sc_hd__o21ai_0 _16880_ (.A1(_05087_),
    .A2(_05860_),
    .B1(_05877_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_1 _16881_ (.A(net194),
    .B(_05860_),
    .Y(_05878_));
 sky130_fd_sc_hd__o21ai_0 _16882_ (.A1(_05095_),
    .A2(_05860_),
    .B1(_05878_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_1 _16883_ (.A(net193),
    .B(_05860_),
    .Y(_05879_));
 sky130_fd_sc_hd__o21ai_0 _16884_ (.A1(_05102_),
    .A2(_05860_),
    .B1(_05879_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _16885_ (.A(net192),
    .B(_05860_),
    .Y(_05880_));
 sky130_fd_sc_hd__o21ai_0 _16886_ (.A1(_05112_),
    .A2(_05860_),
    .B1(_05880_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _16887_ (.A(net191),
    .B(_05860_),
    .Y(_05881_));
 sky130_fd_sc_hd__o21ai_0 _16888_ (.A1(_05121_),
    .A2(_05860_),
    .B1(_05881_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _16889_ (.A(net190),
    .B(_05860_),
    .Y(_05882_));
 sky130_fd_sc_hd__o21ai_0 _16890_ (.A1(_05128_),
    .A2(_05860_),
    .B1(_05882_),
    .Y(_00585_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1240 ();
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(net188),
    .B(_05860_),
    .Y(_05884_));
 sky130_fd_sc_hd__o21ai_0 _16893_ (.A1(_05137_),
    .A2(_05860_),
    .B1(_05884_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _16894_ (.A(net187),
    .B(_05860_),
    .Y(_05885_));
 sky130_fd_sc_hd__o21ai_0 _16895_ (.A1(_05154_),
    .A2(_05860_),
    .B1(_05885_),
    .Y(_00587_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1239 ();
 sky130_fd_sc_hd__nand2_1 _16897_ (.A(net186),
    .B(_05860_),
    .Y(_05887_));
 sky130_fd_sc_hd__o21ai_0 _16898_ (.A1(_05167_),
    .A2(_05860_),
    .B1(_05887_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _16899_ (.A(net185),
    .B(_05860_),
    .Y(_05888_));
 sky130_fd_sc_hd__o21ai_0 _16900_ (.A1(_05175_),
    .A2(_05860_),
    .B1(_05888_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _16901_ (.A(net184),
    .B(_05860_),
    .Y(_05889_));
 sky130_fd_sc_hd__o21ai_0 _16902_ (.A1(_05184_),
    .A2(_05860_),
    .B1(_05889_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand2_1 _16903_ (.A(net183),
    .B(_05860_),
    .Y(_05890_));
 sky130_fd_sc_hd__o21ai_0 _16904_ (.A1(_05196_),
    .A2(_05860_),
    .B1(_05890_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _16905_ (.A(net182),
    .B(_05860_),
    .Y(_05891_));
 sky130_fd_sc_hd__o21ai_0 _16906_ (.A1(_05206_),
    .A2(_05860_),
    .B1(_05891_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _16907_ (.A(net181),
    .B(_05860_),
    .Y(_05892_));
 sky130_fd_sc_hd__o21ai_0 _16908_ (.A1(_05214_),
    .A2(_05860_),
    .B1(_05892_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _16909_ (.A(net180),
    .B(_05860_),
    .Y(_05893_));
 sky130_fd_sc_hd__o21ai_0 _16910_ (.A1(_05224_),
    .A2(_05860_),
    .B1(_05893_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _16911_ (.A(net179),
    .B(_05860_),
    .Y(_05894_));
 sky130_fd_sc_hd__o21ai_0 _16912_ (.A1(_05236_),
    .A2(_05860_),
    .B1(_05894_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _16913_ (.A(net177),
    .B(_05860_),
    .Y(_05895_));
 sky130_fd_sc_hd__o21ai_0 _16914_ (.A1(_05243_),
    .A2(_05860_),
    .B1(_05895_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _16915_ (.A(net176),
    .B(_05860_),
    .Y(_05896_));
 sky130_fd_sc_hd__o21ai_0 _16916_ (.A1(_05251_),
    .A2(_05860_),
    .B1(_05896_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(net175),
    .B(_05860_),
    .Y(_05897_));
 sky130_fd_sc_hd__o21ai_0 _16918_ (.A1(_05260_),
    .A2(_05860_),
    .B1(_05897_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _16919_ (.A(net174),
    .B(_05860_),
    .Y(_05898_));
 sky130_fd_sc_hd__o21ai_0 _16920_ (.A1(_05310_),
    .A2(_05860_),
    .B1(_05898_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_8 _16921_ (.A(_09946_),
    .B(_05313_),
    .Y(_05899_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1237 ();
 sky130_fd_sc_hd__nand2_1 _16924_ (.A(net244),
    .B(_05899_),
    .Y(_05902_));
 sky130_fd_sc_hd__o21ai_0 _16925_ (.A1(_05317_),
    .A2(_05899_),
    .B1(_05902_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _16926_ (.A(net243),
    .B(_05899_),
    .Y(_05903_));
 sky130_fd_sc_hd__o21ai_0 _16927_ (.A1(_05321_),
    .A2(_05899_),
    .B1(_05903_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _16928_ (.A(net242),
    .B(_05899_),
    .Y(_05904_));
 sky130_fd_sc_hd__o21ai_0 _16929_ (.A1(_05324_),
    .A2(_05899_),
    .B1(_05904_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _16930_ (.A(net241),
    .B(_05899_),
    .Y(_05905_));
 sky130_fd_sc_hd__o21ai_0 _16931_ (.A1(_05330_),
    .A2(_05899_),
    .B1(_05905_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _16932_ (.A(net240),
    .B(_05899_),
    .Y(_05906_));
 sky130_fd_sc_hd__o21ai_0 _16933_ (.A1(_05338_),
    .A2(_05899_),
    .B1(_05906_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _16934_ (.A(net239),
    .B(_05899_),
    .Y(_05907_));
 sky130_fd_sc_hd__o21ai_0 _16935_ (.A1(_05347_),
    .A2(_05899_),
    .B1(_05907_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _16936_ (.A(net238),
    .B(_05899_),
    .Y(_05908_));
 sky130_fd_sc_hd__o21ai_0 _16937_ (.A1(_05354_),
    .A2(_05899_),
    .B1(_05908_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _16938_ (.A(net237),
    .B(_05899_),
    .Y(_05909_));
 sky130_fd_sc_hd__o21ai_0 _16939_ (.A1(_05360_),
    .A2(_05899_),
    .B1(_05909_),
    .Y(_00638_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1236 ();
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(net236),
    .B(_05899_),
    .Y(_05911_));
 sky130_fd_sc_hd__o21ai_0 _16942_ (.A1(_05371_),
    .A2(_05899_),
    .B1(_05911_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2_1 _16943_ (.A(net235),
    .B(_05899_),
    .Y(_05912_));
 sky130_fd_sc_hd__o21ai_0 _16944_ (.A1(_05380_),
    .A2(_05899_),
    .B1(_05912_),
    .Y(_00640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1235 ();
 sky130_fd_sc_hd__nand2_1 _16946_ (.A(net233),
    .B(_05899_),
    .Y(_05914_));
 sky130_fd_sc_hd__o21ai_0 _16947_ (.A1(_05388_),
    .A2(_05899_),
    .B1(_05914_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _16948_ (.A(net232),
    .B(_05899_),
    .Y(_05915_));
 sky130_fd_sc_hd__o21ai_0 _16949_ (.A1(_05402_),
    .A2(_05899_),
    .B1(_05915_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _16950_ (.A(net231),
    .B(_05899_),
    .Y(_05916_));
 sky130_fd_sc_hd__o21ai_0 _16951_ (.A1(_05412_),
    .A2(_05899_),
    .B1(_05916_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _16952_ (.A(net230),
    .B(_05899_),
    .Y(_05917_));
 sky130_fd_sc_hd__o21ai_0 _16953_ (.A1(_05419_),
    .A2(_05899_),
    .B1(_05917_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _16954_ (.A(net229),
    .B(_05899_),
    .Y(_05918_));
 sky130_fd_sc_hd__o21ai_0 _16955_ (.A1(_05426_),
    .A2(_05899_),
    .B1(_05918_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _16956_ (.A(net228),
    .B(_05899_),
    .Y(_05919_));
 sky130_fd_sc_hd__o21ai_0 _16957_ (.A1(_05438_),
    .A2(_05899_),
    .B1(_05919_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _16958_ (.A(net227),
    .B(_05899_),
    .Y(_05920_));
 sky130_fd_sc_hd__o21ai_0 _16959_ (.A1(_05447_),
    .A2(_05899_),
    .B1(_05920_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _16960_ (.A(net226),
    .B(_05899_),
    .Y(_05921_));
 sky130_fd_sc_hd__o21ai_0 _16961_ (.A1(_05453_),
    .A2(_05899_),
    .B1(_05921_),
    .Y(_00617_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1234 ();
 sky130_fd_sc_hd__nand2_1 _16963_ (.A(net225),
    .B(_05899_),
    .Y(_05923_));
 sky130_fd_sc_hd__o21ai_0 _16964_ (.A1(_05465_),
    .A2(_05899_),
    .B1(_05923_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand2_1 _16965_ (.A(net224),
    .B(_05899_),
    .Y(_05924_));
 sky130_fd_sc_hd__o21ai_0 _16966_ (.A1(_05480_),
    .A2(_05899_),
    .B1(_05924_),
    .Y(_00619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1233 ();
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(net221),
    .B(_05899_),
    .Y(_05926_));
 sky130_fd_sc_hd__o21ai_0 _16969_ (.A1(_05488_),
    .A2(_05899_),
    .B1(_05926_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(net220),
    .B(_05899_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21ai_0 _16971_ (.A1(_05498_),
    .A2(_05899_),
    .B1(_05927_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _16972_ (.A(net219),
    .B(_05899_),
    .Y(_05928_));
 sky130_fd_sc_hd__o21ai_0 _16973_ (.A1(_05509_),
    .A2(_05899_),
    .B1(_05928_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(net218),
    .B(_05899_),
    .Y(_05929_));
 sky130_fd_sc_hd__o21ai_0 _16975_ (.A1(_05515_),
    .A2(_05899_),
    .B1(_05929_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _16976_ (.A(net217),
    .B(_05899_),
    .Y(_05930_));
 sky130_fd_sc_hd__o21ai_0 _16977_ (.A1(_05523_),
    .A2(_05899_),
    .B1(_05930_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(net216),
    .B(_05899_),
    .Y(_05931_));
 sky130_fd_sc_hd__o21ai_0 _16979_ (.A1(_05535_),
    .A2(_05899_),
    .B1(_05931_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _16980_ (.A(net215),
    .B(_05899_),
    .Y(_05932_));
 sky130_fd_sc_hd__o21ai_0 _16981_ (.A1(_05542_),
    .A2(_05899_),
    .B1(_05932_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _16982_ (.A(net214),
    .B(_05899_),
    .Y(_05933_));
 sky130_fd_sc_hd__o21ai_0 _16983_ (.A1(_05551_),
    .A2(_05899_),
    .B1(_05933_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(net213),
    .B(_05899_),
    .Y(_05934_));
 sky130_fd_sc_hd__o21ai_0 _16985_ (.A1(_05559_),
    .A2(_05899_),
    .B1(_05934_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _16986_ (.A(net212),
    .B(_05899_),
    .Y(_05935_));
 sky130_fd_sc_hd__o21ai_0 _16987_ (.A1(_05567_),
    .A2(_05899_),
    .B1(_05935_),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _16988_ (.A(net210),
    .B(_05899_),
    .Y(_05936_));
 sky130_fd_sc_hd__o21ai_0 _16989_ (.A1(_05573_),
    .A2(_05899_),
    .B1(_05936_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _16990_ (.A(net209),
    .B(_05899_),
    .Y(_05937_));
 sky130_fd_sc_hd__o21ai_0 _16991_ (.A1(_05611_),
    .A2(_05899_),
    .B1(_05937_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_8 _16992_ (.A(_09901_),
    .B(_05614_),
    .Y(_05938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1231 ();
 sky130_fd_sc_hd__nand2_1 _16995_ (.A(net280),
    .B(_05938_),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_0 _16996_ (.A1(_04988_),
    .A2(_05938_),
    .B1(_05941_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(net279),
    .B(_05938_),
    .Y(_05942_));
 sky130_fd_sc_hd__o21ai_0 _16998_ (.A1(_04992_),
    .A2(_05938_),
    .B1(_05942_),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _16999_ (.A(net277),
    .B(_05938_),
    .Y(_05943_));
 sky130_fd_sc_hd__o21ai_0 _17000_ (.A1(_04995_),
    .A2(_05938_),
    .B1(_05943_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2_1 _17001_ (.A(net276),
    .B(_05938_),
    .Y(_05944_));
 sky130_fd_sc_hd__o21ai_0 _17002_ (.A1(_05003_),
    .A2(_05938_),
    .B1(_05944_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _17003_ (.A(net275),
    .B(_05938_),
    .Y(_05945_));
 sky130_fd_sc_hd__o21ai_0 _17004_ (.A1(_05012_),
    .A2(_05938_),
    .B1(_05945_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _17005_ (.A(net274),
    .B(_05938_),
    .Y(_05946_));
 sky130_fd_sc_hd__o21ai_0 _17006_ (.A1(_05021_),
    .A2(_05938_),
    .B1(_05946_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _17007_ (.A(net273),
    .B(_05938_),
    .Y(_05947_));
 sky130_fd_sc_hd__o21ai_0 _17008_ (.A1(_05032_),
    .A2(_05938_),
    .B1(_05947_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _17009_ (.A(net272),
    .B(_05938_),
    .Y(_05948_));
 sky130_fd_sc_hd__o21ai_0 _17010_ (.A1(_05039_),
    .A2(_05938_),
    .B1(_05948_),
    .Y(_00190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1230 ();
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(net271),
    .B(_05938_),
    .Y(_05950_));
 sky130_fd_sc_hd__o21ai_0 _17013_ (.A1(_05048_),
    .A2(_05938_),
    .B1(_05950_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _17014_ (.A(net270),
    .B(_05938_),
    .Y(_05951_));
 sky130_fd_sc_hd__o21ai_0 _17015_ (.A1(_05055_),
    .A2(_05938_),
    .B1(_05951_),
    .Y(_00192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1229 ();
 sky130_fd_sc_hd__nand2_1 _17017_ (.A(net269),
    .B(_05938_),
    .Y(_05953_));
 sky130_fd_sc_hd__o21ai_0 _17018_ (.A1(_05062_),
    .A2(_05938_),
    .B1(_05953_),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _17019_ (.A(net268),
    .B(_05938_),
    .Y(_05954_));
 sky130_fd_sc_hd__o21ai_0 _17020_ (.A1(_05077_),
    .A2(_05938_),
    .B1(_05954_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _17021_ (.A(net266),
    .B(_05938_),
    .Y(_05955_));
 sky130_fd_sc_hd__o21ai_0 _17022_ (.A1(_05087_),
    .A2(_05938_),
    .B1(_05955_),
    .Y(_00164_));
 sky130_fd_sc_hd__nand2_1 _17023_ (.A(net265),
    .B(_05938_),
    .Y(_05956_));
 sky130_fd_sc_hd__o21ai_0 _17024_ (.A1(_05095_),
    .A2(_05938_),
    .B1(_05956_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _17025_ (.A(net264),
    .B(_05938_),
    .Y(_05957_));
 sky130_fd_sc_hd__o21ai_0 _17026_ (.A1(_05102_),
    .A2(_05938_),
    .B1(_05957_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand2_1 _17027_ (.A(net263),
    .B(_05938_),
    .Y(_05958_));
 sky130_fd_sc_hd__o21ai_0 _17028_ (.A1(_05112_),
    .A2(_05938_),
    .B1(_05958_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _17029_ (.A(net262),
    .B(_05938_),
    .Y(_05959_));
 sky130_fd_sc_hd__o21ai_0 _17030_ (.A1(_05121_),
    .A2(_05938_),
    .B1(_05959_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _17031_ (.A(net261),
    .B(_05938_),
    .Y(_05960_));
 sky130_fd_sc_hd__o21ai_0 _17032_ (.A1(_05128_),
    .A2(_05938_),
    .B1(_05960_),
    .Y(_00169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1228 ();
 sky130_fd_sc_hd__nand2_1 _17034_ (.A(net260),
    .B(_05938_),
    .Y(_05962_));
 sky130_fd_sc_hd__o21ai_0 _17035_ (.A1(_05137_),
    .A2(_05938_),
    .B1(_05962_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_1 _17036_ (.A(net259),
    .B(_05938_),
    .Y(_05963_));
 sky130_fd_sc_hd__o21ai_0 _17037_ (.A1(_05154_),
    .A2(_05938_),
    .B1(_05963_),
    .Y(_00171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1227 ();
 sky130_fd_sc_hd__nand2_1 _17039_ (.A(net258),
    .B(_05938_),
    .Y(_05965_));
 sky130_fd_sc_hd__o21ai_0 _17040_ (.A1(_05167_),
    .A2(_05938_),
    .B1(_05965_),
    .Y(_00173_));
 sky130_fd_sc_hd__nand2_1 _17041_ (.A(net257),
    .B(_05938_),
    .Y(_05966_));
 sky130_fd_sc_hd__o21ai_0 _17042_ (.A1(_05175_),
    .A2(_05938_),
    .B1(_05966_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _17043_ (.A(net255),
    .B(_05938_),
    .Y(_05967_));
 sky130_fd_sc_hd__o21ai_0 _17044_ (.A1(_05184_),
    .A2(_05938_),
    .B1(_05967_),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _17045_ (.A(net254),
    .B(_05938_),
    .Y(_05968_));
 sky130_fd_sc_hd__o21ai_0 _17046_ (.A1(_05196_),
    .A2(_05938_),
    .B1(_05968_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand2_1 _17047_ (.A(net253),
    .B(_05938_),
    .Y(_05969_));
 sky130_fd_sc_hd__o21ai_0 _17048_ (.A1(_05206_),
    .A2(_05938_),
    .B1(_05969_),
    .Y(_00177_));
 sky130_fd_sc_hd__nand2_1 _17049_ (.A(net252),
    .B(_05938_),
    .Y(_05970_));
 sky130_fd_sc_hd__o21ai_0 _17050_ (.A1(_05214_),
    .A2(_05938_),
    .B1(_05970_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _17051_ (.A(net251),
    .B(_05938_),
    .Y(_05971_));
 sky130_fd_sc_hd__o21ai_0 _17052_ (.A1(_05224_),
    .A2(_05938_),
    .B1(_05971_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _17053_ (.A(net250),
    .B(_05938_),
    .Y(_05972_));
 sky130_fd_sc_hd__o21ai_0 _17054_ (.A1(_05236_),
    .A2(_05938_),
    .B1(_05972_),
    .Y(_00180_));
 sky130_fd_sc_hd__nand2_1 _17055_ (.A(net249),
    .B(_05938_),
    .Y(_05973_));
 sky130_fd_sc_hd__o21ai_0 _17056_ (.A1(_05243_),
    .A2(_05938_),
    .B1(_05973_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _17057_ (.A(net248),
    .B(_05938_),
    .Y(_05974_));
 sky130_fd_sc_hd__o21ai_0 _17058_ (.A1(_05251_),
    .A2(_05938_),
    .B1(_05974_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _17059_ (.A(net247),
    .B(_05938_),
    .Y(_05975_));
 sky130_fd_sc_hd__o21ai_0 _17060_ (.A1(_05260_),
    .A2(_05938_),
    .B1(_05975_),
    .Y(_00184_));
 sky130_fd_sc_hd__nand2_1 _17061_ (.A(net246),
    .B(_05938_),
    .Y(_05976_));
 sky130_fd_sc_hd__o21ai_0 _17062_ (.A1(_05310_),
    .A2(_05938_),
    .B1(_05976_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_8 _17063_ (.A(_09946_),
    .B(_05655_),
    .Y(_05977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1225 ();
 sky130_fd_sc_hd__nand2_1 _17066_ (.A(net315),
    .B(_05977_),
    .Y(_05980_));
 sky130_fd_sc_hd__o21ai_0 _17067_ (.A1(_05317_),
    .A2(_05977_),
    .B1(_05980_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _17068_ (.A(net314),
    .B(_05977_),
    .Y(_05981_));
 sky130_fd_sc_hd__o21ai_0 _17069_ (.A1(_05321_),
    .A2(_05977_),
    .B1(_05981_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _17070_ (.A(net313),
    .B(_05977_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21ai_0 _17071_ (.A1(_05324_),
    .A2(_05977_),
    .B1(_05982_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _17072_ (.A(net312),
    .B(_05977_),
    .Y(_05983_));
 sky130_fd_sc_hd__o21ai_0 _17073_ (.A1(_05330_),
    .A2(_05977_),
    .B1(_05983_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _17074_ (.A(net310),
    .B(_05977_),
    .Y(_05984_));
 sky130_fd_sc_hd__o21ai_0 _17075_ (.A1(_05338_),
    .A2(_05977_),
    .B1(_05984_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _17076_ (.A(net309),
    .B(_05977_),
    .Y(_05985_));
 sky130_fd_sc_hd__o21ai_0 _17077_ (.A1(_05347_),
    .A2(_05977_),
    .B1(_05985_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _17078_ (.A(net308),
    .B(_05977_),
    .Y(_05986_));
 sky130_fd_sc_hd__o21ai_0 _17079_ (.A1(_05354_),
    .A2(_05977_),
    .B1(_05986_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _17080_ (.A(net307),
    .B(_05977_),
    .Y(_05987_));
 sky130_fd_sc_hd__o21ai_0 _17081_ (.A1(_05360_),
    .A2(_05977_),
    .B1(_05987_),
    .Y(_00222_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1224 ();
 sky130_fd_sc_hd__nand2_1 _17083_ (.A(net306),
    .B(_05977_),
    .Y(_05989_));
 sky130_fd_sc_hd__o21ai_0 _17084_ (.A1(_05371_),
    .A2(_05977_),
    .B1(_05989_),
    .Y(_00223_));
 sky130_fd_sc_hd__nand2_1 _17085_ (.A(net305),
    .B(_05977_),
    .Y(_05990_));
 sky130_fd_sc_hd__o21ai_0 _17086_ (.A1(_05380_),
    .A2(_05977_),
    .B1(_05990_),
    .Y(_00224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1223 ();
 sky130_fd_sc_hd__nand2_1 _17088_ (.A(net304),
    .B(_05977_),
    .Y(_05992_));
 sky130_fd_sc_hd__o21ai_0 _17089_ (.A1(_05388_),
    .A2(_05977_),
    .B1(_05992_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _17090_ (.A(net303),
    .B(_05977_),
    .Y(_05993_));
 sky130_fd_sc_hd__o21ai_0 _17091_ (.A1(_05402_),
    .A2(_05977_),
    .B1(_05993_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _17092_ (.A(net302),
    .B(_05977_),
    .Y(_05994_));
 sky130_fd_sc_hd__o21ai_0 _17093_ (.A1(_05412_),
    .A2(_05977_),
    .B1(_05994_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _17094_ (.A(net301),
    .B(_05977_),
    .Y(_05995_));
 sky130_fd_sc_hd__o21ai_0 _17095_ (.A1(_05419_),
    .A2(_05977_),
    .B1(_05995_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand2_1 _17096_ (.A(net299),
    .B(_05977_),
    .Y(_05996_));
 sky130_fd_sc_hd__o21ai_0 _17097_ (.A1(_05426_),
    .A2(_05977_),
    .B1(_05996_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _17098_ (.A(net298),
    .B(_05977_),
    .Y(_05997_));
 sky130_fd_sc_hd__o21ai_0 _17099_ (.A1(_05438_),
    .A2(_05977_),
    .B1(_05997_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _17100_ (.A(net297),
    .B(_05977_),
    .Y(_05998_));
 sky130_fd_sc_hd__o21ai_0 _17101_ (.A1(_05447_),
    .A2(_05977_),
    .B1(_05998_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _17102_ (.A(net296),
    .B(_05977_),
    .Y(_05999_));
 sky130_fd_sc_hd__o21ai_0 _17103_ (.A1(_05453_),
    .A2(_05977_),
    .B1(_05999_),
    .Y(_00201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1222 ();
 sky130_fd_sc_hd__nand2_1 _17105_ (.A(net295),
    .B(_05977_),
    .Y(_06001_));
 sky130_fd_sc_hd__o21ai_0 _17106_ (.A1(_05465_),
    .A2(_05977_),
    .B1(_06001_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _17107_ (.A(net294),
    .B(_05977_),
    .Y(_06002_));
 sky130_fd_sc_hd__o21ai_0 _17108_ (.A1(_05480_),
    .A2(_05977_),
    .B1(_06002_),
    .Y(_00203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1221 ();
 sky130_fd_sc_hd__nand2_1 _17110_ (.A(net293),
    .B(_05977_),
    .Y(_06004_));
 sky130_fd_sc_hd__o21ai_0 _17111_ (.A1(_05488_),
    .A2(_05977_),
    .B1(_06004_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _17112_ (.A(net292),
    .B(_05977_),
    .Y(_06005_));
 sky130_fd_sc_hd__o21ai_0 _17113_ (.A1(_05498_),
    .A2(_05977_),
    .B1(_06005_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _17114_ (.A(net291),
    .B(_05977_),
    .Y(_06006_));
 sky130_fd_sc_hd__o21ai_0 _17115_ (.A1(_05509_),
    .A2(_05977_),
    .B1(_06006_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_1 _17116_ (.A(net290),
    .B(_05977_),
    .Y(_06007_));
 sky130_fd_sc_hd__o21ai_0 _17117_ (.A1(_05515_),
    .A2(_05977_),
    .B1(_06007_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _17118_ (.A(net288),
    .B(_05977_),
    .Y(_06008_));
 sky130_fd_sc_hd__o21ai_0 _17119_ (.A1(_05523_),
    .A2(_05977_),
    .B1(_06008_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _17120_ (.A(net287),
    .B(_05977_),
    .Y(_06009_));
 sky130_fd_sc_hd__o21ai_0 _17121_ (.A1(_05535_),
    .A2(_05977_),
    .B1(_06009_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _17122_ (.A(net286),
    .B(_05977_),
    .Y(_06010_));
 sky130_fd_sc_hd__o21ai_0 _17123_ (.A1(_05542_),
    .A2(_05977_),
    .B1(_06010_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _17124_ (.A(net285),
    .B(_05977_),
    .Y(_06011_));
 sky130_fd_sc_hd__o21ai_0 _17125_ (.A1(_05551_),
    .A2(_05977_),
    .B1(_06011_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _17126_ (.A(net284),
    .B(_05977_),
    .Y(_06012_));
 sky130_fd_sc_hd__o21ai_0 _17127_ (.A1(_05559_),
    .A2(_05977_),
    .B1(_06012_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _17128_ (.A(net283),
    .B(_05977_),
    .Y(_06013_));
 sky130_fd_sc_hd__o21ai_0 _17129_ (.A1(_05567_),
    .A2(_05977_),
    .B1(_06013_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(net282),
    .B(_05977_),
    .Y(_06014_));
 sky130_fd_sc_hd__o21ai_0 _17131_ (.A1(_05573_),
    .A2(_05977_),
    .B1(_06014_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _17132_ (.A(net281),
    .B(_05977_),
    .Y(_06015_));
 sky130_fd_sc_hd__o21ai_0 _17133_ (.A1(_05611_),
    .A2(_05977_),
    .B1(_06015_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_8 _17134_ (.A(_09901_),
    .B(_05696_),
    .Y(_06016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1219 ();
 sky130_fd_sc_hd__nand2_1 _17137_ (.A(net351),
    .B(_06016_),
    .Y(_06019_));
 sky130_fd_sc_hd__o21ai_0 _17138_ (.A1(_04988_),
    .A2(_06016_),
    .B1(_06019_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _17139_ (.A(net350),
    .B(_06016_),
    .Y(_06020_));
 sky130_fd_sc_hd__o21ai_0 _17140_ (.A1(_04992_),
    .A2(_06016_),
    .B1(_06020_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _17141_ (.A(net349),
    .B(_06016_),
    .Y(_06021_));
 sky130_fd_sc_hd__o21ai_0 _17142_ (.A1(_04995_),
    .A2(_06016_),
    .B1(_06021_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _17143_ (.A(net348),
    .B(_06016_),
    .Y(_06022_));
 sky130_fd_sc_hd__o21ai_0 _17144_ (.A1(_05003_),
    .A2(_06016_),
    .B1(_06022_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _17145_ (.A(net347),
    .B(_06016_),
    .Y(_06023_));
 sky130_fd_sc_hd__o21ai_0 _17146_ (.A1(_05012_),
    .A2(_06016_),
    .B1(_06023_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _17147_ (.A(net346),
    .B(_06016_),
    .Y(_06024_));
 sky130_fd_sc_hd__o21ai_0 _17148_ (.A1(_05021_),
    .A2(_06016_),
    .B1(_06024_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _17149_ (.A(net344),
    .B(_06016_),
    .Y(_06025_));
 sky130_fd_sc_hd__o21ai_0 _17150_ (.A1(_05032_),
    .A2(_06016_),
    .B1(_06025_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _17151_ (.A(net343),
    .B(_06016_),
    .Y(_06026_));
 sky130_fd_sc_hd__o21ai_0 _17152_ (.A1(_05039_),
    .A2(_06016_),
    .B1(_06026_),
    .Y(_00254_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1218 ();
 sky130_fd_sc_hd__nand2_1 _17154_ (.A(net342),
    .B(_06016_),
    .Y(_06028_));
 sky130_fd_sc_hd__o21ai_0 _17155_ (.A1(_05048_),
    .A2(_06016_),
    .B1(_06028_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _17156_ (.A(net341),
    .B(_06016_),
    .Y(_06029_));
 sky130_fd_sc_hd__o21ai_0 _17157_ (.A1(_05055_),
    .A2(_06016_),
    .B1(_06029_),
    .Y(_00256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1217 ();
 sky130_fd_sc_hd__nand2_1 _17159_ (.A(net340),
    .B(_06016_),
    .Y(_06031_));
 sky130_fd_sc_hd__o21ai_0 _17160_ (.A1(_05062_),
    .A2(_06016_),
    .B1(_06031_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _17161_ (.A(net339),
    .B(_06016_),
    .Y(_06032_));
 sky130_fd_sc_hd__o21ai_0 _17162_ (.A1(_05077_),
    .A2(_06016_),
    .B1(_06032_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _17163_ (.A(net338),
    .B(_06016_),
    .Y(_06033_));
 sky130_fd_sc_hd__o21ai_0 _17164_ (.A1(_05087_),
    .A2(_06016_),
    .B1(_06033_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _17165_ (.A(net337),
    .B(_06016_),
    .Y(_06034_));
 sky130_fd_sc_hd__o21ai_0 _17166_ (.A1(_05095_),
    .A2(_06016_),
    .B1(_06034_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _17167_ (.A(net336),
    .B(_06016_),
    .Y(_06035_));
 sky130_fd_sc_hd__o21ai_0 _17168_ (.A1(_05102_),
    .A2(_06016_),
    .B1(_06035_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _17169_ (.A(net335),
    .B(_06016_),
    .Y(_06036_));
 sky130_fd_sc_hd__o21ai_0 _17170_ (.A1(_05112_),
    .A2(_06016_),
    .B1(_06036_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _17171_ (.A(net332),
    .B(_06016_),
    .Y(_06037_));
 sky130_fd_sc_hd__o21ai_0 _17172_ (.A1(_05121_),
    .A2(_06016_),
    .B1(_06037_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _17173_ (.A(net331),
    .B(_06016_),
    .Y(_06038_));
 sky130_fd_sc_hd__o21ai_0 _17174_ (.A1(_05128_),
    .A2(_06016_),
    .B1(_06038_),
    .Y(_00233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1216 ();
 sky130_fd_sc_hd__nand2_1 _17176_ (.A(net330),
    .B(_06016_),
    .Y(_06040_));
 sky130_fd_sc_hd__o21ai_0 _17177_ (.A1(_05137_),
    .A2(_06016_),
    .B1(_06040_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _17178_ (.A(net329),
    .B(_06016_),
    .Y(_06041_));
 sky130_fd_sc_hd__o21ai_0 _17179_ (.A1(_05154_),
    .A2(_06016_),
    .B1(_06041_),
    .Y(_00235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1215 ();
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(net328),
    .B(_06016_),
    .Y(_06043_));
 sky130_fd_sc_hd__o21ai_0 _17182_ (.A1(_05167_),
    .A2(_06016_),
    .B1(_06043_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _17183_ (.A(net327),
    .B(_06016_),
    .Y(_06044_));
 sky130_fd_sc_hd__o21ai_0 _17184_ (.A1(_05175_),
    .A2(_06016_),
    .B1(_06044_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _17185_ (.A(net326),
    .B(_06016_),
    .Y(_06045_));
 sky130_fd_sc_hd__o21ai_0 _17186_ (.A1(_05184_),
    .A2(_06016_),
    .B1(_06045_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _17187_ (.A(net325),
    .B(_06016_),
    .Y(_06046_));
 sky130_fd_sc_hd__o21ai_0 _17188_ (.A1(_05196_),
    .A2(_06016_),
    .B1(_06046_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _17189_ (.A(net324),
    .B(_06016_),
    .Y(_06047_));
 sky130_fd_sc_hd__o21ai_0 _17190_ (.A1(_05206_),
    .A2(_06016_),
    .B1(_06047_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _17191_ (.A(net323),
    .B(_06016_),
    .Y(_06048_));
 sky130_fd_sc_hd__o21ai_0 _17192_ (.A1(_05214_),
    .A2(_06016_),
    .B1(_06048_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _17193_ (.A(net321),
    .B(_06016_),
    .Y(_06049_));
 sky130_fd_sc_hd__o21ai_0 _17194_ (.A1(_05224_),
    .A2(_06016_),
    .B1(_06049_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _17195_ (.A(net320),
    .B(_06016_),
    .Y(_06050_));
 sky130_fd_sc_hd__o21ai_0 _17196_ (.A1(_05236_),
    .A2(_06016_),
    .B1(_06050_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _17197_ (.A(net319),
    .B(_06016_),
    .Y(_06051_));
 sky130_fd_sc_hd__o21ai_0 _17198_ (.A1(_05243_),
    .A2(_06016_),
    .B1(_06051_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _17199_ (.A(net318),
    .B(_06016_),
    .Y(_06052_));
 sky130_fd_sc_hd__o21ai_0 _17200_ (.A1(_05251_),
    .A2(_06016_),
    .B1(_06052_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _17201_ (.A(net317),
    .B(_06016_),
    .Y(_06053_));
 sky130_fd_sc_hd__o21ai_0 _17202_ (.A1(_05260_),
    .A2(_06016_),
    .B1(_06053_),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _17203_ (.A(net316),
    .B(_06016_),
    .Y(_06054_));
 sky130_fd_sc_hd__o21ai_0 _17204_ (.A1(_05310_),
    .A2(_06016_),
    .B1(_06054_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_8 _17205_ (.A(_09946_),
    .B(_05737_),
    .Y(_06055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1213 ();
 sky130_fd_sc_hd__nand2_1 _17208_ (.A(net386),
    .B(_06055_),
    .Y(_06058_));
 sky130_fd_sc_hd__o21ai_0 _17209_ (.A1(_05317_),
    .A2(_06055_),
    .B1(_06058_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _17210_ (.A(net385),
    .B(_06055_),
    .Y(_06059_));
 sky130_fd_sc_hd__o21ai_0 _17211_ (.A1(_05321_),
    .A2(_06055_),
    .B1(_06059_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _17212_ (.A(net384),
    .B(_06055_),
    .Y(_06060_));
 sky130_fd_sc_hd__o21ai_0 _17213_ (.A1(_05324_),
    .A2(_06055_),
    .B1(_06060_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _17214_ (.A(net383),
    .B(_06055_),
    .Y(_06061_));
 sky130_fd_sc_hd__o21ai_0 _17215_ (.A1(_05330_),
    .A2(_06055_),
    .B1(_06061_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _17216_ (.A(net382),
    .B(_06055_),
    .Y(_06062_));
 sky130_fd_sc_hd__o21ai_0 _17217_ (.A1(_05338_),
    .A2(_06055_),
    .B1(_06062_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _17218_ (.A(net381),
    .B(_06055_),
    .Y(_06063_));
 sky130_fd_sc_hd__o21ai_0 _17219_ (.A1(_05347_),
    .A2(_06055_),
    .B1(_06063_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _17220_ (.A(net380),
    .B(_06055_),
    .Y(_06064_));
 sky130_fd_sc_hd__o21ai_0 _17221_ (.A1(_05354_),
    .A2(_06055_),
    .B1(_06064_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _17222_ (.A(net379),
    .B(_06055_),
    .Y(_06065_));
 sky130_fd_sc_hd__o21ai_0 _17223_ (.A1(_05360_),
    .A2(_06055_),
    .B1(_06065_),
    .Y(_00286_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1212 ();
 sky130_fd_sc_hd__nand2_1 _17225_ (.A(net377),
    .B(_06055_),
    .Y(_06067_));
 sky130_fd_sc_hd__o21ai_0 _17226_ (.A1(_05371_),
    .A2(_06055_),
    .B1(_06067_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _17227_ (.A(net376),
    .B(_06055_),
    .Y(_06068_));
 sky130_fd_sc_hd__o21ai_0 _17228_ (.A1(_05380_),
    .A2(_06055_),
    .B1(_06068_),
    .Y(_00288_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1211 ();
 sky130_fd_sc_hd__nand2_1 _17230_ (.A(net375),
    .B(_06055_),
    .Y(_06070_));
 sky130_fd_sc_hd__o21ai_0 _17231_ (.A1(_05388_),
    .A2(_06055_),
    .B1(_06070_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _17232_ (.A(net374),
    .B(_06055_),
    .Y(_06071_));
 sky130_fd_sc_hd__o21ai_0 _17233_ (.A1(_05402_),
    .A2(_06055_),
    .B1(_06071_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _17234_ (.A(net373),
    .B(_06055_),
    .Y(_06072_));
 sky130_fd_sc_hd__o21ai_0 _17235_ (.A1(_05412_),
    .A2(_06055_),
    .B1(_06072_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _17236_ (.A(net372),
    .B(_06055_),
    .Y(_06073_));
 sky130_fd_sc_hd__o21ai_0 _17237_ (.A1(_05419_),
    .A2(_06055_),
    .B1(_06073_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _17238_ (.A(net371),
    .B(_06055_),
    .Y(_06074_));
 sky130_fd_sc_hd__o21ai_0 _17239_ (.A1(_05426_),
    .A2(_06055_),
    .B1(_06074_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _17240_ (.A(net370),
    .B(_06055_),
    .Y(_06075_));
 sky130_fd_sc_hd__o21ai_0 _17241_ (.A1(_05438_),
    .A2(_06055_),
    .B1(_06075_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _17242_ (.A(net369),
    .B(_06055_),
    .Y(_06076_));
 sky130_fd_sc_hd__o21ai_0 _17243_ (.A1(_05447_),
    .A2(_06055_),
    .B1(_06076_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _17244_ (.A(net368),
    .B(_06055_),
    .Y(_06077_));
 sky130_fd_sc_hd__o21ai_0 _17245_ (.A1(_05453_),
    .A2(_06055_),
    .B1(_06077_),
    .Y(_00265_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1210 ();
 sky130_fd_sc_hd__nand2_1 _17247_ (.A(net366),
    .B(_06055_),
    .Y(_06079_));
 sky130_fd_sc_hd__o21ai_0 _17248_ (.A1(_05465_),
    .A2(_06055_),
    .B1(_06079_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_1 _17249_ (.A(net365),
    .B(_06055_),
    .Y(_06080_));
 sky130_fd_sc_hd__o21ai_0 _17250_ (.A1(_05480_),
    .A2(_06055_),
    .B1(_06080_),
    .Y(_00267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1209 ();
 sky130_fd_sc_hd__nand2_1 _17252_ (.A(net364),
    .B(_06055_),
    .Y(_06082_));
 sky130_fd_sc_hd__o21ai_0 _17253_ (.A1(_05488_),
    .A2(_06055_),
    .B1(_06082_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _17254_ (.A(net363),
    .B(_06055_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_0 _17255_ (.A1(_05498_),
    .A2(_06055_),
    .B1(_06083_),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _17256_ (.A(net362),
    .B(_06055_),
    .Y(_06084_));
 sky130_fd_sc_hd__o21ai_0 _17257_ (.A1(_05509_),
    .A2(_06055_),
    .B1(_06084_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _17258_ (.A(net361),
    .B(_06055_),
    .Y(_06085_));
 sky130_fd_sc_hd__o21ai_0 _17259_ (.A1(_05515_),
    .A2(_06055_),
    .B1(_06085_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _17260_ (.A(net360),
    .B(_06055_),
    .Y(_06086_));
 sky130_fd_sc_hd__o21ai_0 _17261_ (.A1(_05523_),
    .A2(_06055_),
    .B1(_06086_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _17262_ (.A(net359),
    .B(_06055_),
    .Y(_06087_));
 sky130_fd_sc_hd__o21ai_0 _17263_ (.A1(_05535_),
    .A2(_06055_),
    .B1(_06087_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _17264_ (.A(net358),
    .B(_06055_),
    .Y(_06088_));
 sky130_fd_sc_hd__o21ai_0 _17265_ (.A1(_05542_),
    .A2(_06055_),
    .B1(_06088_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _17266_ (.A(net357),
    .B(_06055_),
    .Y(_06089_));
 sky130_fd_sc_hd__o21ai_0 _17267_ (.A1(_05551_),
    .A2(_06055_),
    .B1(_06089_),
    .Y(_00276_));
 sky130_fd_sc_hd__nand2_1 _17268_ (.A(net355),
    .B(_06055_),
    .Y(_06090_));
 sky130_fd_sc_hd__o21ai_0 _17269_ (.A1(_05559_),
    .A2(_06055_),
    .B1(_06090_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _17270_ (.A(net354),
    .B(_06055_),
    .Y(_06091_));
 sky130_fd_sc_hd__o21ai_0 _17271_ (.A1(_05567_),
    .A2(_06055_),
    .B1(_06091_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _17272_ (.A(net353),
    .B(_06055_),
    .Y(_06092_));
 sky130_fd_sc_hd__o21ai_0 _17273_ (.A1(_05573_),
    .A2(_06055_),
    .B1(_06092_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _17274_ (.A(net352),
    .B(_06055_),
    .Y(_06093_));
 sky130_fd_sc_hd__o21ai_0 _17275_ (.A1(_05611_),
    .A2(_06055_),
    .B1(_06093_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_8 _17276_ (.A(_09901_),
    .B(_05778_),
    .Y(_06094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1207 ();
 sky130_fd_sc_hd__nand2_1 _17279_ (.A(net421),
    .B(_06094_),
    .Y(_06097_));
 sky130_fd_sc_hd__o21ai_0 _17280_ (.A1(_04988_),
    .A2(_06094_),
    .B1(_06097_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _17281_ (.A(net420),
    .B(_06094_),
    .Y(_06098_));
 sky130_fd_sc_hd__o21ai_0 _17282_ (.A1(_04992_),
    .A2(_06094_),
    .B1(_06098_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _17283_ (.A(net419),
    .B(_06094_),
    .Y(_06099_));
 sky130_fd_sc_hd__o21ai_0 _17284_ (.A1(_04995_),
    .A2(_06094_),
    .B1(_06099_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _17285_ (.A(net418),
    .B(_06094_),
    .Y(_06100_));
 sky130_fd_sc_hd__o21ai_0 _17286_ (.A1(_05003_),
    .A2(_06094_),
    .B1(_06100_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _17287_ (.A(net417),
    .B(_06094_),
    .Y(_06101_));
 sky130_fd_sc_hd__o21ai_0 _17288_ (.A1(_05012_),
    .A2(_06094_),
    .B1(_06101_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _17289_ (.A(net416),
    .B(_06094_),
    .Y(_06102_));
 sky130_fd_sc_hd__o21ai_0 _17290_ (.A1(_05021_),
    .A2(_06094_),
    .B1(_06102_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _17291_ (.A(net415),
    .B(_06094_),
    .Y(_06103_));
 sky130_fd_sc_hd__o21ai_0 _17292_ (.A1(_05032_),
    .A2(_06094_),
    .B1(_06103_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _17293_ (.A(net414),
    .B(_06094_),
    .Y(_06104_));
 sky130_fd_sc_hd__o21ai_0 _17294_ (.A1(_05039_),
    .A2(_06094_),
    .B1(_06104_),
    .Y(_00318_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1206 ();
 sky130_fd_sc_hd__nand2_1 _17296_ (.A(net413),
    .B(_06094_),
    .Y(_06106_));
 sky130_fd_sc_hd__o21ai_0 _17297_ (.A1(_05048_),
    .A2(_06094_),
    .B1(_06106_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _17298_ (.A(net412),
    .B(_06094_),
    .Y(_06107_));
 sky130_fd_sc_hd__o21ai_0 _17299_ (.A1(_05055_),
    .A2(_06094_),
    .B1(_06107_),
    .Y(_00320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1205 ();
 sky130_fd_sc_hd__nand2_1 _17301_ (.A(net410),
    .B(_06094_),
    .Y(_06109_));
 sky130_fd_sc_hd__o21ai_0 _17302_ (.A1(_05062_),
    .A2(_06094_),
    .B1(_06109_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _17303_ (.A(net409),
    .B(_06094_),
    .Y(_06110_));
 sky130_fd_sc_hd__o21ai_0 _17304_ (.A1(_05077_),
    .A2(_06094_),
    .B1(_06110_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _17305_ (.A(net408),
    .B(_06094_),
    .Y(_06111_));
 sky130_fd_sc_hd__o21ai_0 _17306_ (.A1(_05087_),
    .A2(_06094_),
    .B1(_06111_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _17307_ (.A(net407),
    .B(_06094_),
    .Y(_06112_));
 sky130_fd_sc_hd__o21ai_0 _17308_ (.A1(_05095_),
    .A2(_06094_),
    .B1(_06112_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _17309_ (.A(net406),
    .B(_06094_),
    .Y(_06113_));
 sky130_fd_sc_hd__o21ai_0 _17310_ (.A1(_05102_),
    .A2(_06094_),
    .B1(_06113_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(net405),
    .B(_06094_),
    .Y(_06114_));
 sky130_fd_sc_hd__o21ai_0 _17312_ (.A1(_05112_),
    .A2(_06094_),
    .B1(_06114_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _17313_ (.A(net404),
    .B(_06094_),
    .Y(_06115_));
 sky130_fd_sc_hd__o21ai_0 _17314_ (.A1(_05121_),
    .A2(_06094_),
    .B1(_06115_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _17315_ (.A(net403),
    .B(_06094_),
    .Y(_06116_));
 sky130_fd_sc_hd__o21ai_0 _17316_ (.A1(_05128_),
    .A2(_06094_),
    .B1(_06116_),
    .Y(_00297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1204 ();
 sky130_fd_sc_hd__nand2_1 _17318_ (.A(net402),
    .B(_06094_),
    .Y(_06118_));
 sky130_fd_sc_hd__o21ai_0 _17319_ (.A1(_05137_),
    .A2(_06094_),
    .B1(_06118_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _17320_ (.A(net401),
    .B(_06094_),
    .Y(_06119_));
 sky130_fd_sc_hd__o21ai_0 _17321_ (.A1(_05154_),
    .A2(_06094_),
    .B1(_06119_),
    .Y(_00299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1203 ();
 sky130_fd_sc_hd__nand2_1 _17323_ (.A(net399),
    .B(_06094_),
    .Y(_06121_));
 sky130_fd_sc_hd__o21ai_0 _17324_ (.A1(_05167_),
    .A2(_06094_),
    .B1(_06121_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _17325_ (.A(net398),
    .B(_06094_),
    .Y(_06122_));
 sky130_fd_sc_hd__o21ai_0 _17326_ (.A1(_05175_),
    .A2(_06094_),
    .B1(_06122_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _17327_ (.A(net397),
    .B(_06094_),
    .Y(_06123_));
 sky130_fd_sc_hd__o21ai_0 _17328_ (.A1(_05184_),
    .A2(_06094_),
    .B1(_06123_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _17329_ (.A(net396),
    .B(_06094_),
    .Y(_06124_));
 sky130_fd_sc_hd__o21ai_0 _17330_ (.A1(_05196_),
    .A2(_06094_),
    .B1(_06124_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _17331_ (.A(net395),
    .B(_06094_),
    .Y(_06125_));
 sky130_fd_sc_hd__o21ai_0 _17332_ (.A1(_05206_),
    .A2(_06094_),
    .B1(_06125_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _17333_ (.A(net394),
    .B(_06094_),
    .Y(_06126_));
 sky130_fd_sc_hd__o21ai_0 _17334_ (.A1(_05214_),
    .A2(_06094_),
    .B1(_06126_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _17335_ (.A(net393),
    .B(_06094_),
    .Y(_06127_));
 sky130_fd_sc_hd__o21ai_0 _17336_ (.A1(_05224_),
    .A2(_06094_),
    .B1(_06127_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _17337_ (.A(net392),
    .B(_06094_),
    .Y(_06128_));
 sky130_fd_sc_hd__o21ai_0 _17338_ (.A1(_05236_),
    .A2(_06094_),
    .B1(_06128_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _17339_ (.A(net391),
    .B(_06094_),
    .Y(_06129_));
 sky130_fd_sc_hd__o21ai_0 _17340_ (.A1(_05243_),
    .A2(_06094_),
    .B1(_06129_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand2_1 _17341_ (.A(net390),
    .B(_06094_),
    .Y(_06130_));
 sky130_fd_sc_hd__o21ai_0 _17342_ (.A1(_05251_),
    .A2(_06094_),
    .B1(_06130_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _17343_ (.A(net388),
    .B(_06094_),
    .Y(_06131_));
 sky130_fd_sc_hd__o21ai_0 _17344_ (.A1(_05260_),
    .A2(_06094_),
    .B1(_06131_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _17345_ (.A(net387),
    .B(_06094_),
    .Y(_06132_));
 sky130_fd_sc_hd__o21ai_0 _17346_ (.A1(_05310_),
    .A2(_06094_),
    .B1(_06132_),
    .Y(_00313_));
 sky130_fd_sc_hd__nor2b_4 _17347_ (.A(net762),
    .B_N(_13709_),
    .Y(_06133_));
 sky130_fd_sc_hd__nand2_8 _17348_ (.A(_09946_),
    .B(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1201 ();
 sky130_fd_sc_hd__nand2_1 _17351_ (.A(net707),
    .B(_06134_),
    .Y(_06137_));
 sky130_fd_sc_hd__o21ai_0 _17352_ (.A1(_05317_),
    .A2(_06134_),
    .B1(_06137_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _17353_ (.A(net706),
    .B(_06134_),
    .Y(_06138_));
 sky130_fd_sc_hd__o21ai_0 _17354_ (.A1(_05321_),
    .A2(_06134_),
    .B1(_06138_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _17355_ (.A(net704),
    .B(_06134_),
    .Y(_06139_));
 sky130_fd_sc_hd__o21ai_0 _17356_ (.A1(_05324_),
    .A2(_06134_),
    .B1(_06139_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _17357_ (.A(net703),
    .B(_06134_),
    .Y(_06140_));
 sky130_fd_sc_hd__o21ai_0 _17358_ (.A1(_05330_),
    .A2(_06134_),
    .B1(_06140_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _17359_ (.A(net702),
    .B(_06134_),
    .Y(_06141_));
 sky130_fd_sc_hd__o21ai_0 _17360_ (.A1(_05338_),
    .A2(_06134_),
    .B1(_06141_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _17361_ (.A(net452),
    .B(_06134_),
    .Y(_06142_));
 sky130_fd_sc_hd__o21ai_0 _17362_ (.A1(_05347_),
    .A2(_06134_),
    .B1(_06142_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _17363_ (.A(net451),
    .B(_06134_),
    .Y(_06143_));
 sky130_fd_sc_hd__o21ai_0 _17364_ (.A1(_05354_),
    .A2(_06134_),
    .B1(_06143_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _17365_ (.A(net450),
    .B(_06134_),
    .Y(_06144_));
 sky130_fd_sc_hd__o21ai_0 _17366_ (.A1(_05360_),
    .A2(_06134_),
    .B1(_06144_),
    .Y(_00350_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1200 ();
 sky130_fd_sc_hd__nand2_1 _17368_ (.A(net449),
    .B(_06134_),
    .Y(_06146_));
 sky130_fd_sc_hd__o21ai_0 _17369_ (.A1(_05371_),
    .A2(_06134_),
    .B1(_06146_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _17370_ (.A(net448),
    .B(_06134_),
    .Y(_06147_));
 sky130_fd_sc_hd__o21ai_0 _17371_ (.A1(_05380_),
    .A2(_06134_),
    .B1(_06147_),
    .Y(_00352_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1199 ();
 sky130_fd_sc_hd__nand2_1 _17373_ (.A(net447),
    .B(_06134_),
    .Y(_06149_));
 sky130_fd_sc_hd__o21ai_0 _17374_ (.A1(_05388_),
    .A2(_06134_),
    .B1(_06149_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _17375_ (.A(net446),
    .B(_06134_),
    .Y(_06150_));
 sky130_fd_sc_hd__o21ai_0 _17376_ (.A1(_05402_),
    .A2(_06134_),
    .B1(_06150_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _17377_ (.A(net443),
    .B(_06134_),
    .Y(_06151_));
 sky130_fd_sc_hd__o21ai_0 _17378_ (.A1(_05412_),
    .A2(_06134_),
    .B1(_06151_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _17379_ (.A(net442),
    .B(_06134_),
    .Y(_06152_));
 sky130_fd_sc_hd__o21ai_0 _17380_ (.A1(_05419_),
    .A2(_06134_),
    .B1(_06152_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _17381_ (.A(net441),
    .B(_06134_),
    .Y(_06153_));
 sky130_fd_sc_hd__o21ai_0 _17382_ (.A1(_05426_),
    .A2(_06134_),
    .B1(_06153_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _17383_ (.A(net440),
    .B(_06134_),
    .Y(_06154_));
 sky130_fd_sc_hd__o21ai_0 _17384_ (.A1(_05438_),
    .A2(_06134_),
    .B1(_06154_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _17385_ (.A(net439),
    .B(_06134_),
    .Y(_06155_));
 sky130_fd_sc_hd__o21ai_0 _17386_ (.A1(_05447_),
    .A2(_06134_),
    .B1(_06155_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _17387_ (.A(net438),
    .B(_06134_),
    .Y(_06156_));
 sky130_fd_sc_hd__o21ai_0 _17388_ (.A1(_05453_),
    .A2(_06134_),
    .B1(_06156_),
    .Y(_00329_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1198 ();
 sky130_fd_sc_hd__nand2_1 _17390_ (.A(net437),
    .B(_06134_),
    .Y(_06158_));
 sky130_fd_sc_hd__o21ai_0 _17391_ (.A1(_05465_),
    .A2(_06134_),
    .B1(_06158_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _17392_ (.A(net436),
    .B(_06134_),
    .Y(_06159_));
 sky130_fd_sc_hd__o21ai_0 _17393_ (.A1(_05480_),
    .A2(_06134_),
    .B1(_06159_),
    .Y(_00331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1197 ();
 sky130_fd_sc_hd__nand2_1 _17395_ (.A(net435),
    .B(_06134_),
    .Y(_06161_));
 sky130_fd_sc_hd__o21ai_0 _17396_ (.A1(_05488_),
    .A2(_06134_),
    .B1(_06161_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _17397_ (.A(net434),
    .B(_06134_),
    .Y(_06162_));
 sky130_fd_sc_hd__o21ai_0 _17398_ (.A1(_05498_),
    .A2(_06134_),
    .B1(_06162_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _17399_ (.A(net432),
    .B(_06134_),
    .Y(_06163_));
 sky130_fd_sc_hd__o21ai_0 _17400_ (.A1(_05509_),
    .A2(_06134_),
    .B1(_06163_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _17401_ (.A(net431),
    .B(_06134_),
    .Y(_06164_));
 sky130_fd_sc_hd__o21ai_0 _17402_ (.A1(_05515_),
    .A2(_06134_),
    .B1(_06164_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _17403_ (.A(net430),
    .B(_06134_),
    .Y(_06165_));
 sky130_fd_sc_hd__o21ai_0 _17404_ (.A1(_05523_),
    .A2(_06134_),
    .B1(_06165_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _17405_ (.A(net429),
    .B(_06134_),
    .Y(_06166_));
 sky130_fd_sc_hd__o21ai_0 _17406_ (.A1(_05535_),
    .A2(_06134_),
    .B1(_06166_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _17407_ (.A(net428),
    .B(_06134_),
    .Y(_06167_));
 sky130_fd_sc_hd__o21ai_0 _17408_ (.A1(_05542_),
    .A2(_06134_),
    .B1(_06167_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _17409_ (.A(net427),
    .B(_06134_),
    .Y(_06168_));
 sky130_fd_sc_hd__o21ai_0 _17410_ (.A1(_05551_),
    .A2(_06134_),
    .B1(_06168_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_1 _17411_ (.A(net426),
    .B(_06134_),
    .Y(_06169_));
 sky130_fd_sc_hd__o21ai_0 _17412_ (.A1(_05559_),
    .A2(_06134_),
    .B1(_06169_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _17413_ (.A(net425),
    .B(_06134_),
    .Y(_06170_));
 sky130_fd_sc_hd__o21ai_0 _17414_ (.A1(_05567_),
    .A2(_06134_),
    .B1(_06170_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_1 _17415_ (.A(net424),
    .B(_06134_),
    .Y(_06171_));
 sky130_fd_sc_hd__o21ai_0 _17416_ (.A1(_05573_),
    .A2(_06134_),
    .B1(_06171_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _17417_ (.A(net423),
    .B(_06134_),
    .Y(_06172_));
 sky130_fd_sc_hd__o21ai_0 _17418_ (.A1(_05611_),
    .A2(_06134_),
    .B1(_06172_),
    .Y(_00345_));
 sky130_fd_sc_hd__or2_2 _17419_ (.A(\hash.reset ),
    .B(\hash.CA2.f_dash[0] ),
    .X(_12824_));
 sky130_fd_sc_hd__inv_1 _17420_ (.A(_12824_),
    .Y(_00875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1195 ();
 sky130_fd_sc_hd__nor2_2 _17423_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[0] ),
    .Y(_00843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1194 ();
 sky130_fd_sc_hd__nor2_2 _17425_ (.A(net520),
    .B(_12281_),
    .Y(_06176_));
 sky130_fd_sc_hd__clkinvlp_4 _17426_ (.A(_06176_),
    .Y(\hash.CA1.S0.X[2] ));
 sky130_fd_sc_hd__xnor2_1 _17427_ (.A(_13712_),
    .B(_06176_),
    .Y(_00680_));
 sky130_fd_sc_hd__and2b_1 _17428_ (.A_N(_12280_),
    .B(_13423_),
    .X(_06177_));
 sky130_fd_sc_hd__nor2b_1 _17429_ (.A(_13423_),
    .B_N(_12280_),
    .Y(_06178_));
 sky130_fd_sc_hd__or3_4 _17430_ (.A(net520),
    .B(_06177_),
    .C(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__inv_4 _17431_ (.A(_06179_),
    .Y(\hash.CA1.S0.X[3] ));
 sky130_fd_sc_hd__clkinv_2 _17432_ (.A(_00658_),
    .Y(\hash.CA1.S0.X[0] ));
 sky130_fd_sc_hd__nor3_1 _17433_ (.A(_13409_),
    .B(_12281_),
    .C(\hash.CA1.S0.X[0] ),
    .Y(_06180_));
 sky130_fd_sc_hd__xnor2_1 _17434_ (.A(\hash.CA1.S0.X[3] ),
    .B(_06180_),
    .Y(_00683_));
 sky130_fd_sc_hd__a21o_1 _17435_ (.A1(_13408_),
    .A2(_13416_),
    .B1(_13415_),
    .X(_06181_));
 sky130_fd_sc_hd__a21oi_2 _17436_ (.A1(_13423_),
    .A2(_06181_),
    .B1(_13422_),
    .Y(_06182_));
 sky130_fd_sc_hd__xor2_4 _17437_ (.A(_13430_),
    .B(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__nor2_8 _17438_ (.A(net520),
    .B(_06183_),
    .Y(\hash.CA1.S0.X[4] ));
 sky130_fd_sc_hd__nand2_1 _17439_ (.A(_13712_),
    .B(_06176_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _17440_ (.A(\hash.CA1.S0.X[3] ),
    .B(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__xnor2_1 _17441_ (.A(\hash.CA1.S0.X[4] ),
    .B(_06185_),
    .Y(_00684_));
 sky130_fd_sc_hd__o21a_1 _17442_ (.A1(_13422_),
    .A2(_06177_),
    .B1(_13430_),
    .X(_06186_));
 sky130_fd_sc_hd__o21a_1 _17443_ (.A1(_13429_),
    .A2(_06186_),
    .B1(_13437_),
    .X(_06187_));
 sky130_fd_sc_hd__nor3_1 _17444_ (.A(_13437_),
    .B(_13429_),
    .C(_06186_),
    .Y(_06188_));
 sky130_fd_sc_hd__nor2_2 _17445_ (.A(_06187_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nor2_8 _17446_ (.A(net520),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__clkinvlp_4 _17447_ (.A(_06190_),
    .Y(\hash.CA1.S0.X[5] ));
 sky130_fd_sc_hd__nor2_1 _17448_ (.A(_06179_),
    .B(_06180_),
    .Y(_06191_));
 sky130_fd_sc_hd__nand2_1 _17449_ (.A(_06191_),
    .B(\hash.CA1.S0.X[4] ),
    .Y(_06192_));
 sky130_fd_sc_hd__xnor2_1 _17450_ (.A(_06190_),
    .B(_06192_),
    .Y(_00685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1193 ();
 sky130_fd_sc_hd__o21a_2 _17452_ (.A1(_13430_),
    .A2(_13429_),
    .B1(_13437_),
    .X(_06194_));
 sky130_fd_sc_hd__a211o_1 _17453_ (.A1(_13423_),
    .A2(_06181_),
    .B1(_13429_),
    .C1(_13422_),
    .X(_06195_));
 sky130_fd_sc_hd__a21oi_2 _17454_ (.A1(_06194_),
    .A2(_06195_),
    .B1(_13436_),
    .Y(_06196_));
 sky130_fd_sc_hd__xnor2_4 _17455_ (.A(_13444_),
    .B(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__nor2_4 _17456_ (.A(net520),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__clkinv_4 _17457_ (.A(_06198_),
    .Y(\hash.CA1.S0.X[6] ));
 sky130_fd_sc_hd__nor3_2 _17458_ (.A(net520),
    .B(_06183_),
    .C(_06185_),
    .Y(_06199_));
 sky130_fd_sc_hd__nor2_1 _17459_ (.A(\hash.CA1.S0.X[5] ),
    .B(_06199_),
    .Y(_06200_));
 sky130_fd_sc_hd__xnor2_1 _17460_ (.A(_06198_),
    .B(_06200_),
    .Y(_00686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1192 ();
 sky130_fd_sc_hd__o311a_1 _17462_ (.A1(_13422_),
    .A2(_13429_),
    .A3(_06177_),
    .B1(_06194_),
    .C1(_13444_),
    .X(_06202_));
 sky130_fd_sc_hd__a21o_1 _17463_ (.A1(_13444_),
    .A2(_13436_),
    .B1(_13443_),
    .X(_06203_));
 sky130_fd_sc_hd__nor3_1 _17464_ (.A(_13451_),
    .B(_06202_),
    .C(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__o311ai_4 _17465_ (.A1(_13422_),
    .A2(_13429_),
    .A3(_06177_),
    .B1(_06194_),
    .C1(_13444_),
    .Y(_06205_));
 sky130_fd_sc_hd__a21oi_1 _17466_ (.A1(_13444_),
    .A2(_13436_),
    .B1(_13443_),
    .Y(_06206_));
 sky130_fd_sc_hd__a21boi_1 _17467_ (.A1(_06205_),
    .A2(_06206_),
    .B1_N(_13451_),
    .Y(_06207_));
 sky130_fd_sc_hd__nor3_4 _17468_ (.A(net520),
    .B(_06204_),
    .C(_06207_),
    .Y(\hash.CA1.S0.X[7] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1191 ();
 sky130_fd_sc_hd__a2111o_2 _17470_ (.A1(_06191_),
    .A2(\hash.CA1.S0.X[4] ),
    .B1(\hash.CA1.S0.X[5] ),
    .C1(_06197_),
    .D1(net520),
    .X(_06209_));
 sky130_fd_sc_hd__xor2_1 _17471_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06209_),
    .X(_00687_));
 sky130_fd_sc_hd__clkinv_16 _17472_ (.A(net522),
    .Y(_06210_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1190 ();
 sky130_fd_sc_hd__o21a_1 _17474_ (.A1(_13444_),
    .A2(_13443_),
    .B1(_13451_),
    .X(_06212_));
 sky130_fd_sc_hd__nor2_1 _17475_ (.A(_13450_),
    .B(_06212_),
    .Y(_06213_));
 sky130_fd_sc_hd__inv_1 _17476_ (.A(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__a2111o_2 _17477_ (.A1(_06194_),
    .A2(_06195_),
    .B1(_13436_),
    .C1(_13443_),
    .D1(_13450_),
    .X(_06215_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1189 ();
 sky130_fd_sc_hd__a21o_1 _17479_ (.A1(_06214_),
    .A2(_06215_),
    .B1(_13458_),
    .X(_06217_));
 sky130_fd_sc_hd__nand3_1 _17480_ (.A(_13458_),
    .B(_06214_),
    .C(_06215_),
    .Y(_06218_));
 sky130_fd_sc_hd__nand3_4 _17481_ (.A(net519),
    .B(_06217_),
    .C(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__clkinv_4 _17482_ (.A(_06219_),
    .Y(\hash.CA1.S0.X[8] ));
 sky130_fd_sc_hd__o41ai_4 _17483_ (.A1(net520),
    .A2(\hash.CA1.S0.X[5] ),
    .A3(_06197_),
    .A4(_06199_),
    .B1(\hash.CA1.S0.X[7] ),
    .Y(_06220_));
 sky130_fd_sc_hd__xnor2_1 _17484_ (.A(\hash.CA1.S0.X[8] ),
    .B(_06220_),
    .Y(_00688_));
 sky130_fd_sc_hd__a21o_1 _17485_ (.A1(_13458_),
    .A2(_13450_),
    .B1(_13457_),
    .X(_06221_));
 sky130_fd_sc_hd__nand2_1 _17486_ (.A(_13451_),
    .B(_13458_),
    .Y(_06222_));
 sky130_fd_sc_hd__a21oi_1 _17487_ (.A1(_06205_),
    .A2(_06206_),
    .B1(_06222_),
    .Y(_06223_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1188 ();
 sky130_fd_sc_hd__o21a_1 _17489_ (.A1(_06221_),
    .A2(_06223_),
    .B1(_13465_),
    .X(_06225_));
 sky130_fd_sc_hd__nor3_1 _17490_ (.A(_13465_),
    .B(_06221_),
    .C(_06223_),
    .Y(_06226_));
 sky130_fd_sc_hd__o21a_4 _17491_ (.A1(_06225_),
    .A2(_06226_),
    .B1(net519),
    .X(_06227_));
 sky130_fd_sc_hd__inv_2 _17492_ (.A(_06227_),
    .Y(\hash.CA1.S0.X[9] ));
 sky130_fd_sc_hd__nand3_1 _17493_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06209_),
    .C(\hash.CA1.S0.X[8] ),
    .Y(_06228_));
 sky130_fd_sc_hd__xnor2_1 _17494_ (.A(_06227_),
    .B(_06228_),
    .Y(_00689_));
 sky130_fd_sc_hd__inv_1 _17495_ (.A(_13472_),
    .Y(_06229_));
 sky130_fd_sc_hd__or3_1 _17496_ (.A(_06229_),
    .B(_13457_),
    .C(_13464_),
    .X(_06230_));
 sky130_fd_sc_hd__a31oi_1 _17497_ (.A1(_13458_),
    .A2(_06214_),
    .A3(_06215_),
    .B1(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__nor2b_1 _17498_ (.A(_13472_),
    .B_N(_13465_),
    .Y(_06232_));
 sky130_fd_sc_hd__nor3_1 _17499_ (.A(_13465_),
    .B(_06229_),
    .C(_13464_),
    .Y(_06233_));
 sky130_fd_sc_hd__a221oi_1 _17500_ (.A1(_06229_),
    .A2(_13464_),
    .B1(_06232_),
    .B2(_13457_),
    .C1(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__nand4_1 _17501_ (.A(_13458_),
    .B(_06214_),
    .C(_06215_),
    .D(_06232_),
    .Y(_06235_));
 sky130_fd_sc_hd__and4b_4 _17502_ (.A_N(_06231_),
    .B(_06234_),
    .C(_06235_),
    .D(net519),
    .X(_06236_));
 sky130_fd_sc_hd__clkinv_4 _17503_ (.A(_06236_),
    .Y(\hash.CA1.S0.X[10] ));
 sky130_fd_sc_hd__o21ai_0 _17504_ (.A1(_06219_),
    .A2(_06220_),
    .B1(_06227_),
    .Y(_06237_));
 sky130_fd_sc_hd__xnor2_1 _17505_ (.A(\hash.CA1.S0.X[10] ),
    .B(_06237_),
    .Y(_00659_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1187 ();
 sky130_fd_sc_hd__nand4_2 _17507_ (.A(_13451_),
    .B(_13458_),
    .C(_13465_),
    .D(_13472_),
    .Y(_06239_));
 sky130_fd_sc_hd__a21oi_1 _17508_ (.A1(_06205_),
    .A2(_06206_),
    .B1(_06239_),
    .Y(_06240_));
 sky130_fd_sc_hd__a21oi_1 _17509_ (.A1(_13465_),
    .A2(_06221_),
    .B1(_13464_),
    .Y(_06241_));
 sky130_fd_sc_hd__nor2_1 _17510_ (.A(_06229_),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__nor3_4 _17511_ (.A(_13471_),
    .B(_06240_),
    .C(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__xor2_4 _17512_ (.A(_13479_),
    .B(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__nor2_8 _17513_ (.A(net520),
    .B(_06244_),
    .Y(\hash.CA1.S0.X[11] ));
 sky130_fd_sc_hd__a311o_1 _17514_ (.A1(\hash.CA1.S0.X[7] ),
    .A2(_06209_),
    .A3(\hash.CA1.S0.X[8] ),
    .B1(\hash.CA1.S0.X[9] ),
    .C1(\hash.CA1.S0.X[10] ),
    .X(_06245_));
 sky130_fd_sc_hd__xor2_1 _17515_ (.A(\hash.CA1.S0.X[11] ),
    .B(_06245_),
    .X(_00660_));
 sky130_fd_sc_hd__and4_1 _17516_ (.A(_13458_),
    .B(_13465_),
    .C(_13472_),
    .D(_13479_),
    .X(_06246_));
 sky130_fd_sc_hd__a21o_1 _17517_ (.A1(_13465_),
    .A2(_13457_),
    .B1(_13464_),
    .X(_06247_));
 sky130_fd_sc_hd__a21oi_1 _17518_ (.A1(_13472_),
    .A2(_06247_),
    .B1(_13471_),
    .Y(_06248_));
 sky130_fd_sc_hd__nor2b_1 _17519_ (.A(_06248_),
    .B_N(_13479_),
    .Y(_06249_));
 sky130_fd_sc_hd__a311o_2 _17520_ (.A1(_06214_),
    .A2(_06215_),
    .A3(_06246_),
    .B1(_06249_),
    .C1(_13478_),
    .X(_06250_));
 sky130_fd_sc_hd__xnor2_4 _17521_ (.A(_13486_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__nor2_4 _17522_ (.A(net524),
    .B(_06251_),
    .Y(\hash.CA1.S0.X[12] ));
 sky130_fd_sc_hd__o211ai_1 _17523_ (.A1(_06219_),
    .A2(_06220_),
    .B1(_06227_),
    .C1(_06236_),
    .Y(_06252_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(\hash.CA1.S0.X[11] ),
    .B(_06252_),
    .Y(_06253_));
 sky130_fd_sc_hd__xnor2_1 _17525_ (.A(\hash.CA1.S0.X[12] ),
    .B(_06253_),
    .Y(_00661_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1186 ();
 sky130_fd_sc_hd__nand2_1 _17527_ (.A(_13479_),
    .B(_13486_),
    .Y(_06255_));
 sky130_fd_sc_hd__a21oi_1 _17528_ (.A1(_13486_),
    .A2(_13478_),
    .B1(_13485_),
    .Y(_06256_));
 sky130_fd_sc_hd__o21ai_2 _17529_ (.A1(_06243_),
    .A2(_06255_),
    .B1(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__xor2_4 _17530_ (.A(_13493_),
    .B(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__nor2_2 _17531_ (.A(net524),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__inv_1 _17532_ (.A(_06259_),
    .Y(\hash.CA1.S0.X[13] ));
 sky130_fd_sc_hd__nand3_4 _17533_ (.A(\hash.CA1.S0.X[11] ),
    .B(_06245_),
    .C(\hash.CA1.S0.X[12] ),
    .Y(_06260_));
 sky130_fd_sc_hd__xnor2_1 _17534_ (.A(_06259_),
    .B(_06260_),
    .Y(_00662_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1184 ();
 sky130_fd_sc_hd__nor2_1 _17537_ (.A(_13444_),
    .B(_13443_),
    .Y(_06263_));
 sky130_fd_sc_hd__a211oi_2 _17538_ (.A1(_06194_),
    .A2(_06195_),
    .B1(_13436_),
    .C1(_13443_),
    .Y(_06264_));
 sky130_fd_sc_hd__nor3_1 _17539_ (.A(_06263_),
    .B(_06264_),
    .C(_06239_),
    .Y(_06265_));
 sky130_fd_sc_hd__a211o_1 _17540_ (.A1(_13493_),
    .A2(_13485_),
    .B1(_13492_),
    .C1(_13478_),
    .X(_06266_));
 sky130_fd_sc_hd__and4_1 _17541_ (.A(_13458_),
    .B(_13465_),
    .C(_13472_),
    .D(_13450_),
    .X(_06267_));
 sky130_fd_sc_hd__a2111o_2 _17542_ (.A1(_13472_),
    .A2(_06247_),
    .B1(_06266_),
    .C1(_06267_),
    .D1(_13471_),
    .X(_06268_));
 sky130_fd_sc_hd__o211ai_1 _17543_ (.A1(_13479_),
    .A2(_13478_),
    .B1(_13493_),
    .C1(_13486_),
    .Y(_06269_));
 sky130_fd_sc_hd__a21oi_1 _17544_ (.A1(_13493_),
    .A2(_13485_),
    .B1(_13492_),
    .Y(_06270_));
 sky130_fd_sc_hd__nand2_2 _17545_ (.A(_06269_),
    .B(_06270_),
    .Y(_06271_));
 sky130_fd_sc_hd__o21ai_2 _17546_ (.A1(_06265_),
    .A2(_06268_),
    .B1(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__xnor2_4 _17547_ (.A(_13500_),
    .B(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nor2_4 _17548_ (.A(net524),
    .B(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__inv_1 _17549_ (.A(_06274_),
    .Y(\hash.CA1.S0.X[14] ));
 sky130_fd_sc_hd__and3_1 _17550_ (.A(\hash.CA1.S0.X[11] ),
    .B(\hash.CA1.S0.X[12] ),
    .C(_06252_),
    .X(_06275_));
 sky130_fd_sc_hd__nor2_1 _17551_ (.A(\hash.CA1.S0.X[13] ),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__xnor2_1 _17552_ (.A(_06274_),
    .B(_06276_),
    .Y(_00663_));
 sky130_fd_sc_hd__nand2_1 _17553_ (.A(_13493_),
    .B(_13500_),
    .Y(_06277_));
 sky130_fd_sc_hd__nor3_2 _17554_ (.A(_06239_),
    .B(_06255_),
    .C(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__o21ai_4 _17555_ (.A1(_06202_),
    .A2(_06203_),
    .B1(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__a31oi_4 _17556_ (.A1(_13500_),
    .A2(_06271_),
    .A3(_06268_),
    .B1(_13499_),
    .Y(_06280_));
 sky130_fd_sc_hd__nand2_1 _17557_ (.A(_06279_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__xor2_1 _17558_ (.A(_13507_),
    .B(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__nor2_4 _17559_ (.A(net524),
    .B(_06282_),
    .Y(_06283_));
 sky130_fd_sc_hd__inv_1 _17560_ (.A(_06283_),
    .Y(\hash.CA1.S0.X[15] ));
 sky130_fd_sc_hd__nand3_1 _17561_ (.A(_06259_),
    .B(_06260_),
    .C(_06274_),
    .Y(_06284_));
 sky130_fd_sc_hd__xnor2_1 _17562_ (.A(\hash.CA1.S0.X[15] ),
    .B(_06284_),
    .Y(_00664_));
 sky130_fd_sc_hd__nor2b_1 _17563_ (.A(net524),
    .B_N(_13514_),
    .Y(_06285_));
 sky130_fd_sc_hd__nor2_1 _17564_ (.A(net524),
    .B(_13514_),
    .Y(_06286_));
 sky130_fd_sc_hd__nand2_1 _17565_ (.A(_13500_),
    .B(_06271_),
    .Y(_06287_));
 sky130_fd_sc_hd__or4_4 _17566_ (.A(_06263_),
    .B(_06264_),
    .C(_06239_),
    .D(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__nand2_1 _17567_ (.A(_06288_),
    .B(_06280_),
    .Y(_06289_));
 sky130_fd_sc_hd__a21oi_1 _17568_ (.A1(_13507_),
    .A2(_06289_),
    .B1(_13506_),
    .Y(_06290_));
 sky130_fd_sc_hd__mux2_4 _17569_ (.A0(_06285_),
    .A1(_06286_),
    .S(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__inv_1 _17570_ (.A(_06291_),
    .Y(\hash.CA1.S0.X[16] ));
 sky130_fd_sc_hd__nor4_4 _17571_ (.A(net524),
    .B(_06258_),
    .C(_06273_),
    .D(\hash.CA1.S0.X[15] ),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2b_1 _17572_ (.A_N(_06275_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__xnor2_1 _17573_ (.A(\hash.CA1.S0.X[16] ),
    .B(_06293_),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_1 _17574_ (.A(_13513_),
    .Y(_06294_));
 sky130_fd_sc_hd__a21boi_0 _17575_ (.A1(_06279_),
    .A2(_06280_),
    .B1_N(_13507_),
    .Y(_06295_));
 sky130_fd_sc_hd__o21ai_1 _17576_ (.A1(_13506_),
    .A2(_06295_),
    .B1(_13514_),
    .Y(_06296_));
 sky130_fd_sc_hd__a21oi_2 _17577_ (.A1(_06294_),
    .A2(_06296_),
    .B1(_13521_),
    .Y(_06297_));
 sky130_fd_sc_hd__and3_1 _17578_ (.A(_13521_),
    .B(_06294_),
    .C(_06296_),
    .X(_06298_));
 sky130_fd_sc_hd__nor2_1 _17579_ (.A(_06297_),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__nor2_4 _17580_ (.A(net524),
    .B(_06299_),
    .Y(\hash.CA1.S0.X[17] ));
 sky130_fd_sc_hd__nand3_1 _17581_ (.A(_06260_),
    .B(_06291_),
    .C(_06292_),
    .Y(_06300_));
 sky130_fd_sc_hd__xor2_1 _17582_ (.A(\hash.CA1.S0.X[17] ),
    .B(_06300_),
    .X(_00666_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1181 ();
 sky130_fd_sc_hd__and2_0 _17586_ (.A(_13514_),
    .B(_13521_),
    .X(_06304_));
 sky130_fd_sc_hd__nand2_1 _17587_ (.A(_13507_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__a21oi_1 _17588_ (.A1(_06288_),
    .A2(_06280_),
    .B1(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__a21oi_1 _17589_ (.A1(_13521_),
    .A2(_13513_),
    .B1(_13520_),
    .Y(_06307_));
 sky130_fd_sc_hd__nand3_1 _17590_ (.A(_13514_),
    .B(_13521_),
    .C(_13506_),
    .Y(_06308_));
 sky130_fd_sc_hd__nand2_1 _17591_ (.A(_06307_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__o21ai_2 _17592_ (.A1(_06306_),
    .A2(_06309_),
    .B1(_13528_),
    .Y(_06310_));
 sky130_fd_sc_hd__or3_1 _17593_ (.A(_13528_),
    .B(_06306_),
    .C(_06309_),
    .X(_06311_));
 sky130_fd_sc_hd__and3_4 _17594_ (.A(net519),
    .B(_06310_),
    .C(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1178 ();
 sky130_fd_sc_hd__nor3b_1 _17598_ (.A(_06275_),
    .B(\hash.CA1.S0.X[16] ),
    .C_N(_06292_),
    .Y(_06315_));
 sky130_fd_sc_hd__nor3_1 _17599_ (.A(net524),
    .B(_06299_),
    .C(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__xor2_1 _17600_ (.A(_06312_),
    .B(_06316_),
    .X(_00667_));
 sky130_fd_sc_hd__o21ai_0 _17601_ (.A1(_13506_),
    .A2(_06295_),
    .B1(_06304_),
    .Y(_06317_));
 sky130_fd_sc_hd__a21boi_0 _17602_ (.A1(_06307_),
    .A2(_06317_),
    .B1_N(_13528_),
    .Y(_06318_));
 sky130_fd_sc_hd__o21a_1 _17603_ (.A1(_13527_),
    .A2(_06318_),
    .B1(_13535_),
    .X(_06319_));
 sky130_fd_sc_hd__nor3_1 _17604_ (.A(_13535_),
    .B(_13527_),
    .C(_06318_),
    .Y(_06320_));
 sky130_fd_sc_hd__o21a_4 _17605_ (.A1(_06319_),
    .A2(_06320_),
    .B1(net519),
    .X(_06321_));
 sky130_fd_sc_hd__clkinv_2 _17606_ (.A(_06321_),
    .Y(\hash.CA1.S0.X[19] ));
 sky130_fd_sc_hd__o2111ai_4 _17607_ (.A1(_06297_),
    .A2(_06298_),
    .B1(_06310_),
    .C1(_06311_),
    .D1(net519),
    .Y(_06322_));
 sky130_fd_sc_hd__a31oi_4 _17608_ (.A1(_06260_),
    .A2(_06291_),
    .A3(_06292_),
    .B1(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__xnor2_1 _17609_ (.A(\hash.CA1.S0.X[19] ),
    .B(_06323_),
    .Y(_00668_));
 sky130_fd_sc_hd__a21o_1 _17610_ (.A1(_13535_),
    .A2(_13527_),
    .B1(_13534_),
    .X(_06324_));
 sky130_fd_sc_hd__a31o_1 _17611_ (.A1(_13528_),
    .A2(_13535_),
    .A3(_06309_),
    .B1(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__nand2_2 _17612_ (.A(_13542_),
    .B(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__and3_1 _17613_ (.A(_13528_),
    .B(_13535_),
    .C(_06304_),
    .X(_06327_));
 sky130_fd_sc_hd__and3_1 _17614_ (.A(_13542_),
    .B(_13507_),
    .C(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a21bo_4 _17615_ (.A1(_06288_),
    .A2(_06280_),
    .B1_N(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__nand3_1 _17616_ (.A(net519),
    .B(_06326_),
    .C(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__a311o_1 _17617_ (.A1(_13507_),
    .A2(_06289_),
    .A3(_06327_),
    .B1(_06325_),
    .C1(_13542_),
    .X(_06331_));
 sky130_fd_sc_hd__nand2b_2 _17618_ (.A_N(_06330_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__clkinv_4 _17619_ (.A(_06332_),
    .Y(\hash.CA1.S0.X[20] ));
 sky130_fd_sc_hd__o21a_2 _17620_ (.A1(_06315_),
    .A2(_06322_),
    .B1(_06321_),
    .X(_06333_));
 sky130_fd_sc_hd__xnor2_1 _17621_ (.A(\hash.CA1.S0.X[20] ),
    .B(_06333_),
    .Y(_00670_));
 sky130_fd_sc_hd__and2_0 _17622_ (.A(_13542_),
    .B(_06325_),
    .X(_06334_));
 sky130_fd_sc_hd__a21boi_4 _17623_ (.A1(_06280_),
    .A2(_06279_),
    .B1_N(_06328_),
    .Y(_06335_));
 sky130_fd_sc_hd__nor3_2 _17624_ (.A(_13541_),
    .B(_06334_),
    .C(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__xnor2_4 _17625_ (.A(_13549_),
    .B(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__and2_2 _17626_ (.A(net519),
    .B(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1177 ();
 sky130_fd_sc_hd__nor2_1 _17628_ (.A(\hash.CA1.S0.X[19] ),
    .B(_06323_),
    .Y(_06339_));
 sky130_fd_sc_hd__nor2_1 _17629_ (.A(_06339_),
    .B(_06332_),
    .Y(_06340_));
 sky130_fd_sc_hd__xor2_1 _17630_ (.A(_06338_),
    .B(_06340_),
    .X(_00671_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1175 ();
 sky130_fd_sc_hd__inv_1 _17633_ (.A(_13541_),
    .Y(_06343_));
 sky130_fd_sc_hd__inv_1 _17634_ (.A(_13549_),
    .Y(_06344_));
 sky130_fd_sc_hd__a31oi_1 _17635_ (.A1(_06343_),
    .A2(_06326_),
    .A3(_06329_),
    .B1(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__nor2_1 _17636_ (.A(_13541_),
    .B(_13548_),
    .Y(_06346_));
 sky130_fd_sc_hd__o21ai_2 _17637_ (.A1(_13549_),
    .A2(_13548_),
    .B1(_13556_),
    .Y(_06347_));
 sky130_fd_sc_hd__a31o_1 _17638_ (.A1(_06326_),
    .A2(_06329_),
    .A3(_06346_),
    .B1(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__o31a_4 _17639_ (.A1(_13556_),
    .A2(_13548_),
    .A3(_06345_),
    .B1(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1174 ();
 sky130_fd_sc_hd__and2_0 _17641_ (.A(net519),
    .B(_06349_),
    .X(\hash.CA1.S0.X[22] ));
 sky130_fd_sc_hd__nand2_1 _17642_ (.A(\hash.CA1.S0.X[20] ),
    .B(_06338_),
    .Y(_06351_));
 sky130_fd_sc_hd__nor2_1 _17643_ (.A(_06333_),
    .B(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__xor2_1 _17644_ (.A(\hash.CA1.S0.X[22] ),
    .B(_06352_),
    .X(_00672_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1173 ();
 sky130_fd_sc_hd__o21a_1 _17646_ (.A1(_13549_),
    .A2(_13548_),
    .B1(_13556_),
    .X(_06354_));
 sky130_fd_sc_hd__o41a_1 _17647_ (.A1(_13541_),
    .A2(_13548_),
    .A3(_06334_),
    .A4(_06335_),
    .B1(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__nor3_1 _17648_ (.A(_13563_),
    .B(_13555_),
    .C(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__o21a_1 _17649_ (.A1(_13555_),
    .A2(_06355_),
    .B1(_13563_),
    .X(_06357_));
 sky130_fd_sc_hd__nor3_4 _17650_ (.A(net521),
    .B(_06356_),
    .C(_06357_),
    .Y(\hash.CA1.S0.X[23] ));
 sky130_fd_sc_hd__nand3_1 _17651_ (.A(\hash.CA1.S0.X[20] ),
    .B(_06338_),
    .C(_06349_),
    .Y(_06358_));
 sky130_fd_sc_hd__nor2_1 _17652_ (.A(_06339_),
    .B(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__xor2_1 _17653_ (.A(\hash.CA1.S0.X[23] ),
    .B(_06359_),
    .X(_00673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1172 ();
 sky130_fd_sc_hd__nor2b_1 _17655_ (.A(_13570_),
    .B_N(_13563_),
    .Y(_06361_));
 sky130_fd_sc_hd__inv_1 _17656_ (.A(_13570_),
    .Y(_06362_));
 sky130_fd_sc_hd__nor3_1 _17657_ (.A(_06362_),
    .B(_13555_),
    .C(_13562_),
    .Y(_06363_));
 sky130_fd_sc_hd__mux2i_1 _17658_ (.A0(_06361_),
    .A1(_06363_),
    .S(_06348_),
    .Y(_06364_));
 sky130_fd_sc_hd__nor3_1 _17659_ (.A(_13563_),
    .B(_06362_),
    .C(_13562_),
    .Y(_06365_));
 sky130_fd_sc_hd__a221oi_1 _17660_ (.A1(_06362_),
    .A2(_13562_),
    .B1(_06361_),
    .B2(_13555_),
    .C1(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__and2_4 _17661_ (.A(_06364_),
    .B(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nor2_8 _17662_ (.A(net524),
    .B(_06367_),
    .Y(\hash.CA1.S0.X[24] ));
 sky130_fd_sc_hd__and4_1 _17663_ (.A(\hash.CA1.S0.X[20] ),
    .B(_06338_),
    .C(_06349_),
    .D(\hash.CA1.S0.X[23] ),
    .X(_06368_));
 sky130_fd_sc_hd__nand2b_1 _17664_ (.A_N(_06333_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__xnor2_1 _17665_ (.A(\hash.CA1.S0.X[24] ),
    .B(_06369_),
    .Y(_00674_));
 sky130_fd_sc_hd__o21ai_2 _17666_ (.A1(_13562_),
    .A2(_06357_),
    .B1(_13570_),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_1 _17667_ (.A(_13577_),
    .B(_13569_),
    .Y(_06371_));
 sky130_fd_sc_hd__o2111ai_2 _17668_ (.A1(_13555_),
    .A2(_06355_),
    .B1(_13563_),
    .C1(_13570_),
    .D1(_13577_),
    .Y(_06372_));
 sky130_fd_sc_hd__a21o_1 _17669_ (.A1(_13570_),
    .A2(_13562_),
    .B1(_13569_),
    .X(_06373_));
 sky130_fd_sc_hd__nand2_1 _17670_ (.A(_13577_),
    .B(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_2 _17671_ (.A(_06372_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__a21oi_4 _17672_ (.A1(_06370_),
    .A2(_06371_),
    .B1(_06375_),
    .Y(_06376_));
 sky130_fd_sc_hd__nor2_8 _17673_ (.A(net521),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__inv_4 _17674_ (.A(_06377_),
    .Y(\hash.CA1.S0.X[25] ));
 sky130_fd_sc_hd__nand2_1 _17675_ (.A(_06364_),
    .B(_06366_),
    .Y(_06378_));
 sky130_fd_sc_hd__o211ai_4 _17676_ (.A1(\hash.CA1.S0.X[19] ),
    .A2(_06323_),
    .B1(_06378_),
    .C1(_06368_),
    .Y(_06379_));
 sky130_fd_sc_hd__xnor2_1 _17677_ (.A(_06377_),
    .B(_06379_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_1 _17678_ (.A(_13563_),
    .B(_13570_),
    .Y(_06380_));
 sky130_fd_sc_hd__a311oi_4 _17679_ (.A1(_06326_),
    .A2(_06329_),
    .A3(_06346_),
    .B1(_06380_),
    .C1(_06347_),
    .Y(_06381_));
 sky130_fd_sc_hd__a21oi_1 _17680_ (.A1(_13563_),
    .A2(_13555_),
    .B1(_13562_),
    .Y(_06382_));
 sky130_fd_sc_hd__nor2_1 _17681_ (.A(_06362_),
    .B(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__nor2_1 _17682_ (.A(_13569_),
    .B(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__inv_1 _17683_ (.A(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__inv_1 _17684_ (.A(_13576_),
    .Y(_06386_));
 sky130_fd_sc_hd__nand3_1 _17685_ (.A(net519),
    .B(_13584_),
    .C(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__inv_1 _17686_ (.A(_13584_),
    .Y(_06388_));
 sky130_fd_sc_hd__and3_1 _17687_ (.A(net519),
    .B(_13577_),
    .C(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nand2_1 _17688_ (.A(_06381_),
    .B(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__nor2_1 _17689_ (.A(net521),
    .B(_13584_),
    .Y(_06391_));
 sky130_fd_sc_hd__nor4_1 _17690_ (.A(net521),
    .B(_13577_),
    .C(_06388_),
    .D(_13576_),
    .Y(_06392_));
 sky130_fd_sc_hd__a221oi_2 _17691_ (.A1(_06385_),
    .A2(_06389_),
    .B1(_06391_),
    .B2(_13576_),
    .C1(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__o311ai_4 _17692_ (.A1(_06381_),
    .A2(_06385_),
    .A3(_06387_),
    .B1(_06390_),
    .C1(_06393_),
    .Y(\hash.CA1.S0.X[26] ));
 sky130_fd_sc_hd__inv_2 _17693_ (.A(_06368_),
    .Y(_06394_));
 sky130_fd_sc_hd__o31ai_2 _17694_ (.A1(_06333_),
    .A2(_06367_),
    .A3(_06394_),
    .B1(_06377_),
    .Y(_06395_));
 sky130_fd_sc_hd__xor2_1 _17695_ (.A(\hash.CA1.S0.X[26] ),
    .B(_06395_),
    .X(_00676_));
 sky130_fd_sc_hd__nor2_1 _17696_ (.A(_13576_),
    .B(_13583_),
    .Y(_06396_));
 sky130_fd_sc_hd__o21ai_0 _17697_ (.A1(_13584_),
    .A2(_13583_),
    .B1(_13591_),
    .Y(_06397_));
 sky130_fd_sc_hd__a31oi_1 _17698_ (.A1(_06372_),
    .A2(_06374_),
    .A3(_06396_),
    .B1(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__inv_1 _17699_ (.A(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__a31oi_1 _17700_ (.A1(_06372_),
    .A2(_06386_),
    .A3(_06374_),
    .B1(_06388_),
    .Y(_06400_));
 sky130_fd_sc_hd__or3_4 _17701_ (.A(_13591_),
    .B(_13583_),
    .C(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__a21oi_4 _17702_ (.A1(_06399_),
    .A2(_06401_),
    .B1(net521),
    .Y(_06402_));
 sky130_fd_sc_hd__clkinv_2 _17703_ (.A(_06402_),
    .Y(\hash.CA1.S0.X[27] ));
 sky130_fd_sc_hd__nor3_1 _17704_ (.A(_06339_),
    .B(_06367_),
    .C(_06394_),
    .Y(_06403_));
 sky130_fd_sc_hd__o21ai_0 _17705_ (.A1(\hash.CA1.S0.X[25] ),
    .A2(_06403_),
    .B1(\hash.CA1.S0.X[26] ),
    .Y(_06404_));
 sky130_fd_sc_hd__xnor2_1 _17706_ (.A(_06402_),
    .B(_06404_),
    .Y(_00677_));
 sky130_fd_sc_hd__a21oi_1 _17707_ (.A1(_13591_),
    .A2(_13583_),
    .B1(_13590_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand3_1 _17708_ (.A(_06386_),
    .B(_06384_),
    .C(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand2_1 _17709_ (.A(_13584_),
    .B(_13591_),
    .Y(_06407_));
 sky130_fd_sc_hd__nor2_1 _17710_ (.A(_13577_),
    .B(_13576_),
    .Y(_06408_));
 sky130_fd_sc_hd__o21ai_0 _17711_ (.A1(_06407_),
    .A2(_06408_),
    .B1(_06405_),
    .Y(_06409_));
 sky130_fd_sc_hd__o21ai_2 _17712_ (.A1(_06381_),
    .A2(_06406_),
    .B1(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__xnor2_4 _17713_ (.A(_13598_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_8 _17714_ (.A(net519),
    .B(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__inv_1 _17715_ (.A(_06412_),
    .Y(\hash.CA1.S0.X[28] ));
 sky130_fd_sc_hd__a21oi_1 _17716_ (.A1(\hash.CA1.S0.X[26] ),
    .A2(_06395_),
    .B1(\hash.CA1.S0.X[27] ),
    .Y(_06413_));
 sky130_fd_sc_hd__xnor2_1 _17717_ (.A(\hash.CA1.S0.X[28] ),
    .B(_06413_),
    .Y(_00678_));
 sky130_fd_sc_hd__o21a_1 _17718_ (.A1(_13590_),
    .A2(_06398_),
    .B1(_13598_),
    .X(_06414_));
 sky130_fd_sc_hd__nor2_2 _17719_ (.A(_13597_),
    .B(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__xnor2_4 _17720_ (.A(_13605_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__nor2_8 _17721_ (.A(net521),
    .B(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__clkinv_2 _17722_ (.A(_06417_),
    .Y(\hash.CA1.S0.X[29] ));
 sky130_fd_sc_hd__a211oi_2 _17723_ (.A1(_06399_),
    .A2(_06401_),
    .B1(net521),
    .C1(\hash.CA1.S0.X[26] ),
    .Y(_06418_));
 sky130_fd_sc_hd__a311oi_4 _17724_ (.A1(_06377_),
    .A2(_06379_),
    .A3(_06402_),
    .B1(_06412_),
    .C1(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__xor2_1 _17725_ (.A(_06417_),
    .B(_06419_),
    .X(_00679_));
 sky130_fd_sc_hd__nor2_1 _17726_ (.A(net521),
    .B(_13612_),
    .Y(_06420_));
 sky130_fd_sc_hd__nor2b_1 _17727_ (.A(net521),
    .B_N(_13612_),
    .Y(_06421_));
 sky130_fd_sc_hd__o21a_1 _17728_ (.A1(_06381_),
    .A2(_06385_),
    .B1(_13577_),
    .X(_06422_));
 sky130_fd_sc_hd__nor2_1 _17729_ (.A(_13576_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__nand4_1 _17730_ (.A(_13584_),
    .B(_13591_),
    .C(_13598_),
    .D(_13605_),
    .Y(_06424_));
 sky130_fd_sc_hd__inv_1 _17731_ (.A(_13598_),
    .Y(_06425_));
 sky130_fd_sc_hd__o21bai_1 _17732_ (.A1(_06425_),
    .A2(_06405_),
    .B1_N(_13597_),
    .Y(_06426_));
 sky130_fd_sc_hd__a21oi_1 _17733_ (.A1(_13605_),
    .A2(_06426_),
    .B1(_13604_),
    .Y(_06427_));
 sky130_fd_sc_hd__o21ai_2 _17734_ (.A1(_06423_),
    .A2(_06424_),
    .B1(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__mux2i_4 _17735_ (.A0(_06420_),
    .A1(_06421_),
    .S(_06428_),
    .Y(\hash.CA1.S0.X[30] ));
 sky130_fd_sc_hd__o21ai_0 _17736_ (.A1(_06412_),
    .A2(_06413_),
    .B1(_06417_),
    .Y(_06429_));
 sky130_fd_sc_hd__xnor2_1 _17737_ (.A(\hash.CA1.S0.X[30] ),
    .B(_06429_),
    .Y(_00681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1171 ();
 sky130_fd_sc_hd__mux2i_4 _17739_ (.A0(\hash.CA2.f_dash[31] ),
    .A1(\hash.CA2.e_dash[31] ),
    .S(\hash.CA2.S1.X[31] ),
    .Y(_06431_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1168 ();
 sky130_fd_sc_hd__xor2_4 _17743_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA2.S1.X[5] ),
    .X(_06435_));
 sky130_fd_sc_hd__xnor2_2 _17744_ (.A(\hash.CA2.S1.X[24] ),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__xnor2_4 _17745_ (.A(_06431_),
    .B(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__nand3_1 _17746_ (.A(_13595_),
    .B(_13602_),
    .C(_13609_),
    .Y(_06438_));
 sky130_fd_sc_hd__a21o_1 _17747_ (.A1(_13595_),
    .A2(_13587_),
    .B1(_13594_),
    .X(_06439_));
 sky130_fd_sc_hd__a21o_1 _17748_ (.A1(_13602_),
    .A2(_06439_),
    .B1(_13601_),
    .X(_06440_));
 sky130_fd_sc_hd__a21oi_1 _17749_ (.A1(_13609_),
    .A2(_06440_),
    .B1(_13608_),
    .Y(_06441_));
 sky130_fd_sc_hd__nand2_1 _17750_ (.A(_06437_),
    .B(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__a211o_1 _17751_ (.A1(_04930_),
    .A2(_04970_),
    .B1(_04971_),
    .C1(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__nand3_1 _17752_ (.A(_06437_),
    .B(_06441_),
    .C(_06438_),
    .Y(_06444_));
 sky130_fd_sc_hd__o21a_1 _17753_ (.A1(_06437_),
    .A2(_06441_),
    .B1(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__o311ai_4 _17754_ (.A1(_04972_),
    .A2(_06437_),
    .A3(_06438_),
    .B1(_06443_),
    .C1(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__xnor2_1 _17755_ (.A(\hash.CA2.p4[31] ),
    .B(_12532_),
    .Y(_06447_));
 sky130_fd_sc_hd__xnor2_1 _17756_ (.A(_12253_),
    .B(_12528_),
    .Y(_06448_));
 sky130_fd_sc_hd__xnor2_1 _17757_ (.A(_06447_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__xnor2_1 _17758_ (.A(_04786_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__xnor2_1 _17759_ (.A(net1160),
    .B(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__inv_1 _17760_ (.A(_13611_),
    .Y(_06452_));
 sky130_fd_sc_hd__nand3_1 _17761_ (.A(_06386_),
    .B(_06452_),
    .C(_06427_),
    .Y(_06453_));
 sky130_fd_sc_hd__nor2_1 _17762_ (.A(_13612_),
    .B(_13611_),
    .Y(_06454_));
 sky130_fd_sc_hd__a31oi_1 _17763_ (.A1(_06452_),
    .A2(_06427_),
    .A3(_06424_),
    .B1(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__o21ai_2 _17764_ (.A1(_06453_),
    .A2(_06375_),
    .B1(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__xnor2_2 _17765_ (.A(_06451_),
    .B(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__xnor2_4 _17766_ (.A(_06446_),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__or2_1 _17767_ (.A(\hash.CA2.a_dash[31] ),
    .B(_04805_),
    .X(_06459_));
 sky130_fd_sc_hd__and2_1 _17768_ (.A(\hash.CA2.a_dash[31] ),
    .B(_04805_),
    .X(_06460_));
 sky130_fd_sc_hd__a21oi_2 _17769_ (.A1(\hash.CA2.b_dash[31] ),
    .A2(_06459_),
    .B1(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__xnor2_4 _17770_ (.A(_06458_),
    .B(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__nor2_1 _17771_ (.A(net521),
    .B(_06462_),
    .Y(\hash.CA1.S0.X[31] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1166 ();
 sky130_fd_sc_hd__nor3_1 _17774_ (.A(_06416_),
    .B(_06419_),
    .C(\hash.CA1.S0.X[30] ),
    .Y(_06465_));
 sky130_fd_sc_hd__xnor2_1 _17775_ (.A(_06462_),
    .B(_06465_),
    .Y(_06466_));
 sky130_fd_sc_hd__nand2_1 _17776_ (.A(net519),
    .B(_06466_),
    .Y(_00682_));
 sky130_fd_sc_hd__xnor2_2 _17777_ (.A(\hash.CA1.S0.X[3] ),
    .B(_06274_),
    .Y(_06467_));
 sky130_fd_sc_hd__xor2_4 _17778_ (.A(net1127),
    .B(_06467_),
    .X(_13716_));
 sky130_fd_sc_hd__inv_1 _17779_ (.A(_13716_),
    .Y(_13052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1165 ();
 sky130_fd_sc_hd__nor2b_1 _17781_ (.A(net520),
    .B_N(_12253_),
    .Y(\hash.CA1.b[1] ));
 sky130_fd_sc_hd__a21oi_1 _17782_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_13409_),
    .B1(_12253_),
    .Y(_06469_));
 sky130_fd_sc_hd__nor2_1 _17783_ (.A(\hash.CA2.a_dash[1] ),
    .B(_13409_),
    .Y(_06470_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1164 ();
 sky130_fd_sc_hd__o21ai_0 _17785_ (.A1(_06469_),
    .A2(_06470_),
    .B1(net519),
    .Y(_13715_));
 sky130_fd_sc_hd__inv_1 _17786_ (.A(_13715_),
    .Y(_13051_));
 sky130_fd_sc_hd__nor2b_1 _17787_ (.A(net520),
    .B_N(\hash.CA2.a_dash[0] ),
    .Y(\hash.CA1.c[0] ));
 sky130_fd_sc_hd__nand2_1 _17788_ (.A(net519),
    .B(_04840_),
    .Y(\hash.CA1.b[2] ));
 sky130_fd_sc_hd__nor2b_1 _17789_ (.A(net520),
    .B_N(\hash.CA2.a_dash[2] ),
    .Y(_13841_));
 sky130_fd_sc_hd__nor2_1 _17790_ (.A(net520),
    .B(_04646_),
    .Y(\hash.CA1.b[3] ));
 sky130_fd_sc_hd__nor2_2 _17791_ (.A(net520),
    .B(_04662_),
    .Y(_13847_));
 sky130_fd_sc_hd__and2_0 _17792_ (.A(_06210_),
    .B(_04654_),
    .X(\hash.CA1.b[4] ));
 sky130_fd_sc_hd__and2_0 _17793_ (.A(net519),
    .B(_04674_),
    .X(\hash.CA1.b[5] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1163 ();
 sky130_fd_sc_hd__or2_0 _17795_ (.A(net520),
    .B(\hash.CA2.a_dash[5] ),
    .X(_13859_));
 sky130_fd_sc_hd__and2_1 _17796_ (.A(net519),
    .B(_04701_),
    .X(\hash.CA1.b[6] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1162 ();
 sky130_fd_sc_hd__or2_1 _17798_ (.A(net520),
    .B(\hash.CA2.a_dash[6] ),
    .X(_13865_));
 sky130_fd_sc_hd__inv_1 _17799_ (.A(_04724_),
    .Y(_06474_));
 sky130_fd_sc_hd__nand2_1 _17800_ (.A(net519),
    .B(_06474_),
    .Y(\hash.CA1.b[7] ));
 sky130_fd_sc_hd__and2_0 _17801_ (.A(net519),
    .B(_04742_),
    .X(\hash.CA1.b[8] ));
 sky130_fd_sc_hd__nand2_1 _17802_ (.A(net519),
    .B(_04895_),
    .Y(\hash.CA1.b[9] ));
 sky130_fd_sc_hd__nor2_1 _17803_ (.A(net520),
    .B(\hash.CA2.a_dash[9] ),
    .Y(_06475_));
 sky130_fd_sc_hd__inv_1 _17804_ (.A(_06475_),
    .Y(_13884_));
 sky130_fd_sc_hd__o21ai_1 _17805_ (.A1(_04788_),
    .A2(_04790_),
    .B1(_06210_),
    .Y(\hash.CA1.b[10] ));
 sky130_fd_sc_hd__nand2_1 _17806_ (.A(net519),
    .B(_04813_),
    .Y(\hash.CA1.b[11] ));
 sky130_fd_sc_hd__nor2_4 _17807_ (.A(net524),
    .B(net1163),
    .Y(\hash.CA1.b[12] ));
 sky130_fd_sc_hd__nand2_1 _17808_ (.A(net519),
    .B(_04611_),
    .Y(\hash.CA1.b[13] ));
 sky130_fd_sc_hd__or2_0 _17809_ (.A(net524),
    .B(\hash.CA2.a_dash[13] ),
    .X(_13908_));
 sky130_fd_sc_hd__and2_0 _17810_ (.A(net519),
    .B(_04627_),
    .X(\hash.CA1.b[14] ));
 sky130_fd_sc_hd__nor2_1 _17811_ (.A(net524),
    .B(\hash.CA2.a_dash[14] ),
    .Y(_06476_));
 sky130_fd_sc_hd__inv_1 _17812_ (.A(_06476_),
    .Y(_13914_));
 sky130_fd_sc_hd__o21ai_4 _17813_ (.A1(_04657_),
    .A2(_04658_),
    .B1(_06210_),
    .Y(\hash.CA1.b[15] ));
 sky130_fd_sc_hd__or2_2 _17814_ (.A(net524),
    .B(\hash.CA2.a_dash[15] ),
    .X(_13921_));
 sky130_fd_sc_hd__nand2_1 _17815_ (.A(net519),
    .B(net1130),
    .Y(\hash.CA1.b[16] ));
 sky130_fd_sc_hd__nor2_1 _17816_ (.A(net524),
    .B(_04699_),
    .Y(_06477_));
 sky130_fd_sc_hd__inv_1 _17817_ (.A(_06477_),
    .Y(\hash.CA1.b[17] ));
 sky130_fd_sc_hd__or2_0 _17818_ (.A(net524),
    .B(_04721_),
    .X(\hash.CA1.b[18] ));
 sky130_fd_sc_hd__nor2_1 _17819_ (.A(net524),
    .B(_04740_),
    .Y(\hash.CA1.b[19] ));
 sky130_fd_sc_hd__or2_1 _17820_ (.A(net521),
    .B(\hash.CA2.a_dash[19] ),
    .X(_13946_));
 sky130_fd_sc_hd__nor2_1 _17821_ (.A(net524),
    .B(net1140),
    .Y(\hash.CA1.b[20] ));
 sky130_fd_sc_hd__or2_2 _17822_ (.A(net521),
    .B(_04786_),
    .X(_06478_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1161 ();
 sky130_fd_sc_hd__or2_0 _17824_ (.A(net524),
    .B(net1122),
    .X(\hash.CA1.b[22] ));
 sky130_fd_sc_hd__and2_2 _17825_ (.A(net519),
    .B(net1168),
    .X(_06479_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1160 ();
 sky130_fd_sc_hd__or2_0 _17827_ (.A(net521),
    .B(_04652_),
    .X(\hash.CA1.b[24] ));
 sky130_fd_sc_hd__or2_0 _17828_ (.A(net524),
    .B(net1164),
    .X(\hash.CA1.b[25] ));
 sky130_fd_sc_hd__nor3_4 _17829_ (.A(net521),
    .B(_04692_),
    .C(net1125),
    .Y(\hash.CA1.b[26] ));
 sky130_fd_sc_hd__or2_1 _17830_ (.A(net521),
    .B(\hash.CA2.a_dash[26] ),
    .X(_06480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1159 ();
 sky130_fd_sc_hd__or2_1 _17832_ (.A(net521),
    .B(_04716_),
    .X(_06481_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1158 ();
 sky130_fd_sc_hd__or2_0 _17834_ (.A(net521),
    .B(\hash.CA2.a_dash[27] ),
    .X(_13995_));
 sky130_fd_sc_hd__or2_0 _17835_ (.A(net521),
    .B(_04736_),
    .X(\hash.CA1.b[28] ));
 sky130_fd_sc_hd__or2_1 _17836_ (.A(net521),
    .B(\hash.CA2.a_dash[28] ),
    .X(_14002_));
 sky130_fd_sc_hd__or2_1 _17837_ (.A(net521),
    .B(\hash.CA2.a_dash[29] ),
    .X(_14008_));
 sky130_fd_sc_hd__nor2_1 _17838_ (.A(net521),
    .B(net1118),
    .Y(\hash.CA1.b[30] ));
 sky130_fd_sc_hd__or2_0 _17839_ (.A(net521),
    .B(_04805_),
    .X(\hash.CA1.b[31] ));
 sky130_fd_sc_hd__nor2_2 _17840_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[1] ),
    .Y(_12539_));
 sky130_fd_sc_hd__nor2b_2 _17841_ (.A(\hash.reset ),
    .B_N(\hash.CA2.e_dash[2] ),
    .Y(_12546_));
 sky130_fd_sc_hd__nor2_1 _17842_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[3] ),
    .Y(_12554_));
 sky130_fd_sc_hd__clkinv_2 _17843_ (.A(\hash.CA2.e_dash[4] ),
    .Y(_06482_));
 sky130_fd_sc_hd__nor2_1 _17844_ (.A(\hash.reset ),
    .B(_06482_),
    .Y(_12557_));
 sky130_fd_sc_hd__nor2_2 _17845_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[5] ),
    .Y(_12562_));
 sky130_fd_sc_hd__nand2_4 _17846_ (.A(_06210_),
    .B(\hash.CA2.e_dash[6] ),
    .Y(_06483_));
 sky130_fd_sc_hd__inv_1 _17847_ (.A(_06483_),
    .Y(_12565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1157 ();
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[7] ),
    .Y(_12570_));
 sky130_fd_sc_hd__nor2_1 _17850_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[8] ),
    .Y(_12575_));
 sky130_fd_sc_hd__nor2b_4 _17851_ (.A(\hash.reset ),
    .B_N(\hash.CA2.e_dash[9] ),
    .Y(_12578_));
 sky130_fd_sc_hd__nor2b_2 _17852_ (.A(net523),
    .B_N(\hash.CA2.e_dash[10] ),
    .Y(_12581_));
 sky130_fd_sc_hd__nor2_4 _17853_ (.A(net523),
    .B(\hash.CA2.e_dash[11] ),
    .Y(_12586_));
 sky130_fd_sc_hd__nor2_2 _17854_ (.A(net523),
    .B(\hash.CA2.e_dash[12] ),
    .Y(_12591_));
 sky130_fd_sc_hd__nor2b_4 _17855_ (.A(net523),
    .B_N(\hash.CA2.e_dash[13] ),
    .Y(_12594_));
 sky130_fd_sc_hd__nor2_4 _17856_ (.A(net523),
    .B(\hash.CA2.e_dash[14] ),
    .Y(_12599_));
 sky130_fd_sc_hd__nor2_4 _17857_ (.A(net523),
    .B(\hash.CA2.e_dash[15] ),
    .Y(_12604_));
 sky130_fd_sc_hd__nor2_2 _17858_ (.A(net523),
    .B(\hash.CA2.e_dash[16] ),
    .Y(_12609_));
 sky130_fd_sc_hd__nor2_4 _17859_ (.A(net523),
    .B(\hash.CA2.e_dash[17] ),
    .Y(_12614_));
 sky130_fd_sc_hd__nor2b_2 _17860_ (.A(net522),
    .B_N(\hash.CA2.e_dash[18] ),
    .Y(_12617_));
 sky130_fd_sc_hd__nand2_1 _17861_ (.A(_06210_),
    .B(\hash.CA2.e_dash[19] ),
    .Y(_06485_));
 sky130_fd_sc_hd__inv_1 _17862_ (.A(_06485_),
    .Y(_12620_));
 sky130_fd_sc_hd__nor2b_2 _17863_ (.A(net522),
    .B_N(\hash.CA2.e_dash[20] ),
    .Y(_12623_));
 sky130_fd_sc_hd__nor2b_2 _17864_ (.A(net522),
    .B_N(\hash.CA2.e_dash[21] ),
    .Y(_12626_));
 sky130_fd_sc_hd__nor2b_1 _17865_ (.A(net522),
    .B_N(\hash.CA2.e_dash[22] ),
    .Y(_12629_));
 sky130_fd_sc_hd__or2_2 _17866_ (.A(net522),
    .B(\hash.CA2.e_dash[23] ),
    .X(_06486_));
 sky130_fd_sc_hd__inv_1 _17867_ (.A(_06486_),
    .Y(_12634_));
 sky130_fd_sc_hd__nor2_1 _17868_ (.A(net522),
    .B(\hash.CA2.e_dash[24] ),
    .Y(_12639_));
 sky130_fd_sc_hd__nor2_1 _17869_ (.A(net522),
    .B(\hash.CA2.e_dash[25] ),
    .Y(_12644_));
 sky130_fd_sc_hd__nor2_2 _17870_ (.A(net522),
    .B(\hash.CA2.e_dash[26] ),
    .Y(_12649_));
 sky130_fd_sc_hd__nor2_2 _17871_ (.A(net522),
    .B(\hash.CA2.e_dash[27] ),
    .Y(_12654_));
 sky130_fd_sc_hd__nor2_1 _17872_ (.A(net522),
    .B(\hash.CA2.e_dash[28] ),
    .Y(_12659_));
 sky130_fd_sc_hd__nor2b_2 _17873_ (.A(net522),
    .B_N(\hash.CA2.e_dash[29] ),
    .Y(_12662_));
 sky130_fd_sc_hd__nor2b_1 _17874_ (.A(net522),
    .B_N(\hash.CA2.e_dash[30] ),
    .Y(_12665_));
 sky130_fd_sc_hd__nor2b_2 _17875_ (.A(\hash.reset ),
    .B_N(\hash.CA2.f_dash[1] ),
    .Y(_12676_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(_06210_),
    .B(\hash.CA2.f_dash[2] ),
    .Y(_12838_));
 sky130_fd_sc_hd__inv_1 _17877_ (.A(_12838_),
    .Y(_12681_));
 sky130_fd_sc_hd__xor2_1 _17878_ (.A(_14016_),
    .B(_12681_),
    .X(_00896_));
 sky130_fd_sc_hd__nor2_1 _17879_ (.A(\hash.reset ),
    .B(\hash.CA2.f_dash[3] ),
    .Y(_12686_));
 sky130_fd_sc_hd__nand3_1 _17880_ (.A(\hash.CA2.f_dash[0] ),
    .B(\hash.CA2.f_dash[1] ),
    .C(\hash.CA2.f_dash[2] ),
    .Y(_06487_));
 sky130_fd_sc_hd__xnor2_1 _17881_ (.A(\hash.CA2.f_dash[3] ),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__nor2_1 _17882_ (.A(\hash.reset ),
    .B(_06488_),
    .Y(_00899_));
 sky130_fd_sc_hd__nor2_2 _17883_ (.A(\hash.reset ),
    .B(\hash.CA2.f_dash[4] ),
    .Y(_12691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1156 ();
 sky130_fd_sc_hd__a211o_1 _17885_ (.A1(\hash.CA2.f_dash[2] ),
    .A2(_14016_),
    .B1(\hash.CA2.f_dash[4] ),
    .C1(\hash.CA2.f_dash[3] ),
    .X(_06490_));
 sky130_fd_sc_hd__a21o_1 _17886_ (.A1(\hash.CA2.f_dash[2] ),
    .A2(_14016_),
    .B1(\hash.CA2.f_dash[3] ),
    .X(_06491_));
 sky130_fd_sc_hd__nand2_1 _17887_ (.A(\hash.CA2.f_dash[4] ),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__nand3_1 _17888_ (.A(_06210_),
    .B(_06490_),
    .C(_06492_),
    .Y(_00900_));
 sky130_fd_sc_hd__nor2b_4 _17889_ (.A(\hash.reset ),
    .B_N(\hash.CA2.f_dash[5] ),
    .Y(_12696_));
 sky130_fd_sc_hd__nand3b_4 _17890_ (.A_N(\hash.CA2.f_dash[3] ),
    .B(_06487_),
    .C(_12691_),
    .Y(_06493_));
 sky130_fd_sc_hd__xor2_4 _17891_ (.A(_12696_),
    .B(_06493_),
    .X(_00901_));
 sky130_fd_sc_hd__nand2_1 _17892_ (.A(_06210_),
    .B(\hash.CA2.f_dash[6] ),
    .Y(_12864_));
 sky130_fd_sc_hd__inv_1 _17893_ (.A(_12864_),
    .Y(_12701_));
 sky130_fd_sc_hd__nand2_1 _17894_ (.A(\hash.CA2.f_dash[5] ),
    .B(_06490_),
    .Y(_06494_));
 sky130_fd_sc_hd__xor2_4 _17895_ (.A(\hash.CA2.f_dash[6] ),
    .B(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__nor2_1 _17896_ (.A(net520),
    .B(_06495_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_2 _17897_ (.A(_06210_),
    .B(\hash.CA2.f_dash[7] ),
    .Y(_12873_));
 sky130_fd_sc_hd__clkinvlp_4 _17898_ (.A(_12873_),
    .Y(_12706_));
 sky130_fd_sc_hd__nand3_2 _17899_ (.A(\hash.CA2.f_dash[6] ),
    .B(_12696_),
    .C(_06493_),
    .Y(_06496_));
 sky130_fd_sc_hd__xnor2_4 _17900_ (.A(_12706_),
    .B(_06496_),
    .Y(_00903_));
 sky130_fd_sc_hd__nor2_4 _17901_ (.A(\hash.reset ),
    .B(\hash.CA2.f_dash[8] ),
    .Y(_12711_));
 sky130_fd_sc_hd__and4_2 _17902_ (.A(\hash.CA2.f_dash[6] ),
    .B(\hash.CA2.f_dash[7] ),
    .C(_06490_),
    .D(_12696_),
    .X(_06497_));
 sky130_fd_sc_hd__xor2_4 _17903_ (.A(_12711_),
    .B(_06497_),
    .X(_00904_));
 sky130_fd_sc_hd__nand2_1 _17904_ (.A(_06210_),
    .B(\hash.CA2.f_dash[9] ),
    .Y(_12886_));
 sky130_fd_sc_hd__inv_1 _17905_ (.A(_12886_),
    .Y(_12716_));
 sky130_fd_sc_hd__a41oi_4 _17906_ (.A1(\hash.CA2.f_dash[6] ),
    .A2(\hash.CA2.f_dash[7] ),
    .A3(_12696_),
    .A4(_06493_),
    .B1(\hash.CA2.f_dash[8] ),
    .Y(_06498_));
 sky130_fd_sc_hd__xor2_1 _17907_ (.A(\hash.CA2.f_dash[9] ),
    .B(_06498_),
    .X(_06499_));
 sky130_fd_sc_hd__nand2_1 _17908_ (.A(net519),
    .B(_06499_),
    .Y(_00905_));
 sky130_fd_sc_hd__nor2_2 _17909_ (.A(\hash.reset ),
    .B(\hash.CA2.f_dash[10] ),
    .Y(_12721_));
 sky130_fd_sc_hd__o21a_1 _17910_ (.A1(\hash.CA2.f_dash[8] ),
    .A2(_06497_),
    .B1(_12716_),
    .X(_06500_));
 sky130_fd_sc_hd__mux2_2 _17911_ (.A0(_12721_),
    .A1(\hash.CA2.f_dash[10] ),
    .S(_06500_),
    .X(_00876_));
 sky130_fd_sc_hd__nor2_1 _17912_ (.A(net523),
    .B(\hash.CA2.f_dash[11] ),
    .Y(_12726_));
 sky130_fd_sc_hd__clkinv_2 _17913_ (.A(_12726_),
    .Y(_12904_));
 sky130_fd_sc_hd__o21ai_1 _17914_ (.A1(_12886_),
    .A2(_06498_),
    .B1(_12721_),
    .Y(_06501_));
 sky130_fd_sc_hd__xnor2_1 _17915_ (.A(_12904_),
    .B(_06501_),
    .Y(_00877_));
 sky130_fd_sc_hd__nor2b_4 _17916_ (.A(net523),
    .B_N(\hash.CA2.f_dash[12] ),
    .Y(_12731_));
 sky130_fd_sc_hd__or3_2 _17917_ (.A(\hash.CA2.f_dash[10] ),
    .B(_06500_),
    .C(_12904_),
    .X(_06502_));
 sky130_fd_sc_hd__xor2_4 _17918_ (.A(_12731_),
    .B(_06502_),
    .X(_00878_));
 sky130_fd_sc_hd__nor2b_2 _17919_ (.A(net523),
    .B_N(\hash.CA2.f_dash[13] ),
    .Y(_12736_));
 sky130_fd_sc_hd__or2_1 _17920_ (.A(\hash.CA2.f_dash[11] ),
    .B(_06501_),
    .X(_06503_));
 sky130_fd_sc_hd__nand2_1 _17921_ (.A(\hash.CA2.f_dash[12] ),
    .B(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__xor2_4 _17922_ (.A(\hash.CA2.f_dash[13] ),
    .B(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__nor2_1 _17923_ (.A(net524),
    .B(_06505_),
    .Y(_00879_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1155 ();
 sky130_fd_sc_hd__nor2_1 _17925_ (.A(net523),
    .B(\hash.CA2.f_dash[14] ),
    .Y(_12741_));
 sky130_fd_sc_hd__and3_2 _17926_ (.A(\hash.CA2.f_dash[12] ),
    .B(\hash.CA2.f_dash[13] ),
    .C(_06502_),
    .X(_06507_));
 sky130_fd_sc_hd__xor2_4 _17927_ (.A(\hash.CA2.f_dash[14] ),
    .B(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__nor2_1 _17928_ (.A(net524),
    .B(_06508_),
    .Y(_00880_));
 sky130_fd_sc_hd__or2_2 _17929_ (.A(net523),
    .B(\hash.CA2.f_dash[15] ),
    .X(_06509_));
 sky130_fd_sc_hd__inv_1 _17930_ (.A(_06509_),
    .Y(_12746_));
 sky130_fd_sc_hd__a31o_4 _17931_ (.A1(\hash.CA2.f_dash[13] ),
    .A2(_12731_),
    .A3(_06503_),
    .B1(\hash.CA2.f_dash[14] ),
    .X(_06510_));
 sky130_fd_sc_hd__xor2_4 _17932_ (.A(\hash.CA2.f_dash[15] ),
    .B(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__nand2_1 _17933_ (.A(net519),
    .B(_06511_),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2b_4 _17934_ (.A(net523),
    .B_N(\hash.CA2.f_dash[16] ),
    .Y(_12751_));
 sky130_fd_sc_hd__nor3_1 _17935_ (.A(\hash.CA2.f_dash[14] ),
    .B(_06507_),
    .C(_06509_),
    .Y(_06512_));
 sky130_fd_sc_hd__xnor2_2 _17936_ (.A(_12751_),
    .B(_06512_),
    .Y(_00882_));
 sky130_fd_sc_hd__nor2b_4 _17937_ (.A(net523),
    .B_N(\hash.CA2.f_dash[17] ),
    .Y(_12756_));
 sky130_fd_sc_hd__o21ai_2 _17938_ (.A1(\hash.CA2.f_dash[15] ),
    .A2(_06510_),
    .B1(_12751_),
    .Y(_06513_));
 sky130_fd_sc_hd__xnor2_2 _17939_ (.A(_12756_),
    .B(_06513_),
    .Y(_00883_));
 sky130_fd_sc_hd__nor2b_4 _17940_ (.A(net523),
    .B_N(\hash.CA2.f_dash[18] ),
    .Y(_12761_));
 sky130_fd_sc_hd__o311a_2 _17941_ (.A1(\hash.CA2.f_dash[14] ),
    .A2(_06507_),
    .A3(_06509_),
    .B1(_12751_),
    .C1(\hash.CA2.f_dash[17] ),
    .X(_06514_));
 sky130_fd_sc_hd__xor2_2 _17942_ (.A(_12761_),
    .B(_06514_),
    .X(_00884_));
 sky130_fd_sc_hd__nor2b_4 _17943_ (.A(net522),
    .B_N(\hash.CA2.f_dash[19] ),
    .Y(_12766_));
 sky130_fd_sc_hd__o2111ai_4 _17944_ (.A1(_06509_),
    .A2(_06510_),
    .B1(_12751_),
    .C1(\hash.CA2.f_dash[18] ),
    .D1(\hash.CA2.f_dash[17] ),
    .Y(_06515_));
 sky130_fd_sc_hd__xnor2_4 _17945_ (.A(_12766_),
    .B(_06515_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _17946_ (.A(_06210_),
    .B(\hash.CA2.f_dash[20] ),
    .Y(_12965_));
 sky130_fd_sc_hd__inv_1 _17947_ (.A(_12965_),
    .Y(_12771_));
 sky130_fd_sc_hd__nand3_1 _17948_ (.A(\hash.CA2.f_dash[18] ),
    .B(\hash.CA2.f_dash[19] ),
    .C(_06514_),
    .Y(_06516_));
 sky130_fd_sc_hd__xor2_1 _17949_ (.A(\hash.CA2.f_dash[20] ),
    .B(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__nor2_1 _17950_ (.A(net522),
    .B(_06517_),
    .Y(_00886_));
 sky130_fd_sc_hd__nor2_1 _17951_ (.A(net522),
    .B(\hash.CA2.f_dash[21] ),
    .Y(_12776_));
 sky130_fd_sc_hd__clkinv_2 _17952_ (.A(_12776_),
    .Y(_12974_));
 sky130_fd_sc_hd__nand4_1 _17953_ (.A(\hash.CA2.f_dash[18] ),
    .B(\hash.CA2.f_dash[20] ),
    .C(_12756_),
    .D(_12766_),
    .Y(_06518_));
 sky130_fd_sc_hd__nor2_2 _17954_ (.A(_06513_),
    .B(_06518_),
    .Y(_06519_));
 sky130_fd_sc_hd__xnor2_2 _17955_ (.A(_12974_),
    .B(_06519_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_1 _17956_ (.A(net522),
    .B(\hash.CA2.f_dash[22] ),
    .Y(_12781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1154 ();
 sky130_fd_sc_hd__and4_1 _17958_ (.A(\hash.CA2.f_dash[19] ),
    .B(\hash.CA2.f_dash[20] ),
    .C(_12761_),
    .D(_06514_),
    .X(_06521_));
 sky130_fd_sc_hd__or3_1 _17959_ (.A(\hash.CA2.f_dash[21] ),
    .B(\hash.CA2.f_dash[22] ),
    .C(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__o21ai_0 _17960_ (.A1(\hash.CA2.f_dash[21] ),
    .A2(_06521_),
    .B1(\hash.CA2.f_dash[22] ),
    .Y(_06523_));
 sky130_fd_sc_hd__nand3_1 _17961_ (.A(_06210_),
    .B(_06522_),
    .C(_06523_),
    .Y(_00888_));
 sky130_fd_sc_hd__or2_1 _17962_ (.A(net522),
    .B(\hash.CA2.f_dash[23] ),
    .X(_12990_));
 sky130_fd_sc_hd__inv_1 _17963_ (.A(_12990_),
    .Y(_12786_));
 sky130_fd_sc_hd__nor3_1 _17964_ (.A(\hash.CA2.f_dash[21] ),
    .B(\hash.CA2.f_dash[22] ),
    .C(_06519_),
    .Y(_06524_));
 sky130_fd_sc_hd__xnor2_1 _17965_ (.A(\hash.CA2.f_dash[23] ),
    .B(_06524_),
    .Y(_06525_));
 sky130_fd_sc_hd__nand2_1 _17966_ (.A(net519),
    .B(_06525_),
    .Y(_00889_));
 sky130_fd_sc_hd__nor2_1 _17967_ (.A(net522),
    .B(\hash.CA2.f_dash[24] ),
    .Y(_12791_));
 sky130_fd_sc_hd__or3_1 _17968_ (.A(net522),
    .B(\hash.CA2.f_dash[21] ),
    .C(\hash.CA2.f_dash[22] ),
    .X(_06526_));
 sky130_fd_sc_hd__nor3_1 _17969_ (.A(\hash.CA2.f_dash[23] ),
    .B(_06521_),
    .C(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__xnor2_1 _17970_ (.A(\hash.CA2.f_dash[24] ),
    .B(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__nand2_1 _17971_ (.A(net519),
    .B(_06528_),
    .Y(_00890_));
 sky130_fd_sc_hd__nor2_1 _17972_ (.A(net522),
    .B(\hash.CA2.f_dash[25] ),
    .Y(_12796_));
 sky130_fd_sc_hd__inv_1 _17973_ (.A(_12796_),
    .Y(_13006_));
 sky130_fd_sc_hd__or3_1 _17974_ (.A(\hash.CA2.f_dash[24] ),
    .B(_12990_),
    .C(_06526_),
    .X(_06529_));
 sky130_fd_sc_hd__nor2_1 _17975_ (.A(_06519_),
    .B(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__xnor2_1 _17976_ (.A(_12796_),
    .B(_06530_),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2b_2 _17977_ (.A(net522),
    .B_N(\hash.CA2.f_dash[26] ),
    .Y(_12801_));
 sky130_fd_sc_hd__nor2_1 _17978_ (.A(_13006_),
    .B(_06529_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2b_1 _17979_ (.A_N(_06521_),
    .B(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__xor2_1 _17980_ (.A(_12801_),
    .B(_06532_),
    .X(_00892_));
 sky130_fd_sc_hd__nor2_1 _17981_ (.A(net522),
    .B(\hash.CA2.f_dash[27] ),
    .Y(_12806_));
 sky130_fd_sc_hd__inv_1 _17982_ (.A(_12806_),
    .Y(_13021_));
 sky130_fd_sc_hd__nand2b_1 _17983_ (.A_N(_06519_),
    .B(_06531_),
    .Y(_06533_));
 sky130_fd_sc_hd__nand2_1 _17984_ (.A(_12801_),
    .B(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__mux2_1 _17985_ (.A0(\hash.CA2.f_dash[27] ),
    .A1(_12806_),
    .S(_06534_),
    .X(_00893_));
 sky130_fd_sc_hd__or2_1 _17986_ (.A(net522),
    .B(\hash.CA2.f_dash[28] ),
    .X(_13029_));
 sky130_fd_sc_hd__inv_1 _17987_ (.A(_13029_),
    .Y(_12811_));
 sky130_fd_sc_hd__a21oi_1 _17988_ (.A1(\hash.CA2.f_dash[26] ),
    .A2(_06532_),
    .B1(\hash.CA2.f_dash[27] ),
    .Y(_06535_));
 sky130_fd_sc_hd__xnor2_1 _17989_ (.A(\hash.CA2.f_dash[28] ),
    .B(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_1 _17990_ (.A(net519),
    .B(_06536_),
    .Y(_00894_));
 sky130_fd_sc_hd__nor2b_2 _17991_ (.A(net522),
    .B_N(\hash.CA2.f_dash[29] ),
    .Y(_12816_));
 sky130_fd_sc_hd__nor2_1 _17992_ (.A(\hash.CA2.f_dash[27] ),
    .B(_13029_),
    .Y(_06537_));
 sky130_fd_sc_hd__and2_0 _17993_ (.A(_06534_),
    .B(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__xnor2_1 _17994_ (.A(_12816_),
    .B(_06538_),
    .Y(_00895_));
 sky130_fd_sc_hd__or2_1 _17995_ (.A(net522),
    .B(\hash.CA2.f_dash[30] ),
    .X(_13043_));
 sky130_fd_sc_hd__inv_1 _17996_ (.A(_13043_),
    .Y(_12821_));
 sky130_fd_sc_hd__inv_1 _17997_ (.A(_06535_),
    .Y(_06539_));
 sky130_fd_sc_hd__o21ai_1 _17998_ (.A1(\hash.CA2.f_dash[28] ),
    .A2(_06539_),
    .B1(\hash.CA2.f_dash[29] ),
    .Y(_06540_));
 sky130_fd_sc_hd__xnor2_1 _17999_ (.A(\hash.CA2.f_dash[30] ),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__nor2_1 _18000_ (.A(net522),
    .B(_06541_),
    .Y(_00897_));
 sky130_fd_sc_hd__o21ai_1 _18001_ (.A1(\hash.CA2.f_dash[27] ),
    .A2(\hash.CA2.f_dash[28] ),
    .B1(\hash.CA2.f_dash[29] ),
    .Y(_06542_));
 sky130_fd_sc_hd__a41oi_2 _18002_ (.A1(\hash.CA2.f_dash[26] ),
    .A2(\hash.CA2.f_dash[29] ),
    .A3(_06533_),
    .A4(_06537_),
    .B1(_13043_),
    .Y(_06543_));
 sky130_fd_sc_hd__nand3_1 _18003_ (.A(\hash.CA2.f_dash[31] ),
    .B(_06543_),
    .C(_06542_),
    .Y(_06544_));
 sky130_fd_sc_hd__o21a_1 _18004_ (.A1(\hash.CA2.f_dash[31] ),
    .A2(_06542_),
    .B1(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__nor2b_1 _18005_ (.A(net522),
    .B_N(\hash.CA2.f_dash[31] ),
    .Y(_06546_));
 sky130_fd_sc_hd__o22ai_1 _18006_ (.A1(net522),
    .A2(_06545_),
    .B1(_06546_),
    .B2(_06543_),
    .Y(_00898_));
 sky130_fd_sc_hd__xnor2_2 _18007_ (.A(_14017_),
    .B(_12546_),
    .Y(_00865_));
 sky130_fd_sc_hd__o21ai_0 _18008_ (.A1(\hash.CA2.e_dash[0] ),
    .A2(\hash.CA2.e_dash[1] ),
    .B1(\hash.CA2.e_dash[2] ),
    .Y(_06547_));
 sky130_fd_sc_hd__xnor2_1 _18009_ (.A(\hash.CA2.e_dash[3] ),
    .B(_06547_),
    .Y(_06548_));
 sky130_fd_sc_hd__nor2_2 _18010_ (.A(\hash.reset ),
    .B(_06548_),
    .Y(_00868_));
 sky130_fd_sc_hd__inv_1 _18011_ (.A(_14017_),
    .Y(_06549_));
 sky130_fd_sc_hd__a21oi_2 _18012_ (.A1(\hash.CA2.e_dash[2] ),
    .A2(_06549_),
    .B1(\hash.CA2.e_dash[3] ),
    .Y(_06550_));
 sky130_fd_sc_hd__xnor2_1 _18013_ (.A(_06482_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__nand2_2 _18014_ (.A(_06210_),
    .B(_06551_),
    .Y(_00869_));
 sky130_fd_sc_hd__o21a_1 _18015_ (.A1(\hash.CA2.e_dash[0] ),
    .A2(\hash.CA2.e_dash[1] ),
    .B1(_12546_),
    .X(_06552_));
 sky130_fd_sc_hd__o21ai_4 _18016_ (.A1(\hash.CA2.e_dash[3] ),
    .A2(_06552_),
    .B1(\hash.CA2.e_dash[4] ),
    .Y(_06553_));
 sky130_fd_sc_hd__xnor2_4 _18017_ (.A(\hash.CA2.e_dash[5] ),
    .B(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__nor2_1 _18018_ (.A(net520),
    .B(_06554_),
    .Y(_00870_));
 sky130_fd_sc_hd__o21ai_4 _18019_ (.A1(_06482_),
    .A2(_06550_),
    .B1(_12562_),
    .Y(_06555_));
 sky130_fd_sc_hd__xnor2_4 _18020_ (.A(_06483_),
    .B(_06555_),
    .Y(_00871_));
 sky130_fd_sc_hd__inv_1 _18021_ (.A(\hash.CA2.e_dash[5] ),
    .Y(_06556_));
 sky130_fd_sc_hd__a21boi_0 _18022_ (.A1(_06556_),
    .A2(_06553_),
    .B1_N(\hash.CA2.e_dash[6] ),
    .Y(_06557_));
 sky130_fd_sc_hd__xor2_1 _18023_ (.A(\hash.CA2.e_dash[7] ),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__nor2_1 _18024_ (.A(net520),
    .B(_06558_),
    .Y(_00872_));
 sky130_fd_sc_hd__a21oi_2 _18025_ (.A1(\hash.CA2.e_dash[6] ),
    .A2(_06555_),
    .B1(\hash.CA2.e_dash[7] ),
    .Y(_06559_));
 sky130_fd_sc_hd__xnor2_4 _18026_ (.A(\hash.CA2.e_dash[8] ),
    .B(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_1 _18027_ (.A(net519),
    .B(_06560_),
    .Y(_00873_));
 sky130_fd_sc_hd__a21oi_1 _18028_ (.A1(_06556_),
    .A2(_06553_),
    .B1(_06483_),
    .Y(_06561_));
 sky130_fd_sc_hd__or4_2 _18029_ (.A(\hash.reset ),
    .B(\hash.CA2.e_dash[7] ),
    .C(\hash.CA2.e_dash[8] ),
    .D(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__xor2_4 _18030_ (.A(_12578_),
    .B(_06562_),
    .X(_00874_));
 sky130_fd_sc_hd__a211oi_1 _18031_ (.A1(\hash.CA2.e_dash[6] ),
    .A2(_06555_),
    .B1(\hash.CA2.e_dash[8] ),
    .C1(\hash.CA2.e_dash[7] ),
    .Y(_06563_));
 sky130_fd_sc_hd__nand2b_1 _18032_ (.A_N(_06563_),
    .B(_12578_),
    .Y(_06564_));
 sky130_fd_sc_hd__xnor2_2 _18033_ (.A(_12581_),
    .B(_06564_),
    .Y(_00844_));
 sky130_fd_sc_hd__and3_2 _18034_ (.A(\hash.CA2.e_dash[10] ),
    .B(_12578_),
    .C(_06562_),
    .X(_06565_));
 sky130_fd_sc_hd__xor2_4 _18035_ (.A(_12586_),
    .B(_06565_),
    .X(_00845_));
 sky130_fd_sc_hd__a2111oi_1 _18036_ (.A1(\hash.CA2.e_dash[6] ),
    .A2(_06555_),
    .B1(\hash.CA2.e_dash[7] ),
    .C1(\hash.reset ),
    .D1(\hash.CA2.e_dash[8] ),
    .Y(_06566_));
 sky130_fd_sc_hd__nand2_1 _18037_ (.A(\hash.CA2.e_dash[9] ),
    .B(\hash.CA2.e_dash[10] ),
    .Y(_06567_));
 sky130_fd_sc_hd__o21ai_0 _18038_ (.A1(_06566_),
    .A2(_06567_),
    .B1(_12586_),
    .Y(_06568_));
 sky130_fd_sc_hd__xor2_1 _18039_ (.A(_12591_),
    .B(_06568_),
    .X(_00846_));
 sky130_fd_sc_hd__nor4_4 _18040_ (.A(net523),
    .B(\hash.CA2.e_dash[11] ),
    .C(\hash.CA2.e_dash[12] ),
    .D(_06565_),
    .Y(_06569_));
 sky130_fd_sc_hd__xnor2_4 _18041_ (.A(_12594_),
    .B(_06569_),
    .Y(_00847_));
 sky130_fd_sc_hd__and3b_1 _18042_ (.A_N(_06563_),
    .B(_12581_),
    .C(_12578_),
    .X(_06570_));
 sky130_fd_sc_hd__o311a_2 _18043_ (.A1(\hash.CA2.e_dash[11] ),
    .A2(\hash.CA2.e_dash[12] ),
    .A3(_06570_),
    .B1(\hash.CA2.e_dash[13] ),
    .C1(_06210_),
    .X(_06571_));
 sky130_fd_sc_hd__xor2_4 _18044_ (.A(_12599_),
    .B(_06571_),
    .X(_00848_));
 sky130_fd_sc_hd__o31ai_1 _18045_ (.A1(\hash.CA2.e_dash[11] ),
    .A2(\hash.CA2.e_dash[12] ),
    .A3(_06565_),
    .B1(\hash.CA2.e_dash[13] ),
    .Y(_06572_));
 sky130_fd_sc_hd__nand2_1 _18046_ (.A(_12599_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__xor2_4 _18047_ (.A(_12604_),
    .B(_06573_),
    .X(_00849_));
 sky130_fd_sc_hd__nor4_2 _18048_ (.A(net523),
    .B(\hash.CA2.e_dash[14] ),
    .C(\hash.CA2.e_dash[15] ),
    .D(_06571_),
    .Y(_06574_));
 sky130_fd_sc_hd__xnor2_2 _18049_ (.A(_12609_),
    .B(_06574_),
    .Y(_00850_));
 sky130_fd_sc_hd__inv_1 _18050_ (.A(_06569_),
    .Y(_06575_));
 sky130_fd_sc_hd__or4_2 _18051_ (.A(net523),
    .B(\hash.CA2.e_dash[14] ),
    .C(\hash.CA2.e_dash[15] ),
    .D(\hash.CA2.e_dash[16] ),
    .X(_06576_));
 sky130_fd_sc_hd__a21oi_4 _18052_ (.A1(\hash.CA2.e_dash[13] ),
    .A2(_06575_),
    .B1(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__xnor2_2 _18053_ (.A(_12614_),
    .B(_06577_),
    .Y(_00851_));
 sky130_fd_sc_hd__clkinvlp_4 _18054_ (.A(_12617_),
    .Y(_06578_));
 sky130_fd_sc_hd__or3_4 _18055_ (.A(\hash.CA2.e_dash[17] ),
    .B(_06571_),
    .C(_06576_),
    .X(_06579_));
 sky130_fd_sc_hd__xnor2_2 _18056_ (.A(_06578_),
    .B(_06579_),
    .Y(_00852_));
 sky130_fd_sc_hd__a21oi_1 _18057_ (.A1(_12614_),
    .A2(_06577_),
    .B1(_06578_),
    .Y(_06580_));
 sky130_fd_sc_hd__mux2i_1 _18058_ (.A0(_06485_),
    .A1(\hash.CA2.e_dash[19] ),
    .S(_06580_),
    .Y(_00853_));
 sky130_fd_sc_hd__and3_1 _18059_ (.A(\hash.CA2.e_dash[19] ),
    .B(_12617_),
    .C(_06579_),
    .X(_06581_));
 sky130_fd_sc_hd__xor2_2 _18060_ (.A(_12623_),
    .B(_06581_),
    .X(_00855_));
 sky130_fd_sc_hd__nand3_1 _18061_ (.A(\hash.CA2.e_dash[19] ),
    .B(\hash.CA2.e_dash[20] ),
    .C(_06580_),
    .Y(_06582_));
 sky130_fd_sc_hd__xnor2_1 _18062_ (.A(_12626_),
    .B(_06582_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand3_1 _18063_ (.A(\hash.CA2.e_dash[20] ),
    .B(\hash.CA2.e_dash[21] ),
    .C(_06581_),
    .Y(_06583_));
 sky130_fd_sc_hd__xor2_1 _18064_ (.A(\hash.CA2.e_dash[22] ),
    .B(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__nor2_1 _18065_ (.A(net522),
    .B(_06584_),
    .Y(_00857_));
 sky130_fd_sc_hd__nand3_1 _18066_ (.A(\hash.CA2.e_dash[20] ),
    .B(\hash.CA2.e_dash[22] ),
    .C(_12626_),
    .Y(_06585_));
 sky130_fd_sc_hd__a2111oi_4 _18067_ (.A1(_12614_),
    .A2(_06577_),
    .B1(_06585_),
    .C1(_06578_),
    .D1(_06485_),
    .Y(_06586_));
 sky130_fd_sc_hd__xnor2_1 _18068_ (.A(_06486_),
    .B(_06586_),
    .Y(_00858_));
 sky130_fd_sc_hd__nand4_2 _18069_ (.A(\hash.CA2.e_dash[20] ),
    .B(\hash.CA2.e_dash[22] ),
    .C(_12626_),
    .D(_06581_),
    .Y(_06587_));
 sky130_fd_sc_hd__nor2b_1 _18070_ (.A(\hash.CA2.e_dash[23] ),
    .B_N(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__xnor2_1 _18071_ (.A(\hash.CA2.e_dash[24] ),
    .B(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__nand2_1 _18072_ (.A(_06210_),
    .B(_06589_),
    .Y(_00859_));
 sky130_fd_sc_hd__nor3_1 _18073_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .C(_06586_),
    .Y(_06590_));
 sky130_fd_sc_hd__xnor2_1 _18074_ (.A(\hash.CA2.e_dash[25] ),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__nand2_1 _18075_ (.A(_06210_),
    .B(_06591_),
    .Y(_00860_));
 sky130_fd_sc_hd__or4_1 _18076_ (.A(net522),
    .B(\hash.CA2.e_dash[23] ),
    .C(\hash.CA2.e_dash[24] ),
    .D(\hash.CA2.e_dash[25] ),
    .X(_06592_));
 sky130_fd_sc_hd__nor2b_1 _18077_ (.A(_06592_),
    .B_N(_06587_),
    .Y(_06593_));
 sky130_fd_sc_hd__xnor2_1 _18078_ (.A(_12649_),
    .B(_06593_),
    .Y(_00861_));
 sky130_fd_sc_hd__nor3_1 _18079_ (.A(\hash.CA2.e_dash[26] ),
    .B(_06586_),
    .C(_06592_),
    .Y(_06594_));
 sky130_fd_sc_hd__xnor2_1 _18080_ (.A(_12654_),
    .B(_06594_),
    .Y(_00862_));
 sky130_fd_sc_hd__nor2_1 _18081_ (.A(\hash.CA2.e_dash[26] ),
    .B(_06592_),
    .Y(_06595_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(_12654_),
    .B(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__o21bai_1 _18083_ (.A1(_06486_),
    .A2(_06587_),
    .B1_N(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__xor2_1 _18084_ (.A(_12659_),
    .B(_06597_),
    .X(_00863_));
 sky130_fd_sc_hd__nor3_1 _18085_ (.A(\hash.CA2.e_dash[28] ),
    .B(_06586_),
    .C(_06596_),
    .Y(_06598_));
 sky130_fd_sc_hd__xnor2_1 _18086_ (.A(_12662_),
    .B(_06598_),
    .Y(_00864_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1153 ();
 sky130_fd_sc_hd__o21ai_0 _18088_ (.A1(\hash.CA2.e_dash[28] ),
    .A2(_06597_),
    .B1(\hash.CA2.e_dash[29] ),
    .Y(_06600_));
 sky130_fd_sc_hd__xor2_1 _18089_ (.A(\hash.CA2.e_dash[30] ),
    .B(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__nor2_1 _18090_ (.A(net522),
    .B(_06601_),
    .Y(_00866_));
 sky130_fd_sc_hd__nor2b_4 _18091_ (.A(net522),
    .B_N(\hash.CA2.e_dash[31] ),
    .Y(_06602_));
 sky130_fd_sc_hd__nand3b_1 _18092_ (.A_N(_06598_),
    .B(_12662_),
    .C(\hash.CA2.e_dash[30] ),
    .Y(_06603_));
 sky130_fd_sc_hd__xnor2_1 _18093_ (.A(_06602_),
    .B(_06603_),
    .Y(_00867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1152 ();
 sky130_fd_sc_hd__nor2b_2 _18095_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[4] ),
    .Y(\hash.CA1.f[4] ));
 sky130_fd_sc_hd__xnor2_2 _18096_ (.A(_14020_),
    .B(\hash.CA1.f[4] ),
    .Y(_00835_));
 sky130_fd_sc_hd__nor2b_1 _18097_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[5] ),
    .Y(\hash.CA1.f[5] ));
 sky130_fd_sc_hd__o21ai_2 _18098_ (.A1(\hash.CA2.S1.X[2] ),
    .A2(\hash.CA2.S1.X[3] ),
    .B1(\hash.CA2.S1.X[4] ),
    .Y(_06605_));
 sky130_fd_sc_hd__xor2_4 _18099_ (.A(\hash.CA2.S1.X[5] ),
    .B(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__nor2_1 _18100_ (.A(net520),
    .B(_06606_),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2b_1 _18101_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[6] ),
    .Y(\hash.CA1.f[6] ));
 sky130_fd_sc_hd__inv_1 _18102_ (.A(net1091),
    .Y(_06607_));
 sky130_fd_sc_hd__nand3b_2 _18103_ (.A_N(_14020_),
    .B(\hash.CA2.S1.X[5] ),
    .C(\hash.CA2.S1.X[4] ),
    .Y(_06608_));
 sky130_fd_sc_hd__xnor2_2 _18104_ (.A(_06607_),
    .B(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__nor2_1 _18105_ (.A(net520),
    .B(_06609_),
    .Y(_00837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1151 ();
 sky130_fd_sc_hd__inv_1 _18107_ (.A(\hash.CA2.S1.X[7] ),
    .Y(_06611_));
 sky130_fd_sc_hd__nand2_1 _18108_ (.A(_06210_),
    .B(_06611_),
    .Y(\hash.CA1.f[7] ));
 sky130_fd_sc_hd__o211a_1 _18109_ (.A1(\hash.CA2.S1.X[2] ),
    .A2(\hash.CA2.S1.X[3] ),
    .B1(\hash.CA2.S1.X[4] ),
    .C1(\hash.CA2.S1.X[5] ),
    .X(_06612_));
 sky130_fd_sc_hd__and3_1 _18110_ (.A(_06611_),
    .B(net1092),
    .C(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__a21oi_1 _18111_ (.A1(net1093),
    .A2(_06612_),
    .B1(_06611_),
    .Y(_06614_));
 sky130_fd_sc_hd__nor3_2 _18112_ (.A(\hash.reset ),
    .B(_06613_),
    .C(_06614_),
    .Y(_00838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1150 ();
 sky130_fd_sc_hd__nor2b_1 _18114_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[8] ),
    .Y(\hash.CA1.f[8] ));
 sky130_fd_sc_hd__o31a_2 _18115_ (.A1(\hash.reset ),
    .A2(_06607_),
    .A3(_06608_),
    .B1(_06611_),
    .X(_06616_));
 sky130_fd_sc_hd__xor2_4 _18116_ (.A(\hash.CA2.S1.X[8] ),
    .B(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__nand2_1 _18117_ (.A(net519),
    .B(_06617_),
    .Y(_00839_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1149 ();
 sky130_fd_sc_hd__nor2b_1 _18119_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[9] ),
    .Y(\hash.CA1.f[9] ));
 sky130_fd_sc_hd__nand2_1 _18120_ (.A(\hash.CA1.f[6] ),
    .B(_06612_),
    .Y(_06619_));
 sky130_fd_sc_hd__nand2_1 _18121_ (.A(_06611_),
    .B(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__nand2_1 _18122_ (.A(\hash.CA2.S1.X[8] ),
    .B(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__xor2_1 _18123_ (.A(\hash.CA2.S1.X[9] ),
    .B(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__nor2_2 _18124_ (.A(\hash.reset ),
    .B(_06622_),
    .Y(_00840_));
 sky130_fd_sc_hd__nand2_1 _18125_ (.A(_06210_),
    .B(\hash.CA2.S1.X[10] ),
    .Y(_06623_));
 sky130_fd_sc_hd__inv_1 _18126_ (.A(_06623_),
    .Y(\hash.CA1.f[10] ));
 sky130_fd_sc_hd__nand2_1 _18127_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA1.f[9] ),
    .Y(_06624_));
 sky130_fd_sc_hd__nor2_1 _18128_ (.A(_06616_),
    .B(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__xnor2_1 _18129_ (.A(_06623_),
    .B(_06625_),
    .Y(_00841_));
 sky130_fd_sc_hd__nor2_1 _18130_ (.A(\hash.reset ),
    .B(\hash.CA2.S1.X[11] ),
    .Y(_06626_));
 sky130_fd_sc_hd__inv_1 _18131_ (.A(_06626_),
    .Y(\hash.CA1.f[11] ));
 sky130_fd_sc_hd__and4_2 _18132_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[10] ),
    .C(\hash.CA1.f[9] ),
    .D(_06620_),
    .X(_06627_));
 sky130_fd_sc_hd__xnor2_4 _18133_ (.A(\hash.CA1.f[11] ),
    .B(_06627_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2b_2 _18134_ (.A(net523),
    .B_N(\hash.CA2.S1.X[12] ),
    .Y(\hash.CA1.f[12] ));
 sky130_fd_sc_hd__o31ai_2 _18135_ (.A1(_06616_),
    .A2(_06623_),
    .A3(_06624_),
    .B1(_06626_),
    .Y(_06628_));
 sky130_fd_sc_hd__nor2_1 _18136_ (.A(\hash.CA2.S1.X[12] ),
    .B(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__a21oi_1 _18137_ (.A1(\hash.CA1.f[12] ),
    .A2(_06628_),
    .B1(_06629_),
    .Y(_00814_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1148 ();
 sky130_fd_sc_hd__inv_1 _18139_ (.A(\hash.CA2.S1.X[13] ),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_1 _18140_ (.A(_06210_),
    .B(_06631_),
    .Y(\hash.CA1.f[13] ));
 sky130_fd_sc_hd__o21ai_4 _18141_ (.A1(\hash.CA2.S1.X[11] ),
    .A2(_06627_),
    .B1(\hash.CA1.f[12] ),
    .Y(_06632_));
 sky130_fd_sc_hd__mux2i_4 _18142_ (.A0(_06631_),
    .A1(\hash.CA1.f[13] ),
    .S(_06632_),
    .Y(_00815_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1147 ();
 sky130_fd_sc_hd__or2_0 _18144_ (.A(net523),
    .B(\hash.CA2.S1.X[14] ),
    .X(\hash.CA1.f[14] ));
 sky130_fd_sc_hd__a21o_1 _18145_ (.A1(\hash.CA1.f[10] ),
    .A2(_06625_),
    .B1(\hash.CA2.S1.X[11] ),
    .X(_06634_));
 sky130_fd_sc_hd__a21oi_1 _18146_ (.A1(\hash.CA2.S1.X[12] ),
    .A2(_06634_),
    .B1(\hash.CA2.S1.X[13] ),
    .Y(_06635_));
 sky130_fd_sc_hd__xnor2_1 _18147_ (.A(\hash.CA2.S1.X[14] ),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__nand2_1 _18148_ (.A(_06210_),
    .B(_06636_),
    .Y(_00816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1146 ();
 sky130_fd_sc_hd__nand2_2 _18150_ (.A(_06210_),
    .B(\hash.CA2.S1.X[15] ),
    .Y(_06638_));
 sky130_fd_sc_hd__inv_1 _18151_ (.A(_06638_),
    .Y(\hash.CA1.f[15] ));
 sky130_fd_sc_hd__nor2_2 _18152_ (.A(\hash.CA2.S1.X[14] ),
    .B(\hash.CA1.f[13] ),
    .Y(_06639_));
 sky130_fd_sc_hd__a21oi_2 _18153_ (.A1(_06632_),
    .A2(_06639_),
    .B1(_06638_),
    .Y(_06640_));
 sky130_fd_sc_hd__and3_1 _18154_ (.A(_06632_),
    .B(_06638_),
    .C(_06639_),
    .X(_06641_));
 sky130_fd_sc_hd__nor2_2 _18155_ (.A(_06640_),
    .B(_06641_),
    .Y(_00817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1145 ();
 sky130_fd_sc_hd__inv_1 _18157_ (.A(\hash.CA2.S1.X[16] ),
    .Y(_06643_));
 sky130_fd_sc_hd__nand2_2 _18158_ (.A(_06210_),
    .B(_06643_),
    .Y(\hash.CA1.f[16] ));
 sky130_fd_sc_hd__nand2_1 _18159_ (.A(\hash.CA2.S1.X[12] ),
    .B(_06628_),
    .Y(_06644_));
 sky130_fd_sc_hd__a21oi_4 _18160_ (.A1(_06639_),
    .A2(_06644_),
    .B1(_06638_),
    .Y(_06645_));
 sky130_fd_sc_hd__xnor2_4 _18161_ (.A(\hash.CA1.f[16] ),
    .B(_06645_),
    .Y(_00818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1144 ();
 sky130_fd_sc_hd__nor2b_2 _18163_ (.A(net523),
    .B_N(\hash.CA2.S1.X[17] ),
    .Y(\hash.CA1.f[17] ));
 sky130_fd_sc_hd__nor2_2 _18164_ (.A(_06640_),
    .B(\hash.CA1.f[16] ),
    .Y(_06647_));
 sky130_fd_sc_hd__xnor2_4 _18165_ (.A(\hash.CA1.f[17] ),
    .B(_06647_),
    .Y(_00819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1143 ();
 sky130_fd_sc_hd__nor2_2 _18167_ (.A(net522),
    .B(\hash.CA2.S1.X[18] ),
    .Y(_06649_));
 sky130_fd_sc_hd__inv_1 _18168_ (.A(_06649_),
    .Y(\hash.CA1.f[18] ));
 sky130_fd_sc_hd__inv_1 _18169_ (.A(\hash.CA2.S1.X[18] ),
    .Y(_06650_));
 sky130_fd_sc_hd__o21ai_2 _18170_ (.A1(\hash.CA2.S1.X[16] ),
    .A2(_06645_),
    .B1(\hash.CA1.f[17] ),
    .Y(_06651_));
 sky130_fd_sc_hd__nand2_2 _18171_ (.A(_06649_),
    .B(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__o21ai_2 _18172_ (.A1(_06650_),
    .A2(_06651_),
    .B1(_06652_),
    .Y(_00820_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1142 ();
 sky130_fd_sc_hd__nor2b_2 _18174_ (.A(net522),
    .B_N(\hash.CA2.S1.X[19] ),
    .Y(\hash.CA1.f[19] ));
 sky130_fd_sc_hd__o21ai_1 _18175_ (.A1(\hash.CA2.S1.X[16] ),
    .A2(_06640_),
    .B1(\hash.CA2.S1.X[17] ),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_2 _18176_ (.A(_06649_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__xor2_1 _18177_ (.A(\hash.CA1.f[19] ),
    .B(_06655_),
    .X(_00821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1141 ();
 sky130_fd_sc_hd__nor2b_1 _18179_ (.A(net522),
    .B_N(\hash.CA2.S1.X[20] ),
    .Y(\hash.CA1.f[20] ));
 sky130_fd_sc_hd__nand2_1 _18180_ (.A(\hash.CA2.S1.X[19] ),
    .B(_06652_),
    .Y(_06657_));
 sky130_fd_sc_hd__xor2_2 _18181_ (.A(\hash.CA2.S1.X[20] ),
    .B(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__nor2_1 _18182_ (.A(net522),
    .B(_06658_),
    .Y(_00822_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1140 ();
 sky130_fd_sc_hd__nor2b_1 _18184_ (.A(net522),
    .B_N(\hash.CA2.S1.X[21] ),
    .Y(\hash.CA1.f[21] ));
 sky130_fd_sc_hd__nand3_1 _18185_ (.A(\hash.CA2.S1.X[20] ),
    .B(\hash.CA1.f[19] ),
    .C(_06655_),
    .Y(_06660_));
 sky130_fd_sc_hd__xnor2_1 _18186_ (.A(\hash.CA1.f[21] ),
    .B(_06660_),
    .Y(_00823_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1139 ();
 sky130_fd_sc_hd__nand2_1 _18188_ (.A(_06210_),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_06662_));
 sky130_fd_sc_hd__inv_1 _18189_ (.A(_06662_),
    .Y(\hash.CA1.f[22] ));
 sky130_fd_sc_hd__nand3_1 _18190_ (.A(\hash.CA2.S1.X[20] ),
    .B(\hash.CA2.S1.X[21] ),
    .C(\hash.CA1.f[19] ),
    .Y(_06663_));
 sky130_fd_sc_hd__a21oi_1 _18191_ (.A1(_06650_),
    .A2(_06651_),
    .B1(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__xnor2_1 _18192_ (.A(_06662_),
    .B(_06664_),
    .Y(_00825_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1138 ();
 sky130_fd_sc_hd__nor2b_1 _18194_ (.A(net522),
    .B_N(\hash.CA2.S1.X[23] ),
    .Y(\hash.CA1.f[23] ));
 sky130_fd_sc_hd__nor2_2 _18195_ (.A(_06662_),
    .B(_06663_),
    .Y(_06666_));
 sky130_fd_sc_hd__nand2_1 _18196_ (.A(_06655_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__xnor2_1 _18197_ (.A(\hash.CA1.f[23] ),
    .B(_06667_),
    .Y(_00826_));
 sky130_fd_sc_hd__or2_1 _18198_ (.A(net522),
    .B(\hash.CA2.S1.X[24] ),
    .X(_06668_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1137 ();
 sky130_fd_sc_hd__nand3_1 _18200_ (.A(\hash.CA2.S1.X[23] ),
    .B(_06652_),
    .C(_06666_),
    .Y(_06669_));
 sky130_fd_sc_hd__xor2_2 _18201_ (.A(_06668_),
    .B(_06669_),
    .X(_00827_));
 sky130_fd_sc_hd__inv_1 _18202_ (.A(net1032),
    .Y(_06670_));
 sky130_fd_sc_hd__nand2_1 _18203_ (.A(_06210_),
    .B(_06670_),
    .Y(\hash.CA1.f[25] ));
 sky130_fd_sc_hd__a31oi_4 _18204_ (.A1(\hash.CA2.S1.X[23] ),
    .A2(_06655_),
    .A3(_06666_),
    .B1(\hash.CA2.S1.X[24] ),
    .Y(_06671_));
 sky130_fd_sc_hd__xnor2_2 _18205_ (.A(net1022),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_1 _18206_ (.A(net519),
    .B(_06672_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_2 _18207_ (.A(_06210_),
    .B(\hash.CA2.S1.X[26] ),
    .Y(_06673_));
 sky130_fd_sc_hd__inv_1 _18208_ (.A(_06673_),
    .Y(\hash.CA1.f[26] ));
 sky130_fd_sc_hd__a311o_2 _18209_ (.A1(\hash.CA2.S1.X[23] ),
    .A2(_06652_),
    .A3(_06666_),
    .B1(_06668_),
    .C1(net1031),
    .X(_06674_));
 sky130_fd_sc_hd__xnor2_1 _18210_ (.A(_06673_),
    .B(_06674_),
    .Y(_00829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1136 ();
 sky130_fd_sc_hd__or2_0 _18212_ (.A(net522),
    .B(net1152),
    .X(\hash.CA1.f[27] ));
 sky130_fd_sc_hd__a21oi_2 _18213_ (.A1(_06670_),
    .A2(_06671_),
    .B1(_06673_),
    .Y(_06676_));
 sky130_fd_sc_hd__xnor2_1 _18214_ (.A(\hash.CA1.f[27] ),
    .B(_06676_),
    .Y(_00830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1135 ();
 sky130_fd_sc_hd__or2_1 _18216_ (.A(net522),
    .B(\hash.CA2.S1.X[28] ),
    .X(\hash.CA1.f[28] ));
 sky130_fd_sc_hd__a21oi_1 _18217_ (.A1(\hash.CA2.S1.X[26] ),
    .A2(_06674_),
    .B1(net1150),
    .Y(_06678_));
 sky130_fd_sc_hd__xnor2_1 _18218_ (.A(\hash.CA2.S1.X[28] ),
    .B(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__nand2_1 _18219_ (.A(_06210_),
    .B(_06679_),
    .Y(_00831_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1134 ();
 sky130_fd_sc_hd__nor2b_1 _18221_ (.A(net522),
    .B_N(\hash.CA2.S1.X[29] ),
    .Y(\hash.CA1.f[29] ));
 sky130_fd_sc_hd__or3_1 _18222_ (.A(net1151),
    .B(_06676_),
    .C(\hash.CA1.f[28] ),
    .X(_06681_));
 sky130_fd_sc_hd__xor2_1 _18223_ (.A(\hash.CA1.f[29] ),
    .B(_06681_),
    .X(_00832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1133 ();
 sky130_fd_sc_hd__nor2b_1 _18225_ (.A(net522),
    .B_N(\hash.CA2.S1.X[30] ),
    .Y(\hash.CA1.f[30] ));
 sky130_fd_sc_hd__inv_1 _18226_ (.A(_06678_),
    .Y(_06683_));
 sky130_fd_sc_hd__o21ai_0 _18227_ (.A1(\hash.CA2.S1.X[28] ),
    .A2(_06683_),
    .B1(\hash.CA2.S1.X[29] ),
    .Y(_06684_));
 sky130_fd_sc_hd__xor2_1 _18228_ (.A(\hash.CA2.S1.X[30] ),
    .B(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__nor2_1 _18229_ (.A(net522),
    .B(_06685_),
    .Y(_00833_));
 sky130_fd_sc_hd__or2_1 _18230_ (.A(net522),
    .B(\hash.CA2.S1.X[31] ),
    .X(\hash.CA1.f[31] ));
 sky130_fd_sc_hd__nand3_1 _18231_ (.A(\hash.CA2.S1.X[29] ),
    .B(_06681_),
    .C(\hash.CA1.f[30] ),
    .Y(_06686_));
 sky130_fd_sc_hd__xor2_1 _18232_ (.A(\hash.CA1.f[31] ),
    .B(_06686_),
    .X(_00834_));
 sky130_fd_sc_hd__xnor2_2 _18233_ (.A(_12535_),
    .B(_13617_),
    .Y(_06687_));
 sky130_fd_sc_hd__and2_4 _18234_ (.A(_06210_),
    .B(_06687_),
    .X(_06688_));
 sky130_fd_sc_hd__inv_2 _18235_ (.A(_06688_),
    .Y(\hash.CA1.S1.X[2] ));
 sky130_fd_sc_hd__xnor2_2 _18236_ (.A(_14023_),
    .B(_06688_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand2_4 _18237_ (.A(_06210_),
    .B(_12536_),
    .Y(\hash.CA1.S1.X[1] ));
 sky130_fd_sc_hd__inv_1 _18238_ (.A(_00781_),
    .Y(\hash.CA1.S1.X[0] ));
 sky130_fd_sc_hd__a21o_1 _18239_ (.A1(_12534_),
    .A2(_13615_),
    .B1(_13614_),
    .X(_06689_));
 sky130_fd_sc_hd__a21oi_2 _18240_ (.A1(_13617_),
    .A2(_06689_),
    .B1(_13616_),
    .Y(_06690_));
 sky130_fd_sc_hd__xnor2_4 _18241_ (.A(_13619_),
    .B(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__nor2_8 _18242_ (.A(\hash.reset ),
    .B(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__clkinv_4 _18243_ (.A(_06692_),
    .Y(\hash.CA1.S1.X[3] ));
 sky130_fd_sc_hd__and3_1 _18244_ (.A(_12536_),
    .B(_00781_),
    .C(_06687_),
    .X(_06693_));
 sky130_fd_sc_hd__xnor2_2 _18245_ (.A(_06692_),
    .B(_06693_),
    .Y(_00806_));
 sky130_fd_sc_hd__clkinv_2 _18246_ (.A(_13621_),
    .Y(_06694_));
 sky130_fd_sc_hd__inv_1 _18247_ (.A(_13619_),
    .Y(_06695_));
 sky130_fd_sc_hd__a21oi_2 _18248_ (.A1(_12535_),
    .A2(_13617_),
    .B1(_13616_),
    .Y(_06696_));
 sky130_fd_sc_hd__o21bai_2 _18249_ (.A1(_06695_),
    .A2(_06696_),
    .B1_N(_13618_),
    .Y(_06697_));
 sky130_fd_sc_hd__xnor2_4 _18250_ (.A(_06694_),
    .B(_06697_),
    .Y(_06698_));
 sky130_fd_sc_hd__nor2_8 _18251_ (.A(\hash.reset ),
    .B(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__inv_1 _18252_ (.A(_06699_),
    .Y(\hash.CA1.S1.X[4] ));
 sky130_fd_sc_hd__and3_2 _18253_ (.A(_06210_),
    .B(_14023_),
    .C(_06687_),
    .X(_06700_));
 sky130_fd_sc_hd__nand2_1 _18254_ (.A(_06692_),
    .B(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__xnor2_2 _18255_ (.A(\hash.CA1.S1.X[4] ),
    .B(_06701_),
    .Y(_00807_));
 sky130_fd_sc_hd__a211oi_4 _18256_ (.A1(_12534_),
    .A2(_13615_),
    .B1(_13614_),
    .C1(_13616_),
    .Y(_06702_));
 sky130_fd_sc_hd__o211ai_4 _18257_ (.A1(_13617_),
    .A2(_13616_),
    .B1(_13621_),
    .C1(_13619_),
    .Y(_06703_));
 sky130_fd_sc_hd__a21oi_4 _18258_ (.A1(_13621_),
    .A2(_13618_),
    .B1(_13620_),
    .Y(_06704_));
 sky130_fd_sc_hd__o21ai_2 _18259_ (.A1(_06702_),
    .A2(_06703_),
    .B1(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__xor2_4 _18260_ (.A(_13623_),
    .B(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__nor2_8 _18261_ (.A(\hash.reset ),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__inv_1 _18262_ (.A(_06707_),
    .Y(\hash.CA1.S1.X[5] ));
 sky130_fd_sc_hd__nand3b_1 _18263_ (.A_N(_06698_),
    .B(_06693_),
    .C(_06692_),
    .Y(_06708_));
 sky130_fd_sc_hd__xnor2_2 _18264_ (.A(\hash.CA1.S1.X[5] ),
    .B(_06708_),
    .Y(_00808_));
 sky130_fd_sc_hd__nor2b_1 _18265_ (.A(\hash.reset ),
    .B_N(_13625_),
    .Y(_06709_));
 sky130_fd_sc_hd__nor2_1 _18266_ (.A(\hash.reset ),
    .B(_13625_),
    .Y(_06710_));
 sky130_fd_sc_hd__o31ai_1 _18267_ (.A1(_06695_),
    .A2(_06694_),
    .A3(_06696_),
    .B1(_06704_),
    .Y(_06711_));
 sky130_fd_sc_hd__a21oi_1 _18268_ (.A1(_13623_),
    .A2(_06711_),
    .B1(_13622_),
    .Y(_06712_));
 sky130_fd_sc_hd__mux2_8 _18269_ (.A0(_06709_),
    .A1(_06710_),
    .S(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__clkinv_4 _18270_ (.A(_06713_),
    .Y(\hash.CA1.S1.X[6] ));
 sky130_fd_sc_hd__nor4_4 _18271_ (.A(\hash.reset ),
    .B(_06691_),
    .C(_06698_),
    .D(_06706_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand2_1 _18272_ (.A(_06700_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__xnor2_2 _18273_ (.A(\hash.CA1.S1.X[6] ),
    .B(_06715_),
    .Y(_00809_));
 sky130_fd_sc_hd__o21a_1 _18274_ (.A1(_13623_),
    .A2(_13622_),
    .B1(_13625_),
    .X(_06716_));
 sky130_fd_sc_hd__nor2_1 _18275_ (.A(_13624_),
    .B(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__nor2_1 _18276_ (.A(_13622_),
    .B(_13624_),
    .Y(_06718_));
 sky130_fd_sc_hd__o211a_1 _18277_ (.A1(_06702_),
    .A2(_06703_),
    .B1(_06704_),
    .C1(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__o21a_1 _18278_ (.A1(_06717_),
    .A2(_06719_),
    .B1(_13627_),
    .X(_06720_));
 sky130_fd_sc_hd__nor3_1 _18279_ (.A(_13627_),
    .B(_06717_),
    .C(_06719_),
    .Y(_06721_));
 sky130_fd_sc_hd__o21ai_4 _18280_ (.A1(_06720_),
    .A2(_06721_),
    .B1(_06210_),
    .Y(_06722_));
 sky130_fd_sc_hd__clkinv_4 _18281_ (.A(_06722_),
    .Y(\hash.CA1.S1.X[7] ));
 sky130_fd_sc_hd__nand3_2 _18282_ (.A(_06693_),
    .B(_06713_),
    .C(_06714_),
    .Y(_06723_));
 sky130_fd_sc_hd__xnor2_2 _18283_ (.A(_06722_),
    .B(_06723_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor3_1 _18284_ (.A(_13623_),
    .B(_13622_),
    .C(_13624_),
    .Y(_06724_));
 sky130_fd_sc_hd__o21ai_1 _18285_ (.A1(_13625_),
    .A2(_13624_),
    .B1(_13627_),
    .Y(_06725_));
 sky130_fd_sc_hd__o21bai_2 _18286_ (.A1(_06724_),
    .A2(_06725_),
    .B1_N(_13626_),
    .Y(_06726_));
 sky130_fd_sc_hd__nor3_1 _18287_ (.A(_13622_),
    .B(_13624_),
    .C(_13626_),
    .Y(_06727_));
 sky130_fd_sc_hd__o311ai_4 _18288_ (.A1(_06695_),
    .A2(_06694_),
    .A3(_06696_),
    .B1(_06704_),
    .C1(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__a21oi_1 _18289_ (.A1(_06726_),
    .A2(_06728_),
    .B1(_13629_),
    .Y(_06729_));
 sky130_fd_sc_hd__and3_1 _18290_ (.A(_13629_),
    .B(_06726_),
    .C(_06728_),
    .X(_06730_));
 sky130_fd_sc_hd__or3_4 _18291_ (.A(net524),
    .B(_06729_),
    .C(_06730_),
    .X(_06731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1132 ();
 sky130_fd_sc_hd__clkinv_4 _18293_ (.A(_06731_),
    .Y(\hash.CA1.S1.X[8] ));
 sky130_fd_sc_hd__o21ai_1 _18294_ (.A1(\hash.CA1.S1.X[6] ),
    .A2(_06715_),
    .B1(\hash.CA1.S1.X[7] ),
    .Y(_06733_));
 sky130_fd_sc_hd__xnor2_2 _18295_ (.A(\hash.CA1.S1.X[8] ),
    .B(_06733_),
    .Y(_00811_));
 sky130_fd_sc_hd__o211ai_1 _18296_ (.A1(_13624_),
    .A2(_06716_),
    .B1(_13627_),
    .C1(_13629_),
    .Y(_06734_));
 sky130_fd_sc_hd__a21oi_2 _18297_ (.A1(_13629_),
    .A2(_13626_),
    .B1(_13628_),
    .Y(_06735_));
 sky130_fd_sc_hd__o21ai_1 _18298_ (.A1(_06719_),
    .A2(_06734_),
    .B1(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__xor2_2 _18299_ (.A(_13631_),
    .B(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__nor2_8 _18300_ (.A(net524),
    .B(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__clkinv_2 _18301_ (.A(_06738_),
    .Y(\hash.CA1.S1.X[9] ));
 sky130_fd_sc_hd__nand3_2 _18302_ (.A(\hash.CA1.S1.X[7] ),
    .B(_06723_),
    .C(\hash.CA1.S1.X[8] ),
    .Y(_06739_));
 sky130_fd_sc_hd__xnor2_1 _18303_ (.A(_06738_),
    .B(_06739_),
    .Y(_00812_));
 sky130_fd_sc_hd__nor4b_2 _18304_ (.A(_13628_),
    .B(_13630_),
    .C(_06730_),
    .D_N(_13633_),
    .Y(_06740_));
 sky130_fd_sc_hd__nor2b_1 _18305_ (.A(_13633_),
    .B_N(_13631_),
    .Y(_06741_));
 sky130_fd_sc_hd__and2_0 _18306_ (.A(_06730_),
    .B(_06741_),
    .X(_06742_));
 sky130_fd_sc_hd__inv_1 _18307_ (.A(_13630_),
    .Y(_06743_));
 sky130_fd_sc_hd__nor3b_1 _18308_ (.A(_13631_),
    .B(_13630_),
    .C_N(_13633_),
    .Y(_06744_));
 sky130_fd_sc_hd__a21oi_1 _18309_ (.A1(_13628_),
    .A2(_06741_),
    .B1(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__o21ai_2 _18310_ (.A1(_13633_),
    .A2(_06743_),
    .B1(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__nor3_4 _18311_ (.A(_06740_),
    .B(_06742_),
    .C(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__nor2_8 _18312_ (.A(net524),
    .B(_06747_),
    .Y(\hash.CA1.S1.X[10] ));
 sky130_fd_sc_hd__a311oi_4 _18313_ (.A1(_06700_),
    .A2(_06713_),
    .A3(_06714_),
    .B1(_06722_),
    .C1(_06731_),
    .Y(_06748_));
 sky130_fd_sc_hd__nor2_1 _18314_ (.A(\hash.CA1.S1.X[9] ),
    .B(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__xnor2_2 _18315_ (.A(\hash.CA1.S1.X[10] ),
    .B(_06749_),
    .Y(_00782_));
 sky130_fd_sc_hd__o211ai_4 _18316_ (.A1(_06702_),
    .A2(_06703_),
    .B1(_06704_),
    .C1(_06718_),
    .Y(_06750_));
 sky130_fd_sc_hd__and3_1 _18317_ (.A(_13631_),
    .B(_13629_),
    .C(_13633_),
    .X(_06751_));
 sky130_fd_sc_hd__nor3b_2 _18318_ (.A(_06724_),
    .B(_06725_),
    .C_N(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__nand2_1 _18319_ (.A(_13631_),
    .B(_13633_),
    .Y(_06753_));
 sky130_fd_sc_hd__a21oi_1 _18320_ (.A1(_13633_),
    .A2(_13630_),
    .B1(_13632_),
    .Y(_06754_));
 sky130_fd_sc_hd__o21ai_4 _18321_ (.A1(_06735_),
    .A2(_06753_),
    .B1(_06754_),
    .Y(_06755_));
 sky130_fd_sc_hd__a21oi_1 _18322_ (.A1(_06750_),
    .A2(_06752_),
    .B1(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__xnor2_1 _18323_ (.A(_13635_),
    .B(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_4 _18324_ (.A(_06210_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__clkinv_2 _18325_ (.A(_06758_),
    .Y(\hash.CA1.S1.X[11] ));
 sky130_fd_sc_hd__nand2_1 _18326_ (.A(_06738_),
    .B(_06739_),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_1 _18327_ (.A(_06759_),
    .B(\hash.CA1.S1.X[10] ),
    .Y(_06760_));
 sky130_fd_sc_hd__xnor2_1 _18328_ (.A(\hash.CA1.S1.X[11] ),
    .B(_06760_),
    .Y(_00783_));
 sky130_fd_sc_hd__nor2b_1 _18329_ (.A(net524),
    .B_N(_13637_),
    .Y(_06761_));
 sky130_fd_sc_hd__nor2_1 _18330_ (.A(net524),
    .B(_13637_),
    .Y(_06762_));
 sky130_fd_sc_hd__clkinvlp_4 _18331_ (.A(_13635_),
    .Y(_06763_));
 sky130_fd_sc_hd__a31oi_4 _18332_ (.A1(_06726_),
    .A2(_06728_),
    .A3(_06751_),
    .B1(_13632_),
    .Y(_06764_));
 sky130_fd_sc_hd__nand2_1 _18333_ (.A(_13631_),
    .B(_13628_),
    .Y(_06765_));
 sky130_fd_sc_hd__nand2_1 _18334_ (.A(_06743_),
    .B(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__a31oi_4 _18335_ (.A1(_13633_),
    .A2(_13635_),
    .A3(_06766_),
    .B1(_13634_),
    .Y(_06767_));
 sky130_fd_sc_hd__o21a_1 _18336_ (.A1(_06763_),
    .A2(_06764_),
    .B1(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__mux2i_4 _18337_ (.A0(_06761_),
    .A1(_06762_),
    .S(_06768_),
    .Y(\hash.CA1.S1.X[12] ));
 sky130_fd_sc_hd__or3_4 _18338_ (.A(_06740_),
    .B(_06742_),
    .C(_06746_),
    .X(_06769_));
 sky130_fd_sc_hd__o211ai_4 _18339_ (.A1(\hash.CA1.S1.X[9] ),
    .A2(_06748_),
    .B1(\hash.CA1.S1.X[11] ),
    .C1(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__xor2_2 _18340_ (.A(\hash.CA1.S1.X[12] ),
    .B(_06770_),
    .X(_00784_));
 sky130_fd_sc_hd__nand2_1 _18341_ (.A(_13637_),
    .B(_13635_),
    .Y(_06771_));
 sky130_fd_sc_hd__a21oi_1 _18342_ (.A1(_13637_),
    .A2(_13634_),
    .B1(_13636_),
    .Y(_06772_));
 sky130_fd_sc_hd__o21ai_0 _18343_ (.A1(_06756_),
    .A2(_06771_),
    .B1(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__xor2_1 _18344_ (.A(_13639_),
    .B(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__nand2_2 _18345_ (.A(_06210_),
    .B(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__clkinv_4 _18346_ (.A(_06775_),
    .Y(\hash.CA1.S1.X[13] ));
 sky130_fd_sc_hd__a31oi_1 _18347_ (.A1(_06759_),
    .A2(_06769_),
    .A3(\hash.CA1.S1.X[11] ),
    .B1(\hash.CA1.S1.X[12] ),
    .Y(_06776_));
 sky130_fd_sc_hd__xnor2_1 _18348_ (.A(\hash.CA1.S1.X[13] ),
    .B(_06776_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand3_1 _18349_ (.A(_13637_),
    .B(_13641_),
    .C(_13639_),
    .Y(_06777_));
 sky130_fd_sc_hd__a21oi_1 _18350_ (.A1(_13639_),
    .A2(_13636_),
    .B1(_13638_),
    .Y(_06778_));
 sky130_fd_sc_hd__nor2_1 _18351_ (.A(net524),
    .B(_13641_),
    .Y(_06779_));
 sky130_fd_sc_hd__o2111ai_2 _18352_ (.A1(_06763_),
    .A2(_06764_),
    .B1(_06778_),
    .C1(_06779_),
    .D1(_06767_),
    .Y(_06780_));
 sky130_fd_sc_hd__a21o_1 _18353_ (.A1(_13639_),
    .A2(_13636_),
    .B1(_13638_),
    .X(_06781_));
 sky130_fd_sc_hd__a2111oi_1 _18354_ (.A1(_13637_),
    .A2(_13639_),
    .B1(_06781_),
    .C1(_13641_),
    .D1(net524),
    .Y(_06782_));
 sky130_fd_sc_hd__a31oi_2 _18355_ (.A1(_06210_),
    .A2(_13641_),
    .A3(_06781_),
    .B1(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__o311ai_4 _18356_ (.A1(net524),
    .A2(_06768_),
    .A3(_06777_),
    .B1(_06780_),
    .C1(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__clkinv_2 _18357_ (.A(_06784_),
    .Y(\hash.CA1.S1.X[14] ));
 sky130_fd_sc_hd__nand2b_1 _18358_ (.A_N(\hash.CA1.S1.X[12] ),
    .B(_06770_),
    .Y(_06785_));
 sky130_fd_sc_hd__nand2_1 _18359_ (.A(_06785_),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_06786_));
 sky130_fd_sc_hd__xnor2_2 _18360_ (.A(_06784_),
    .B(_06786_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand2_1 _18361_ (.A(_13641_),
    .B(_13639_),
    .Y(_06787_));
 sky130_fd_sc_hd__a21oi_1 _18362_ (.A1(_13641_),
    .A2(_13638_),
    .B1(_13640_),
    .Y(_06788_));
 sky130_fd_sc_hd__o21a_1 _18363_ (.A1(_06772_),
    .A2(_06787_),
    .B1(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__o31a_1 _18364_ (.A1(_06763_),
    .A2(_06756_),
    .A3(_06777_),
    .B1(_06789_),
    .X(_06790_));
 sky130_fd_sc_hd__xnor2_2 _18365_ (.A(_13643_),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__nand2_8 _18366_ (.A(_06210_),
    .B(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__a2111oi_0 _18367_ (.A1(_06738_),
    .A2(_06739_),
    .B1(_06747_),
    .C1(_06758_),
    .D1(_06775_),
    .Y(_06793_));
 sky130_fd_sc_hd__a211o_2 _18368_ (.A1(\hash.CA1.S1.X[12] ),
    .A2(\hash.CA1.S1.X[13] ),
    .B1(\hash.CA1.S1.X[14] ),
    .C1(_06793_),
    .X(_06794_));
 sky130_fd_sc_hd__xnor2_2 _18369_ (.A(_06792_),
    .B(_06794_),
    .Y(_00787_));
 sky130_fd_sc_hd__inv_1 _18370_ (.A(_13643_),
    .Y(_06795_));
 sky130_fd_sc_hd__o21ai_0 _18371_ (.A1(_13637_),
    .A2(_13636_),
    .B1(_13639_),
    .Y(_06796_));
 sky130_fd_sc_hd__nand2b_1 _18372_ (.A_N(_13638_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__a21oi_1 _18373_ (.A1(_13641_),
    .A2(_06797_),
    .B1(_13640_),
    .Y(_06798_));
 sky130_fd_sc_hd__o21bai_2 _18374_ (.A1(_06795_),
    .A2(_06798_),
    .B1_N(_13642_),
    .Y(_06799_));
 sky130_fd_sc_hd__a211oi_2 _18375_ (.A1(_13643_),
    .A2(_13640_),
    .B1(_13642_),
    .C1(_06781_),
    .Y(_06800_));
 sky130_fd_sc_hd__o211ai_4 _18376_ (.A1(_06763_),
    .A2(_06764_),
    .B1(_06800_),
    .C1(_06767_),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_1 _18377_ (.A(_06799_),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__xnor2_1 _18378_ (.A(_13645_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__and2_4 _18379_ (.A(_06210_),
    .B(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1131 ();
 sky130_fd_sc_hd__nor2_1 _18381_ (.A(\hash.CA1.S1.X[12] ),
    .B(\hash.CA1.S1.X[14] ),
    .Y(_06805_));
 sky130_fd_sc_hd__a22o_2 _18382_ (.A1(_06775_),
    .A2(_06784_),
    .B1(_06805_),
    .B2(_06770_),
    .X(_06806_));
 sky130_fd_sc_hd__nor2_1 _18383_ (.A(_06806_),
    .B(_06792_),
    .Y(_06807_));
 sky130_fd_sc_hd__xor2_2 _18384_ (.A(_06804_),
    .B(_06807_),
    .X(_00788_));
 sky130_fd_sc_hd__inv_2 _18385_ (.A(_06792_),
    .Y(\hash.CA1.S1.X[15] ));
 sky130_fd_sc_hd__a21o_1 _18386_ (.A1(_13645_),
    .A2(_13642_),
    .B1(_13644_),
    .X(_06808_));
 sky130_fd_sc_hd__nor3_4 _18387_ (.A(_06795_),
    .B(_06771_),
    .C(_06787_),
    .Y(_06809_));
 sky130_fd_sc_hd__nand3_2 _18388_ (.A(_06750_),
    .B(_06752_),
    .C(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__o21ai_1 _18389_ (.A1(_06772_),
    .A2(_06787_),
    .B1(_06788_),
    .Y(_06811_));
 sky130_fd_sc_hd__a22oi_4 _18390_ (.A1(_13643_),
    .A2(_06811_),
    .B1(_06809_),
    .B2(_06755_),
    .Y(_06812_));
 sky130_fd_sc_hd__a21boi_0 _18391_ (.A1(_06810_),
    .A2(_06812_),
    .B1_N(_13649_),
    .Y(_06813_));
 sky130_fd_sc_hd__o21ai_1 _18392_ (.A1(_06808_),
    .A2(_06813_),
    .B1(_13647_),
    .Y(_06814_));
 sky130_fd_sc_hd__or3_1 _18393_ (.A(_13647_),
    .B(_06808_),
    .C(_06813_),
    .X(_06815_));
 sky130_fd_sc_hd__a21oi_4 _18394_ (.A1(_06814_),
    .A2(_06815_),
    .B1(net523),
    .Y(_06816_));
 sky130_fd_sc_hd__inv_1 _18395_ (.A(_06816_),
    .Y(\hash.CA1.S1.X[17] ));
 sky130_fd_sc_hd__nand3_1 _18396_ (.A(\hash.CA1.S1.X[15] ),
    .B(_06794_),
    .C(_06804_),
    .Y(_06817_));
 sky130_fd_sc_hd__xnor2_2 _18397_ (.A(_06816_),
    .B(_06817_),
    .Y(_00789_));
 sky130_fd_sc_hd__a31o_1 _18398_ (.A1(_13649_),
    .A2(_06799_),
    .A3(_06801_),
    .B1(_13644_),
    .X(_06818_));
 sky130_fd_sc_hd__a21o_2 _18399_ (.A1(_13647_),
    .A2(_06818_),
    .B1(_13646_),
    .X(_06819_));
 sky130_fd_sc_hd__xor2_4 _18400_ (.A(_13651_),
    .B(_06819_),
    .X(_06820_));
 sky130_fd_sc_hd__nor2_4 _18401_ (.A(net523),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__inv_1 _18402_ (.A(_06821_),
    .Y(\hash.CA1.S1.X[18] ));
 sky130_fd_sc_hd__nand3_1 _18403_ (.A(_06210_),
    .B(\hash.CA1.S1.X[15] ),
    .C(_06803_),
    .Y(_06822_));
 sky130_fd_sc_hd__o21ai_1 _18404_ (.A1(_06806_),
    .A2(_06822_),
    .B1(_06816_),
    .Y(_06823_));
 sky130_fd_sc_hd__xor2_2 _18405_ (.A(_06821_),
    .B(_06823_),
    .X(_00790_));
 sky130_fd_sc_hd__a21o_1 _18406_ (.A1(_13647_),
    .A2(_06808_),
    .B1(_13646_),
    .X(_06824_));
 sky130_fd_sc_hd__a21o_1 _18407_ (.A1(_13651_),
    .A2(_06824_),
    .B1(_13650_),
    .X(_06825_));
 sky130_fd_sc_hd__and3_1 _18408_ (.A(_13647_),
    .B(_13649_),
    .C(_13651_),
    .X(_06826_));
 sky130_fd_sc_hd__a21boi_4 _18409_ (.A1(_06810_),
    .A2(_06812_),
    .B1_N(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__o21ai_1 _18410_ (.A1(_06825_),
    .A2(_06827_),
    .B1(_13653_),
    .Y(_06828_));
 sky130_fd_sc_hd__or3_1 _18411_ (.A(_13653_),
    .B(_06825_),
    .C(_06827_),
    .X(_06829_));
 sky130_fd_sc_hd__a21oi_4 _18412_ (.A1(_06828_),
    .A2(_06829_),
    .B1(net523),
    .Y(_06830_));
 sky130_fd_sc_hd__inv_1 _18413_ (.A(_06830_),
    .Y(\hash.CA1.S1.X[19] ));
 sky130_fd_sc_hd__a31oi_4 _18414_ (.A1(\hash.CA1.S1.X[15] ),
    .A2(_06794_),
    .A3(_06804_),
    .B1(_06820_),
    .Y(_06831_));
 sky130_fd_sc_hd__nand2_1 _18415_ (.A(_06816_),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__xnor2_2 _18416_ (.A(\hash.CA1.S1.X[19] ),
    .B(_06832_),
    .Y(_00791_));
 sky130_fd_sc_hd__a21oi_1 _18417_ (.A1(_13647_),
    .A2(_13644_),
    .B1(_13646_),
    .Y(_06833_));
 sky130_fd_sc_hd__nor2b_1 _18418_ (.A(_06833_),
    .B_N(_13651_),
    .Y(_06834_));
 sky130_fd_sc_hd__o21ai_0 _18419_ (.A1(_13650_),
    .A2(_06834_),
    .B1(_13653_),
    .Y(_06835_));
 sky130_fd_sc_hd__nand2b_1 _18420_ (.A_N(_13652_),
    .B(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__a41o_2 _18421_ (.A1(_13653_),
    .A2(_06799_),
    .A3(_06801_),
    .A4(_06826_),
    .B1(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__xnor2_2 _18422_ (.A(_13655_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_8 _18423_ (.A(net523),
    .B(_06838_),
    .Y(\hash.CA1.S1.X[20] ));
 sky130_fd_sc_hd__xnor2_2 _18424_ (.A(_13651_),
    .B(_06819_),
    .Y(_06839_));
 sky130_fd_sc_hd__and2_2 _18425_ (.A(_06816_),
    .B(_06830_),
    .X(_06840_));
 sky130_fd_sc_hd__o211a_2 _18426_ (.A1(_06806_),
    .A2(_06822_),
    .B1(_06839_),
    .C1(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__xnor2_1 _18427_ (.A(\hash.CA1.S1.X[20] ),
    .B(_06841_),
    .Y(_00793_));
 sky130_fd_sc_hd__inv_1 _18428_ (.A(_13657_),
    .Y(_06842_));
 sky130_fd_sc_hd__a21oi_4 _18429_ (.A1(_13655_),
    .A2(_13652_),
    .B1(_13654_),
    .Y(_06843_));
 sky130_fd_sc_hd__nand2_1 _18430_ (.A(_13653_),
    .B(_13659_),
    .Y(_06844_));
 sky130_fd_sc_hd__o21bai_1 _18431_ (.A1(_06825_),
    .A2(_06827_),
    .B1_N(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__and3_1 _18432_ (.A(_06842_),
    .B(_06843_),
    .C(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__a21oi_1 _18433_ (.A1(_06843_),
    .A2(_06845_),
    .B1(_06842_),
    .Y(_06847_));
 sky130_fd_sc_hd__nor3_4 _18434_ (.A(net523),
    .B(_06846_),
    .C(_06847_),
    .Y(\hash.CA1.S1.X[21] ));
 sky130_fd_sc_hd__nand2_1 _18435_ (.A(_06831_),
    .B(_06840_),
    .Y(_06848_));
 sky130_fd_sc_hd__nand2_1 _18436_ (.A(\hash.CA1.S1.X[20] ),
    .B(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__xnor2_2 _18437_ (.A(\hash.CA1.S1.X[21] ),
    .B(_06849_),
    .Y(_00794_));
 sky130_fd_sc_hd__a21oi_1 _18438_ (.A1(_13657_),
    .A2(_13654_),
    .B1(_13656_),
    .Y(_06850_));
 sky130_fd_sc_hd__inv_1 _18439_ (.A(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__a31oi_2 _18440_ (.A1(_13659_),
    .A2(_13663_),
    .A3(_06837_),
    .B1(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__xnor2_2 _18441_ (.A(net1025),
    .B(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__and2_4 _18442_ (.A(_06210_),
    .B(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1130 ();
 sky130_fd_sc_hd__nand2_1 _18444_ (.A(\hash.CA1.S1.X[20] ),
    .B(\hash.CA1.S1.X[21] ),
    .Y(_06855_));
 sky130_fd_sc_hd__nor2_1 _18445_ (.A(_06841_),
    .B(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__xor2_2 _18446_ (.A(_06854_),
    .B(_06856_),
    .X(_00795_));
 sky130_fd_sc_hd__nand2_2 _18447_ (.A(_13663_),
    .B(_13667_),
    .Y(_06857_));
 sky130_fd_sc_hd__nor2_4 _18448_ (.A(_06844_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__a21oi_2 _18449_ (.A1(_13656_),
    .A2(_13661_),
    .B1(_13660_),
    .Y(_06859_));
 sky130_fd_sc_hd__o21ai_2 _18450_ (.A1(_06843_),
    .A2(_06857_),
    .B1(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__a21o_1 _18451_ (.A1(_06825_),
    .A2(_06858_),
    .B1(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__a21oi_4 _18452_ (.A1(_06827_),
    .A2(_06858_),
    .B1(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__xnor2_2 _18453_ (.A(_13665_),
    .B(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__nand2_4 _18454_ (.A(_06210_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__clkinv_2 _18455_ (.A(_06864_),
    .Y(\hash.CA1.S1.X[23] ));
 sky130_fd_sc_hd__nand4_1 _18456_ (.A(_06210_),
    .B(\hash.CA1.S1.X[20] ),
    .C(\hash.CA1.S1.X[21] ),
    .D(_06853_),
    .Y(_06865_));
 sky130_fd_sc_hd__nand2b_1 _18457_ (.A_N(_06865_),
    .B(_06848_),
    .Y(_06866_));
 sky130_fd_sc_hd__xnor2_2 _18458_ (.A(\hash.CA1.S1.X[23] ),
    .B(_06866_),
    .Y(_00796_));
 sky130_fd_sc_hd__nor2b_1 _18459_ (.A(net523),
    .B_N(_13669_),
    .Y(_06867_));
 sky130_fd_sc_hd__nor2_1 _18460_ (.A(net523),
    .B(_13669_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand2_1 _18461_ (.A(_13659_),
    .B(_13663_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand2_1 _18462_ (.A(_13667_),
    .B(_13671_),
    .Y(_06870_));
 sky130_fd_sc_hd__nor2_1 _18463_ (.A(_06869_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__a21oi_1 _18464_ (.A1(_13665_),
    .A2(_13660_),
    .B1(_13664_),
    .Y(_06872_));
 sky130_fd_sc_hd__o21ai_1 _18465_ (.A1(_06850_),
    .A2(_06870_),
    .B1(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__a21oi_4 _18466_ (.A1(_06837_),
    .A2(_06871_),
    .B1(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__mux2i_4 _18467_ (.A0(_06867_),
    .A1(_06868_),
    .S(net1110),
    .Y(\hash.CA1.S1.X[24] ));
 sky130_fd_sc_hd__nor3_2 _18468_ (.A(_06841_),
    .B(_06864_),
    .C(_06865_),
    .Y(_06875_));
 sky130_fd_sc_hd__xnor2_1 _18469_ (.A(\hash.CA1.S1.X[24] ),
    .B(_06875_),
    .Y(_00797_));
 sky130_fd_sc_hd__a211oi_1 _18470_ (.A1(_06831_),
    .A2(_06840_),
    .B1(_06864_),
    .C1(_06865_),
    .Y(_06876_));
 sky130_fd_sc_hd__nor2_1 _18471_ (.A(\hash.CA1.S1.X[24] ),
    .B(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__nand2_1 _18472_ (.A(_13669_),
    .B(_13671_),
    .Y(_06878_));
 sky130_fd_sc_hd__a21oi_1 _18473_ (.A1(_13669_),
    .A2(_13664_),
    .B1(_13668_),
    .Y(_06879_));
 sky130_fd_sc_hd__o21ai_4 _18474_ (.A1(_06862_),
    .A2(_06878_),
    .B1(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__xnor2_4 _18475_ (.A(net1107),
    .B(_13673_),
    .Y(_06881_));
 sky130_fd_sc_hd__nor2_8 _18476_ (.A(net523),
    .B(_06881_),
    .Y(\hash.CA1.S1.X[25] ));
 sky130_fd_sc_hd__xnor2_1 _18477_ (.A(_06877_),
    .B(net1020),
    .Y(_00798_));
 sky130_fd_sc_hd__nand2_1 _18478_ (.A(_13669_),
    .B(_13677_),
    .Y(_06882_));
 sky130_fd_sc_hd__a21oi_1 _18479_ (.A1(_13673_),
    .A2(_13668_),
    .B1(_13672_),
    .Y(_06883_));
 sky130_fd_sc_hd__o21ai_2 _18480_ (.A1(_06874_),
    .A2(_06882_),
    .B1(_06883_),
    .Y(_06884_));
 sky130_fd_sc_hd__xor2_2 _18481_ (.A(_13675_),
    .B(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__nand2_8 _18482_ (.A(_06210_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__clkinv_4 _18483_ (.A(_06886_),
    .Y(\hash.CA1.S1.X[26] ));
 sky130_fd_sc_hd__o21ai_1 _18484_ (.A1(\hash.CA1.S1.X[24] ),
    .A2(_06875_),
    .B1(\hash.CA1.S1.X[25] ),
    .Y(_06887_));
 sky130_fd_sc_hd__xnor2_1 _18485_ (.A(\hash.CA1.S1.X[26] ),
    .B(_06887_),
    .Y(_00799_));
 sky130_fd_sc_hd__a21o_1 _18486_ (.A1(_13675_),
    .A2(_13672_),
    .B1(_13674_),
    .X(_06888_));
 sky130_fd_sc_hd__a311oi_2 _18487_ (.A1(_13677_),
    .A2(_06880_),
    .A3(_13681_),
    .B1(_06888_),
    .C1(_13679_),
    .Y(_06889_));
 sky130_fd_sc_hd__nand2_1 _18488_ (.A(_13677_),
    .B(_13681_),
    .Y(_06890_));
 sky130_fd_sc_hd__nor2_1 _18489_ (.A(_06878_),
    .B(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2_1 _18490_ (.A(_13679_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__nor3b_2 _18491_ (.A(_06879_),
    .B(_06890_),
    .C_N(_13679_),
    .Y(_06893_));
 sky130_fd_sc_hd__a21oi_2 _18492_ (.A1(_13679_),
    .A2(_06888_),
    .B1(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__o21ai_4 _18493_ (.A1(net1108),
    .A2(_06892_),
    .B1(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__or3_4 _18494_ (.A(net523),
    .B(_06889_),
    .C(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1129 ();
 sky130_fd_sc_hd__inv_1 _18496_ (.A(net1027),
    .Y(\hash.CA1.S1.X[27] ));
 sky130_fd_sc_hd__nand2_1 _18497_ (.A(net1020),
    .B(\hash.CA1.S1.X[26] ),
    .Y(_06898_));
 sky130_fd_sc_hd__nor2_1 _18498_ (.A(_06877_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__xnor2_1 _18499_ (.A(net1026),
    .B(_06899_),
    .Y(_00800_));
 sky130_fd_sc_hd__a21o_1 _18500_ (.A1(_13679_),
    .A2(_13674_),
    .B1(_13678_),
    .X(_06900_));
 sky130_fd_sc_hd__a31oi_4 _18501_ (.A1(_06884_),
    .A2(_13679_),
    .A3(_13675_),
    .B1(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__xnor2_4 _18502_ (.A(_13683_),
    .B(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__nor2_8 _18503_ (.A(net522),
    .B(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__clkinvlp_4 _18504_ (.A(_06903_),
    .Y(\hash.CA1.S1.X[28] ));
 sky130_fd_sc_hd__nor3_1 _18505_ (.A(_06886_),
    .B(_06887_),
    .C(net1027),
    .Y(_06904_));
 sky130_fd_sc_hd__xnor2_1 _18506_ (.A(\hash.CA1.S1.X[28] ),
    .B(_06904_),
    .Y(_00801_));
 sky130_fd_sc_hd__o21ai_1 _18507_ (.A1(_13678_),
    .A2(_06895_),
    .B1(_13683_),
    .Y(_06905_));
 sky130_fd_sc_hd__nor2_1 _18508_ (.A(_13685_),
    .B(_13682_),
    .Y(_06906_));
 sky130_fd_sc_hd__nor2_1 _18509_ (.A(_13678_),
    .B(_13682_),
    .Y(_06907_));
 sky130_fd_sc_hd__o211ai_2 _18510_ (.A1(net1108),
    .A2(_06892_),
    .B1(_06907_),
    .C1(_06894_),
    .Y(_06908_));
 sky130_fd_sc_hd__o21a_1 _18511_ (.A1(_13683_),
    .A2(_13682_),
    .B1(_13685_),
    .X(_06909_));
 sky130_fd_sc_hd__a221o_4 _18512_ (.A1(_06906_),
    .A2(_06905_),
    .B1(_06909_),
    .B2(_06908_),
    .C1(net523),
    .X(_06910_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1128 ();
 sky130_fd_sc_hd__o31ai_1 _18514_ (.A1(_06877_),
    .A2(net1027),
    .A3(_06898_),
    .B1(_06903_),
    .Y(_06912_));
 sky130_fd_sc_hd__xnor2_1 _18515_ (.A(_06910_),
    .B(_06912_),
    .Y(_00802_));
 sky130_fd_sc_hd__inv_1 _18516_ (.A(_06910_),
    .Y(\hash.CA1.S1.X[29] ));
 sky130_fd_sc_hd__nand2_1 _18517_ (.A(_13685_),
    .B(_13683_),
    .Y(_06913_));
 sky130_fd_sc_hd__a21oi_1 _18518_ (.A1(_13685_),
    .A2(_13682_),
    .B1(_13684_),
    .Y(_06914_));
 sky130_fd_sc_hd__o21ai_1 _18519_ (.A1(_06901_),
    .A2(_06913_),
    .B1(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__xor2_2 _18520_ (.A(_13687_),
    .B(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__nor2_8 _18521_ (.A(net522),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__inv_1 _18522_ (.A(_06917_),
    .Y(\hash.CA1.S1.X[30] ));
 sky130_fd_sc_hd__o21a_1 _18523_ (.A1(\hash.CA1.S1.X[28] ),
    .A2(_06904_),
    .B1(\hash.CA1.S1.X[29] ),
    .X(_06918_));
 sky130_fd_sc_hd__xnor2_1 _18524_ (.A(\hash.CA1.S1.X[30] ),
    .B(_06918_),
    .Y(_00804_));
 sky130_fd_sc_hd__a21o_1 _18525_ (.A1(_06908_),
    .A2(_06909_),
    .B1(_13684_),
    .X(_06919_));
 sky130_fd_sc_hd__a21oi_2 _18526_ (.A1(_06919_),
    .A2(_13687_),
    .B1(_13686_),
    .Y(_06920_));
 sky130_fd_sc_hd__xor3_1 _18527_ (.A(\hash.CA2.p5[31] ),
    .B(_06446_),
    .C(_06920_),
    .X(_06921_));
 sky130_fd_sc_hd__and2_4 _18528_ (.A(_06210_),
    .B(_06921_),
    .X(_06922_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1127 ();
 sky130_fd_sc_hd__nand4_1 _18530_ (.A(net1020),
    .B(\hash.CA1.S1.X[26] ),
    .C(\hash.CA1.S1.X[27] ),
    .D(\hash.CA1.S1.X[29] ),
    .Y(_06923_));
 sky130_fd_sc_hd__o221a_1 _18531_ (.A1(_06903_),
    .A2(_06910_),
    .B1(_06923_),
    .B2(_06877_),
    .C1(_06917_),
    .X(_06924_));
 sky130_fd_sc_hd__xnor2_1 _18532_ (.A(_06922_),
    .B(_06924_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand2_2 _18533_ (.A(net519),
    .B(\hash.CA2.b_dash[2] ),
    .Y(_12837_));
 sky130_fd_sc_hd__inv_1 _18534_ (.A(_12837_),
    .Y(_14025_));
 sky130_fd_sc_hd__nor2_4 _18535_ (.A(net520),
    .B(\hash.CA2.b_dash[3] ),
    .Y(_12845_));
 sky130_fd_sc_hd__xor2_1 _18536_ (.A(_14026_),
    .B(_12845_),
    .X(_00772_));
 sky130_fd_sc_hd__nor2_2 _18537_ (.A(net520),
    .B(\hash.CA2.b_dash[4] ),
    .Y(_12850_));
 sky130_fd_sc_hd__a21oi_1 _18538_ (.A1(\hash.CA2.b_dash[1] ),
    .A2(\hash.CA2.b_dash[2] ),
    .B1(\hash.CA2.b_dash[3] ),
    .Y(_06925_));
 sky130_fd_sc_hd__xnor2_1 _18539_ (.A(\hash.CA2.b_dash[4] ),
    .B(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__nand2_1 _18540_ (.A(net519),
    .B(_06926_),
    .Y(_00774_));
 sky130_fd_sc_hd__or2_4 _18541_ (.A(net520),
    .B(\hash.CA2.b_dash[5] ),
    .X(_12855_));
 sky130_fd_sc_hd__nor4_1 _18542_ (.A(net520),
    .B(\hash.CA2.b_dash[3] ),
    .C(\hash.CA2.b_dash[4] ),
    .D(_14026_),
    .Y(_06927_));
 sky130_fd_sc_hd__xor2_1 _18543_ (.A(_12855_),
    .B(_06927_),
    .X(_00775_));
 sky130_fd_sc_hd__nand2b_4 _18544_ (.A_N(net520),
    .B(\hash.CA2.b_dash[6] ),
    .Y(_12863_));
 sky130_fd_sc_hd__nor3_1 _18545_ (.A(net520),
    .B(\hash.CA2.b_dash[3] ),
    .C(\hash.CA2.b_dash[4] ),
    .Y(_06928_));
 sky130_fd_sc_hd__a21oi_1 _18546_ (.A1(\hash.CA2.b_dash[1] ),
    .A2(\hash.CA2.b_dash[2] ),
    .B1(\hash.CA2.b_dash[5] ),
    .Y(_06929_));
 sky130_fd_sc_hd__nand2_1 _18547_ (.A(_06928_),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__xnor2_1 _18548_ (.A(_12863_),
    .B(_06930_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand2b_4 _18549_ (.A_N(net520),
    .B(\hash.CA2.b_dash[7] ),
    .Y(_12872_));
 sky130_fd_sc_hd__nor4_2 _18550_ (.A(\hash.CA2.b_dash[3] ),
    .B(\hash.CA2.b_dash[4] ),
    .C(\hash.CA2.b_dash[5] ),
    .D(_14026_),
    .Y(_06931_));
 sky130_fd_sc_hd__nor2_1 _18551_ (.A(_12863_),
    .B(_06931_),
    .Y(_06932_));
 sky130_fd_sc_hd__mux2i_1 _18552_ (.A0(_12872_),
    .A1(\hash.CA2.b_dash[7] ),
    .S(_06932_),
    .Y(_00777_));
 sky130_fd_sc_hd__nor2_4 _18553_ (.A(net520),
    .B(\hash.CA2.b_dash[8] ),
    .Y(_12879_));
 sky130_fd_sc_hd__inv_1 _18554_ (.A(\hash.CA2.b_dash[7] ),
    .Y(_06933_));
 sky130_fd_sc_hd__a211oi_2 _18555_ (.A1(_06928_),
    .A2(_06929_),
    .B1(_12863_),
    .C1(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__xor2_1 _18556_ (.A(_12879_),
    .B(_06934_),
    .X(_00778_));
 sky130_fd_sc_hd__nand2b_1 _18557_ (.A_N(\hash.CA2.b_dash[5] ),
    .B(_06927_),
    .Y(_06935_));
 sky130_fd_sc_hd__nand3_1 _18558_ (.A(\hash.CA2.b_dash[6] ),
    .B(\hash.CA2.b_dash[7] ),
    .C(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__nand2_4 _18559_ (.A(net519),
    .B(\hash.CA2.b_dash[9] ),
    .Y(_12885_));
 sky130_fd_sc_hd__a21oi_1 _18560_ (.A1(_12879_),
    .A2(_06936_),
    .B1(_12885_),
    .Y(_06937_));
 sky130_fd_sc_hd__nand2_1 _18561_ (.A(_12879_),
    .B(_06936_),
    .Y(_06938_));
 sky130_fd_sc_hd__nor2_1 _18562_ (.A(\hash.CA2.b_dash[9] ),
    .B(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__nor2_1 _18563_ (.A(_06937_),
    .B(_06939_),
    .Y(_00779_));
 sky130_fd_sc_hd__nor2_4 _18564_ (.A(net520),
    .B(\hash.CA2.b_dash[10] ),
    .Y(_12894_));
 sky130_fd_sc_hd__o21bai_1 _18565_ (.A1(\hash.CA2.b_dash[8] ),
    .A2(_06934_),
    .B1_N(_12885_),
    .Y(_06940_));
 sky130_fd_sc_hd__xnor2_1 _18566_ (.A(_12894_),
    .B(_06940_),
    .Y(_00780_));
 sky130_fd_sc_hd__nor2_4 _18567_ (.A(net520),
    .B(_04826_),
    .Y(_12903_));
 sky130_fd_sc_hd__inv_1 _18568_ (.A(\hash.CA2.b_dash[8] ),
    .Y(_06941_));
 sky130_fd_sc_hd__o31ai_1 _18569_ (.A1(_12863_),
    .A2(_06931_),
    .A3(_12872_),
    .B1(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__a211o_1 _18570_ (.A1(\hash.CA2.b_dash[9] ),
    .A2(_06942_),
    .B1(\hash.CA2.b_dash[10] ),
    .C1(net520),
    .X(_06943_));
 sky130_fd_sc_hd__xor2_1 _18571_ (.A(_12903_),
    .B(_06943_),
    .X(_00752_));
 sky130_fd_sc_hd__nor2_1 _18572_ (.A(net520),
    .B(\hash.CA2.b_dash[12] ),
    .Y(_06944_));
 sky130_fd_sc_hd__inv_2 _18573_ (.A(_06944_),
    .Y(_12911_));
 sky130_fd_sc_hd__nand2b_1 _18574_ (.A_N(\hash.CA2.b_dash[10] ),
    .B(_06940_),
    .Y(_06945_));
 sky130_fd_sc_hd__nand2_2 _18575_ (.A(_12903_),
    .B(_06945_),
    .Y(_06946_));
 sky130_fd_sc_hd__xnor2_1 _18576_ (.A(_06944_),
    .B(_06946_),
    .Y(_00753_));
 sky130_fd_sc_hd__or2_4 _18577_ (.A(net524),
    .B(\hash.CA2.b_dash[13] ),
    .X(_12917_));
 sky130_fd_sc_hd__a21oi_1 _18578_ (.A1(\hash.CA2.b_dash[9] ),
    .A2(_06938_),
    .B1(\hash.CA2.b_dash[10] ),
    .Y(_06947_));
 sky130_fd_sc_hd__o21ai_2 _18579_ (.A1(_04826_),
    .A2(_06947_),
    .B1(_06944_),
    .Y(_06948_));
 sky130_fd_sc_hd__nor2_2 _18580_ (.A(\hash.CA2.b_dash[12] ),
    .B(_12917_),
    .Y(_06949_));
 sky130_fd_sc_hd__o21ai_1 _18581_ (.A1(\hash.CA2.b_dash[10] ),
    .A2(_06937_),
    .B1(\hash.CA2.b_dash[11] ),
    .Y(_06950_));
 sky130_fd_sc_hd__a22o_1 _18582_ (.A1(_12917_),
    .A2(_06948_),
    .B1(_06949_),
    .B2(_06950_),
    .X(_00754_));
 sky130_fd_sc_hd__nor2_4 _18583_ (.A(net524),
    .B(\hash.CA2.b_dash[14] ),
    .Y(_12923_));
 sky130_fd_sc_hd__nand2_1 _18584_ (.A(\hash.CA2.b_dash[11] ),
    .B(_06945_),
    .Y(_06951_));
 sky130_fd_sc_hd__nand2_1 _18585_ (.A(_06949_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__xor2_1 _18586_ (.A(_12923_),
    .B(_06952_),
    .X(_00755_));
 sky130_fd_sc_hd__nor2_4 _18587_ (.A(net524),
    .B(\hash.CA2.b_dash[15] ),
    .Y(_12930_));
 sky130_fd_sc_hd__nand2_1 _18588_ (.A(_12903_),
    .B(_06943_),
    .Y(_06953_));
 sky130_fd_sc_hd__nand3_2 _18589_ (.A(_06953_),
    .B(_06949_),
    .C(_12923_),
    .Y(_06954_));
 sky130_fd_sc_hd__mux2i_1 _18590_ (.A0(\hash.CA2.b_dash[15] ),
    .A1(_12930_),
    .S(_06954_),
    .Y(_00756_));
 sky130_fd_sc_hd__nand2_4 _18591_ (.A(net519),
    .B(_04863_),
    .Y(_12938_));
 sky130_fd_sc_hd__nor3_1 _18592_ (.A(net524),
    .B(\hash.CA2.b_dash[14] ),
    .C(\hash.CA2.b_dash[15] ),
    .Y(_06955_));
 sky130_fd_sc_hd__nand3_1 _18593_ (.A(_06946_),
    .B(_06949_),
    .C(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__xnor2_1 _18594_ (.A(_12938_),
    .B(_06956_),
    .Y(_00757_));
 sky130_fd_sc_hd__nor2_1 _18595_ (.A(net524),
    .B(\hash.CA2.b_dash[17] ),
    .Y(_06957_));
 sky130_fd_sc_hd__nor4b_1 _18596_ (.A(\hash.CA2.b_dash[13] ),
    .B(_06948_),
    .C(_12938_),
    .D_N(_06955_),
    .Y(_06958_));
 sky130_fd_sc_hd__xnor2_1 _18597_ (.A(_06957_),
    .B(_06958_),
    .Y(_00758_));
 sky130_fd_sc_hd__or2_4 _18598_ (.A(net524),
    .B(\hash.CA2.b_dash[18] ),
    .X(_12951_));
 sky130_fd_sc_hd__nand2_1 _18599_ (.A(_12930_),
    .B(_06957_),
    .Y(_06959_));
 sky130_fd_sc_hd__nor4_1 _18600_ (.A(\hash.CA2.b_dash[14] ),
    .B(\hash.CA2.b_dash[16] ),
    .C(_06952_),
    .D(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__xor2_1 _18601_ (.A(_12951_),
    .B(_06960_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_4 _18602_ (.A(net524),
    .B(\hash.CA2.b_dash[19] ),
    .X(_12957_));
 sky130_fd_sc_hd__or3_1 _18603_ (.A(net524),
    .B(\hash.CA2.b_dash[16] ),
    .C(\hash.CA2.b_dash[18] ),
    .X(_06961_));
 sky130_fd_sc_hd__nor3_1 _18604_ (.A(_06954_),
    .B(_06959_),
    .C(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__xor2_1 _18605_ (.A(_12957_),
    .B(_06962_),
    .X(_00760_));
 sky130_fd_sc_hd__nor3_2 _18606_ (.A(\hash.CA2.b_dash[17] ),
    .B(_12957_),
    .C(_06961_),
    .Y(_06963_));
 sky130_fd_sc_hd__nand4_4 _18607_ (.A(_06946_),
    .B(_06949_),
    .C(_06955_),
    .D(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__nand2_2 _18608_ (.A(_06210_),
    .B(\hash.CA2.b_dash[20] ),
    .Y(_12964_));
 sky130_fd_sc_hd__xnor2_2 _18609_ (.A(_06964_),
    .B(_12964_),
    .Y(_00761_));
 sky130_fd_sc_hd__nor2b_2 _18610_ (.A(net521),
    .B_N(\hash.CA2.b_dash[21] ),
    .Y(_12973_));
 sky130_fd_sc_hd__o41a_2 _18611_ (.A1(\hash.CA2.b_dash[19] ),
    .A2(_06954_),
    .A3(_06959_),
    .A4(_06961_),
    .B1(\hash.CA2.b_dash[20] ),
    .X(_06965_));
 sky130_fd_sc_hd__xnor2_1 _18612_ (.A(\hash.CA2.b_dash[21] ),
    .B(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__nor2_1 _18613_ (.A(net521),
    .B(_06966_),
    .Y(_00762_));
 sky130_fd_sc_hd__nor2_2 _18614_ (.A(net521),
    .B(\hash.CA2.b_dash[22] ),
    .Y(_12981_));
 sky130_fd_sc_hd__and4_1 _18615_ (.A(_06210_),
    .B(\hash.CA2.b_dash[20] ),
    .C(\hash.CA2.b_dash[21] ),
    .D(_06964_),
    .X(_06967_));
 sky130_fd_sc_hd__xor2_1 _18616_ (.A(_12981_),
    .B(_06967_),
    .X(_00763_));
 sky130_fd_sc_hd__nor2b_4 _18617_ (.A(net521),
    .B_N(\hash.CA2.b_dash[23] ),
    .Y(_12989_));
 sky130_fd_sc_hd__a211o_1 _18618_ (.A1(\hash.CA2.b_dash[21] ),
    .A2(_06965_),
    .B1(\hash.CA2.b_dash[22] ),
    .C1(net521),
    .X(_06968_));
 sky130_fd_sc_hd__xor2_1 _18619_ (.A(_12989_),
    .B(_06968_),
    .X(_00764_));
 sky130_fd_sc_hd__nor2_2 _18620_ (.A(net521),
    .B(\hash.CA2.b_dash[24] ),
    .Y(_12997_));
 sky130_fd_sc_hd__or2_0 _18621_ (.A(\hash.CA2.b_dash[22] ),
    .B(_06967_),
    .X(_06969_));
 sky130_fd_sc_hd__nand2_1 _18622_ (.A(_12989_),
    .B(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__xnor2_1 _18623_ (.A(_12997_),
    .B(_06970_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand2_1 _18624_ (.A(_06210_),
    .B(\hash.CA2.b_dash[25] ),
    .Y(_06971_));
 sky130_fd_sc_hd__clkinvlp_4 _18625_ (.A(_06971_),
    .Y(_13005_));
 sky130_fd_sc_hd__a21boi_0 _18626_ (.A1(_12989_),
    .A2(_06968_),
    .B1_N(_12997_),
    .Y(_06972_));
 sky130_fd_sc_hd__xnor2_1 _18627_ (.A(_13005_),
    .B(_06972_),
    .Y(_00766_));
 sky130_fd_sc_hd__a21oi_1 _18628_ (.A1(\hash.CA2.b_dash[23] ),
    .A2(_06969_),
    .B1(\hash.CA2.b_dash[24] ),
    .Y(_06973_));
 sky130_fd_sc_hd__nor2_1 _18629_ (.A(net521),
    .B(\hash.CA2.b_dash[26] ),
    .Y(_06974_));
 sky130_fd_sc_hd__o21ai_1 _18630_ (.A1(_06971_),
    .A2(_06973_),
    .B1(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__nor2_1 _18631_ (.A(_06971_),
    .B(_06973_),
    .Y(_06976_));
 sky130_fd_sc_hd__inv_1 _18632_ (.A(_06974_),
    .Y(_13013_));
 sky130_fd_sc_hd__nand2_1 _18633_ (.A(_06976_),
    .B(_13013_),
    .Y(_06977_));
 sky130_fd_sc_hd__nand2_1 _18634_ (.A(_06975_),
    .B(_06977_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2b_2 _18635_ (.A(net521),
    .B_N(\hash.CA2.b_dash[27] ),
    .Y(_13020_));
 sky130_fd_sc_hd__inv_1 _18636_ (.A(\hash.CA2.b_dash[25] ),
    .Y(_06978_));
 sky130_fd_sc_hd__a21oi_1 _18637_ (.A1(\hash.CA2.b_dash[23] ),
    .A2(_06968_),
    .B1(\hash.CA2.b_dash[24] ),
    .Y(_06979_));
 sky130_fd_sc_hd__o21ai_1 _18638_ (.A1(_06978_),
    .A2(_06979_),
    .B1(_06974_),
    .Y(_06980_));
 sky130_fd_sc_hd__xor2_1 _18639_ (.A(_13020_),
    .B(_06980_),
    .X(_00768_));
 sky130_fd_sc_hd__nor2b_1 _18640_ (.A(net523),
    .B_N(\hash.CA2.b_dash[28] ),
    .Y(_13028_));
 sky130_fd_sc_hd__o21ai_0 _18641_ (.A1(\hash.CA2.b_dash[26] ),
    .A2(_06976_),
    .B1(\hash.CA2.b_dash[27] ),
    .Y(_06981_));
 sky130_fd_sc_hd__xor2_1 _18642_ (.A(\hash.CA2.b_dash[28] ),
    .B(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__nor2_1 _18643_ (.A(net521),
    .B(_06982_),
    .Y(_00769_));
 sky130_fd_sc_hd__or2_2 _18644_ (.A(net521),
    .B(\hash.CA2.b_dash[29] ),
    .X(_13035_));
 sky130_fd_sc_hd__and3_1 _18645_ (.A(\hash.CA2.b_dash[28] ),
    .B(_13020_),
    .C(_06980_),
    .X(_06983_));
 sky130_fd_sc_hd__xnor2_1 _18646_ (.A(_13035_),
    .B(_06983_),
    .Y(_00770_));
 sky130_fd_sc_hd__nor2b_2 _18647_ (.A(net521),
    .B_N(\hash.CA2.b_dash[30] ),
    .Y(_13042_));
 sky130_fd_sc_hd__a31oi_1 _18648_ (.A1(\hash.CA2.b_dash[28] ),
    .A2(_06975_),
    .A3(_13020_),
    .B1(_13035_),
    .Y(_06984_));
 sky130_fd_sc_hd__xnor2_1 _18649_ (.A(_13042_),
    .B(_06984_),
    .Y(_00771_));
 sky130_fd_sc_hd__o21ai_1 _18650_ (.A1(\hash.CA2.b_dash[29] ),
    .A2(_06983_),
    .B1(\hash.CA2.b_dash[30] ),
    .Y(_06985_));
 sky130_fd_sc_hd__xnor2_1 _18651_ (.A(\hash.CA2.b_dash[31] ),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__nor2_1 _18652_ (.A(net521),
    .B(_06986_),
    .Y(_00773_));
 sky130_fd_sc_hd__xor2_1 _18653_ (.A(_14027_),
    .B(_13847_),
    .X(_00742_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1126 ();
 sky130_fd_sc_hd__nand3_1 _18655_ (.A(\hash.CA2.a_dash[1] ),
    .B(\hash.CA2.a_dash[2] ),
    .C(\hash.CA2.a_dash[3] ),
    .Y(_06988_));
 sky130_fd_sc_hd__xnor2_1 _18656_ (.A(\hash.CA2.a_dash[4] ),
    .B(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__nor2_1 _18657_ (.A(net520),
    .B(_06989_),
    .Y(_00744_));
 sky130_fd_sc_hd__or2_0 _18658_ (.A(net520),
    .B(\hash.CA2.a_dash[4] ),
    .X(_13853_));
 sky130_fd_sc_hd__a21oi_1 _18659_ (.A1(\hash.CA2.a_dash[3] ),
    .A2(_14027_),
    .B1(\hash.CA2.a_dash[4] ),
    .Y(_06990_));
 sky130_fd_sc_hd__xnor2_1 _18660_ (.A(\hash.CA2.a_dash[5] ),
    .B(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand2_1 _18661_ (.A(net519),
    .B(_06991_),
    .Y(_00745_));
 sky130_fd_sc_hd__nor3_1 _18662_ (.A(net520),
    .B(\hash.CA2.a_dash[4] ),
    .C(\hash.CA2.a_dash[5] ),
    .Y(_06992_));
 sky130_fd_sc_hd__nand2_1 _18663_ (.A(_06988_),
    .B(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__xnor2_1 _18664_ (.A(_13865_),
    .B(_06993_),
    .Y(_00746_));
 sky130_fd_sc_hd__a21oi_1 _18665_ (.A1(\hash.CA2.a_dash[3] ),
    .A2(_14027_),
    .B1(\hash.CA2.a_dash[6] ),
    .Y(_06994_));
 sky130_fd_sc_hd__nand2_1 _18666_ (.A(_06992_),
    .B(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__nand2_1 _18667_ (.A(net519),
    .B(\hash.CA2.a_dash[7] ),
    .Y(_06996_));
 sky130_fd_sc_hd__xnor2_1 _18668_ (.A(_06995_),
    .B(_06996_),
    .Y(_00747_));
 sky130_fd_sc_hd__or2_1 _18669_ (.A(net520),
    .B(\hash.CA2.a_dash[8] ),
    .X(_13878_));
 sky130_fd_sc_hd__o21ai_0 _18670_ (.A1(\hash.CA2.a_dash[6] ),
    .A2(_06993_),
    .B1(\hash.CA2.a_dash[7] ),
    .Y(_06997_));
 sky130_fd_sc_hd__xnor2_1 _18671_ (.A(\hash.CA2.a_dash[8] ),
    .B(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__nor2_1 _18672_ (.A(net520),
    .B(_06998_),
    .Y(_00748_));
 sky130_fd_sc_hd__a21oi_2 _18673_ (.A1(\hash.CA2.a_dash[7] ),
    .A2(_06995_),
    .B1(\hash.CA2.a_dash[8] ),
    .Y(_06999_));
 sky130_fd_sc_hd__xnor2_1 _18674_ (.A(\hash.CA2.a_dash[9] ),
    .B(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand2_1 _18675_ (.A(net519),
    .B(_07000_),
    .Y(_00749_));
 sky130_fd_sc_hd__nor2b_2 _18676_ (.A(net520),
    .B_N(\hash.CA2.a_dash[10] ),
    .Y(_13889_));
 sky130_fd_sc_hd__nor2_1 _18677_ (.A(\hash.CA2.a_dash[6] ),
    .B(_06993_),
    .Y(_07001_));
 sky130_fd_sc_hd__nor2_1 _18678_ (.A(\hash.CA2.a_dash[9] ),
    .B(_13878_),
    .Y(_07002_));
 sky130_fd_sc_hd__o21ai_1 _18679_ (.A1(_06996_),
    .A2(_07001_),
    .B1(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__xor2_1 _18680_ (.A(_13889_),
    .B(_07003_),
    .X(_00750_));
 sky130_fd_sc_hd__nor2_2 _18681_ (.A(net520),
    .B(_04827_),
    .Y(_13895_));
 sky130_fd_sc_hd__nand2_1 _18682_ (.A(_06475_),
    .B(_06999_),
    .Y(_07004_));
 sky130_fd_sc_hd__nand2_1 _18683_ (.A(_13889_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__xnor2_1 _18684_ (.A(_13895_),
    .B(_07005_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand2_2 _18685_ (.A(net519),
    .B(_04833_),
    .Y(_13902_));
 sky130_fd_sc_hd__nand2_1 _18686_ (.A(\hash.CA2.a_dash[11] ),
    .B(_13889_),
    .Y(_07006_));
 sky130_fd_sc_hd__nor2b_1 _18687_ (.A(_07006_),
    .B_N(_07003_),
    .Y(_07007_));
 sky130_fd_sc_hd__xnor2_1 _18688_ (.A(_13902_),
    .B(_07007_),
    .Y(_00723_));
 sky130_fd_sc_hd__a21oi_2 _18689_ (.A1(_06475_),
    .A2(_06999_),
    .B1(_07006_),
    .Y(_07008_));
 sky130_fd_sc_hd__or3_1 _18690_ (.A(\hash.CA2.a_dash[12] ),
    .B(\hash.CA2.a_dash[13] ),
    .C(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__o21ai_0 _18691_ (.A1(\hash.CA2.a_dash[12] ),
    .A2(_07008_),
    .B1(\hash.CA2.a_dash[13] ),
    .Y(_07010_));
 sky130_fd_sc_hd__nand3_1 _18692_ (.A(net519),
    .B(_07009_),
    .C(_07010_),
    .Y(_00724_));
 sky130_fd_sc_hd__nor3_1 _18693_ (.A(\hash.CA2.a_dash[13] ),
    .B(_13902_),
    .C(_07007_),
    .Y(_07011_));
 sky130_fd_sc_hd__xnor2_1 _18694_ (.A(_06476_),
    .B(_07011_),
    .Y(_00725_));
 sky130_fd_sc_hd__or4_2 _18695_ (.A(\hash.CA2.a_dash[13] ),
    .B(_13914_),
    .C(_13902_),
    .D(_07008_),
    .X(_07012_));
 sky130_fd_sc_hd__xnor2_1 _18696_ (.A(_13921_),
    .B(_07012_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand2_2 _18697_ (.A(net519),
    .B(\hash.CA2.a_dash[16] ),
    .Y(_07013_));
 sky130_fd_sc_hd__nor2_1 _18698_ (.A(\hash.CA2.a_dash[14] ),
    .B(_13921_),
    .Y(_07014_));
 sky130_fd_sc_hd__nand2_1 _18699_ (.A(_07011_),
    .B(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__xnor2_1 _18700_ (.A(_07013_),
    .B(_07015_),
    .Y(_00727_));
 sky130_fd_sc_hd__or2_0 _18701_ (.A(net523),
    .B(\hash.CA2.a_dash[17] ),
    .X(_13935_));
 sky130_fd_sc_hd__o21ai_0 _18702_ (.A1(\hash.CA2.a_dash[15] ),
    .A2(_07012_),
    .B1(\hash.CA2.a_dash[16] ),
    .Y(_07016_));
 sky130_fd_sc_hd__xnor2_1 _18703_ (.A(\hash.CA2.a_dash[17] ),
    .B(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__nor2_1 _18704_ (.A(net524),
    .B(_07017_),
    .Y(_00728_));
 sky130_fd_sc_hd__or2_2 _18705_ (.A(net524),
    .B(\hash.CA2.a_dash[18] ),
    .X(_13941_));
 sky130_fd_sc_hd__a21o_1 _18706_ (.A1(\hash.CA2.a_dash[16] ),
    .A2(_07015_),
    .B1(\hash.CA2.a_dash[17] ),
    .X(_07018_));
 sky130_fd_sc_hd__xor2_1 _18707_ (.A(\hash.CA2.a_dash[18] ),
    .B(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__nand2_1 _18708_ (.A(net519),
    .B(_07019_),
    .Y(_00729_));
 sky130_fd_sc_hd__nor2_1 _18709_ (.A(\hash.CA2.a_dash[15] ),
    .B(_07012_),
    .Y(_07020_));
 sky130_fd_sc_hd__nor2_1 _18710_ (.A(\hash.CA2.a_dash[17] ),
    .B(_13941_),
    .Y(_07021_));
 sky130_fd_sc_hd__o21ai_2 _18711_ (.A1(_07013_),
    .A2(_07020_),
    .B1(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__xnor2_2 _18712_ (.A(_13946_),
    .B(_07022_),
    .Y(_00730_));
 sky130_fd_sc_hd__nor3_1 _18713_ (.A(\hash.CA2.a_dash[18] ),
    .B(\hash.CA2.a_dash[19] ),
    .C(_07018_),
    .Y(_07023_));
 sky130_fd_sc_hd__xnor2_2 _18714_ (.A(_04898_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__nand2_1 _18715_ (.A(net519),
    .B(_07024_),
    .Y(_00731_));
 sky130_fd_sc_hd__or2_0 _18716_ (.A(net521),
    .B(\hash.CA2.a_dash[21] ),
    .X(_13956_));
 sky130_fd_sc_hd__or2_1 _18717_ (.A(\hash.CA2.a_dash[19] ),
    .B(_07022_),
    .X(_07025_));
 sky130_fd_sc_hd__nand2_1 _18718_ (.A(\hash.CA2.a_dash[20] ),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__xnor2_2 _18719_ (.A(\hash.CA2.a_dash[21] ),
    .B(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__nor2_1 _18720_ (.A(net521),
    .B(_07027_),
    .Y(_00732_));
 sky130_fd_sc_hd__or2_2 _18721_ (.A(net521),
    .B(\hash.CA2.a_dash[22] ),
    .X(_13961_));
 sky130_fd_sc_hd__o31ai_1 _18722_ (.A1(\hash.CA2.a_dash[19] ),
    .A2(_13941_),
    .A3(_07018_),
    .B1(\hash.CA2.a_dash[20] ),
    .Y(_07028_));
 sky130_fd_sc_hd__nand2b_2 _18723_ (.A_N(\hash.CA2.a_dash[21] ),
    .B(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__xor2_1 _18724_ (.A(\hash.CA2.a_dash[22] ),
    .B(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__nand2_1 _18725_ (.A(net519),
    .B(_07030_),
    .Y(_00733_));
 sky130_fd_sc_hd__nor2b_2 _18726_ (.A(net521),
    .B_N(\hash.CA2.a_dash[23] ),
    .Y(_13967_));
 sky130_fd_sc_hd__nor2_1 _18727_ (.A(net521),
    .B(_04898_),
    .Y(_13951_));
 sky130_fd_sc_hd__a211oi_4 _18728_ (.A1(_07025_),
    .A2(_13951_),
    .B1(_13961_),
    .C1(\hash.CA2.a_dash[21] ),
    .Y(_07031_));
 sky130_fd_sc_hd__xnor2_1 _18729_ (.A(_13967_),
    .B(_07031_),
    .Y(_00734_));
 sky130_fd_sc_hd__o21ai_0 _18730_ (.A1(\hash.CA2.a_dash[22] ),
    .A2(_07029_),
    .B1(\hash.CA2.a_dash[23] ),
    .Y(_07032_));
 sky130_fd_sc_hd__xor2_1 _18731_ (.A(\hash.CA2.a_dash[24] ),
    .B(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__nor2_1 _18732_ (.A(net524),
    .B(_07033_),
    .Y(_00735_));
 sky130_fd_sc_hd__nor2b_1 _18733_ (.A(net521),
    .B_N(\hash.CA2.a_dash[25] ),
    .Y(_13981_));
 sky130_fd_sc_hd__nand2_1 _18734_ (.A(\hash.CA2.a_dash[24] ),
    .B(_13967_),
    .Y(_07034_));
 sky130_fd_sc_hd__nor2_1 _18735_ (.A(_07031_),
    .B(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__xor2_1 _18736_ (.A(_13981_),
    .B(_07035_),
    .X(_00736_));
 sky130_fd_sc_hd__nand3_1 _18737_ (.A(\hash.CA2.a_dash[24] ),
    .B(_13967_),
    .C(_13981_),
    .Y(_07036_));
 sky130_fd_sc_hd__o21ba_1 _18738_ (.A1(_13961_),
    .A2(_07029_),
    .B1_N(_07036_),
    .X(_07037_));
 sky130_fd_sc_hd__xnor2_1 _18739_ (.A(_06480_),
    .B(_07037_),
    .Y(_00737_));
 sky130_fd_sc_hd__nor2_2 _18740_ (.A(_07031_),
    .B(_07036_),
    .Y(_07038_));
 sky130_fd_sc_hd__or3_1 _18741_ (.A(\hash.CA2.a_dash[26] ),
    .B(\hash.CA2.a_dash[27] ),
    .C(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__o21ai_0 _18742_ (.A1(\hash.CA2.a_dash[26] ),
    .A2(_07038_),
    .B1(\hash.CA2.a_dash[27] ),
    .Y(_07040_));
 sky130_fd_sc_hd__nand3_1 _18743_ (.A(net519),
    .B(_07039_),
    .C(_07040_),
    .Y(_00738_));
 sky130_fd_sc_hd__nor3_1 _18744_ (.A(\hash.CA2.a_dash[27] ),
    .B(_06480_),
    .C(_07037_),
    .Y(_07041_));
 sky130_fd_sc_hd__xor2_1 _18745_ (.A(_14002_),
    .B(_07041_),
    .X(_00739_));
 sky130_fd_sc_hd__or3_1 _18746_ (.A(\hash.CA2.a_dash[27] ),
    .B(\hash.CA2.a_dash[28] ),
    .C(_06480_),
    .X(_07042_));
 sky130_fd_sc_hd__nor2_1 _18747_ (.A(_07038_),
    .B(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__xor2_1 _18748_ (.A(_14008_),
    .B(_07043_),
    .X(_00740_));
 sky130_fd_sc_hd__nor2_1 _18749_ (.A(net521),
    .B(_04976_),
    .Y(_14013_));
 sky130_fd_sc_hd__nor3_1 _18750_ (.A(\hash.CA2.a_dash[29] ),
    .B(_07037_),
    .C(_07042_),
    .Y(_07044_));
 sky130_fd_sc_hd__xnor2_1 _18751_ (.A(_14013_),
    .B(_07044_),
    .Y(_00741_));
 sky130_fd_sc_hd__o31ai_1 _18752_ (.A1(\hash.CA2.a_dash[29] ),
    .A2(_07038_),
    .A3(_07042_),
    .B1(\hash.CA2.a_dash[30] ),
    .Y(_07045_));
 sky130_fd_sc_hd__xor2_1 _18753_ (.A(\hash.CA2.a_dash[31] ),
    .B(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__nor2_1 _18754_ (.A(net521),
    .B(_07046_),
    .Y(_00743_));
 sky130_fd_sc_hd__xnor2_1 _18755_ (.A(_14028_),
    .B(\hash.CA1.b[2] ),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(_13090_),
    .B(_12253_),
    .Y(_07047_));
 sky130_fd_sc_hd__nand2_2 _18757_ (.A(_04840_),
    .B(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__xor2_1 _18758_ (.A(_04646_),
    .B(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__nand2_1 _18759_ (.A(net519),
    .B(_07049_),
    .Y(_00714_));
 sky130_fd_sc_hd__nor2_2 _18760_ (.A(_14028_),
    .B(_04592_),
    .Y(_07050_));
 sky130_fd_sc_hd__o21ai_0 _18761_ (.A1(_04646_),
    .A2(_07050_),
    .B1(_04654_),
    .Y(_07051_));
 sky130_fd_sc_hd__or3_1 _18762_ (.A(_04646_),
    .B(_04654_),
    .C(_07050_),
    .X(_07052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1125 ();
 sky130_fd_sc_hd__a21oi_1 _18764_ (.A1(_07051_),
    .A2(_07052_),
    .B1(net520),
    .Y(_00715_));
 sky130_fd_sc_hd__nor3b_1 _18765_ (.A(net520),
    .B(_04646_),
    .C_N(_04654_),
    .Y(_07054_));
 sky130_fd_sc_hd__nand2_1 _18766_ (.A(_07048_),
    .B(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__xnor2_1 _18767_ (.A(\hash.CA1.b[5] ),
    .B(_07055_),
    .Y(_00716_));
 sky130_fd_sc_hd__and2_0 _18768_ (.A(_04674_),
    .B(_07054_),
    .X(_07056_));
 sky130_fd_sc_hd__nor2b_1 _18769_ (.A(_07050_),
    .B_N(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__xor2_1 _18770_ (.A(\hash.CA1.b[6] ),
    .B(_07057_),
    .X(_00717_));
 sky130_fd_sc_hd__nand3_2 _18771_ (.A(\hash.CA1.b[6] ),
    .B(_07048_),
    .C(_07056_),
    .Y(_07058_));
 sky130_fd_sc_hd__xor2_1 _18772_ (.A(\hash.CA1.b[7] ),
    .B(_07058_),
    .X(_00718_));
 sky130_fd_sc_hd__and4b_1 _18773_ (.A_N(_07050_),
    .B(_07054_),
    .C(_04674_),
    .D(_04701_),
    .X(_07059_));
 sky130_fd_sc_hd__nor3_1 _18774_ (.A(_04724_),
    .B(_04742_),
    .C(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__o21ai_4 _18775_ (.A1(_04724_),
    .A2(_07059_),
    .B1(_04742_),
    .Y(_07061_));
 sky130_fd_sc_hd__nand2b_1 _18776_ (.A_N(_07060_),
    .B(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__nand2_1 _18777_ (.A(net519),
    .B(_07062_),
    .Y(_00719_));
 sky130_fd_sc_hd__a21boi_4 _18778_ (.A1(_06474_),
    .A2(_07058_),
    .B1_N(\hash.CA1.b[8] ),
    .Y(_07063_));
 sky130_fd_sc_hd__nand2_1 _18779_ (.A(_04773_),
    .B(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__o21ai_0 _18780_ (.A1(\hash.CA1.b[9] ),
    .A2(_07063_),
    .B1(_07064_),
    .Y(_00720_));
 sky130_fd_sc_hd__and3_1 _18781_ (.A(_04895_),
    .B(_04791_),
    .C(_07061_),
    .X(_07065_));
 sky130_fd_sc_hd__a21oi_1 _18782_ (.A1(_04895_),
    .A2(_07061_),
    .B1(_04791_),
    .Y(_07066_));
 sky130_fd_sc_hd__o21ai_0 _18783_ (.A1(_07065_),
    .A2(_07066_),
    .B1(net519),
    .Y(_00691_));
 sky130_fd_sc_hd__nor3_1 _18784_ (.A(_04791_),
    .B(\hash.CA1.b[9] ),
    .C(_07063_),
    .Y(_07067_));
 sky130_fd_sc_hd__xor2_1 _18785_ (.A(\hash.CA1.b[11] ),
    .B(_07067_),
    .X(_00692_));
 sky130_fd_sc_hd__o2111a_1 _18786_ (.A1(_04788_),
    .A2(_04790_),
    .B1(_04813_),
    .C1(_04895_),
    .D1(_06210_),
    .X(_07068_));
 sky130_fd_sc_hd__nand2_1 _18787_ (.A(_07061_),
    .B(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__xor2_1 _18788_ (.A(\hash.CA1.b[12] ),
    .B(_07069_),
    .X(_00693_));
 sky130_fd_sc_hd__a21oi_1 _18789_ (.A1(_04813_),
    .A2(_07067_),
    .B1(net1162),
    .Y(_07070_));
 sky130_fd_sc_hd__xnor2_1 _18790_ (.A(_04611_),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__nor2_1 _18791_ (.A(net520),
    .B(_07071_),
    .Y(_00694_));
 sky130_fd_sc_hd__a21oi_2 _18792_ (.A1(_07061_),
    .A2(_07068_),
    .B1(net1162),
    .Y(_07072_));
 sky130_fd_sc_hd__o21a_1 _18793_ (.A1(_04842_),
    .A2(_07072_),
    .B1(_04627_),
    .X(_07073_));
 sky130_fd_sc_hd__nor3_1 _18794_ (.A(_04842_),
    .B(_04627_),
    .C(_07072_),
    .Y(_07074_));
 sky130_fd_sc_hd__o21ai_0 _18795_ (.A1(_07073_),
    .A2(_07074_),
    .B1(net519),
    .Y(_00695_));
 sky130_fd_sc_hd__nand4b_2 _18796_ (.A_N(_04791_),
    .B(_04611_),
    .C(_04895_),
    .D(_04813_),
    .Y(_07075_));
 sky130_fd_sc_hd__o221ai_2 _18797_ (.A1(_04842_),
    .A2(\hash.CA1.b[12] ),
    .B1(_07063_),
    .B2(_07075_),
    .C1(\hash.CA1.b[14] ),
    .Y(_07076_));
 sky130_fd_sc_hd__xor2_1 _18798_ (.A(\hash.CA1.b[15] ),
    .B(_07076_),
    .X(_00696_));
 sky130_fd_sc_hd__nand2_1 _18799_ (.A(\hash.CA1.b[12] ),
    .B(_07069_),
    .Y(_07077_));
 sky130_fd_sc_hd__nand2_1 _18800_ (.A(_04611_),
    .B(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__a21oi_1 _18801_ (.A1(_04627_),
    .A2(_07078_),
    .B1(_04659_),
    .Y(_07079_));
 sky130_fd_sc_hd__xor2_1 _18802_ (.A(net1129),
    .B(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__nand2_1 _18803_ (.A(net519),
    .B(_07080_),
    .Y(_00697_));
 sky130_fd_sc_hd__o221ai_4 _18804_ (.A1(_04842_),
    .A2(\hash.CA1.b[12] ),
    .B1(_07063_),
    .B2(_07075_),
    .C1(_04627_),
    .Y(_07081_));
 sky130_fd_sc_hd__and3b_1 _18805_ (.A_N(\hash.CA1.b[15] ),
    .B(_07081_),
    .C(net1130),
    .X(_07082_));
 sky130_fd_sc_hd__xnor2_1 _18806_ (.A(_06477_),
    .B(_07082_),
    .Y(_00698_));
 sky130_fd_sc_hd__o21ai_4 _18807_ (.A1(\hash.CA1.b[13] ),
    .A2(_07072_),
    .B1(_04627_),
    .Y(_07083_));
 sky130_fd_sc_hd__nand4b_1 _18808_ (.A_N(\hash.CA1.b[15] ),
    .B(_06477_),
    .C(_07083_),
    .D(net1132),
    .Y(_07084_));
 sky130_fd_sc_hd__xnor2_1 _18809_ (.A(\hash.CA1.b[18] ),
    .B(_07084_),
    .Y(_00699_));
 sky130_fd_sc_hd__nor4b_2 _18810_ (.A(_04699_),
    .B(\hash.CA1.b[15] ),
    .C(_04721_),
    .D_N(net1130),
    .Y(_07085_));
 sky130_fd_sc_hd__nand2_1 _18811_ (.A(_07081_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__xor2_1 _18812_ (.A(\hash.CA1.b[19] ),
    .B(_07086_),
    .X(_00700_));
 sky130_fd_sc_hd__a21oi_1 _18813_ (.A1(_07083_),
    .A2(_07085_),
    .B1(_04740_),
    .Y(_07087_));
 sky130_fd_sc_hd__xor2_1 _18814_ (.A(net1142),
    .B(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__nor2_1 _18815_ (.A(net524),
    .B(_07088_),
    .Y(_00701_));
 sky130_fd_sc_hd__or3_1 _18816_ (.A(net524),
    .B(_04740_),
    .C(net1141),
    .X(_07089_));
 sky130_fd_sc_hd__a21oi_2 _18817_ (.A1(_07081_),
    .A2(_07085_),
    .B1(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__xnor2_1 _18818_ (.A(_06478_),
    .B(_07090_),
    .Y(_00702_));
 sky130_fd_sc_hd__a21oi_2 _18819_ (.A1(_07083_),
    .A2(_07085_),
    .B1(_07089_),
    .Y(_07091_));
 sky130_fd_sc_hd__nor2_1 _18820_ (.A(_06478_),
    .B(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__nor2_1 _18821_ (.A(\hash.CA1.b[22] ),
    .B(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__a21oi_1 _18822_ (.A1(net1123),
    .A2(_07092_),
    .B1(_07093_),
    .Y(_00703_));
 sky130_fd_sc_hd__or2_0 _18823_ (.A(net1122),
    .B(_06478_),
    .X(_07094_));
 sky130_fd_sc_hd__or2_2 _18824_ (.A(_07090_),
    .B(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__xor2_1 _18825_ (.A(_06479_),
    .B(_07095_),
    .X(_00704_));
 sky130_fd_sc_hd__o21ai_0 _18826_ (.A1(_07091_),
    .A2(_07094_),
    .B1(net1169),
    .Y(_07096_));
 sky130_fd_sc_hd__xnor2_1 _18827_ (.A(net1134),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__nor2_1 _18828_ (.A(net524),
    .B(_07097_),
    .Y(_00705_));
 sky130_fd_sc_hd__a21oi_1 _18829_ (.A1(net1169),
    .A2(_07095_),
    .B1(net1134),
    .Y(_07098_));
 sky130_fd_sc_hd__xnor2_1 _18830_ (.A(net1164),
    .B(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__nand2_1 _18831_ (.A(net519),
    .B(_07099_),
    .Y(_00706_));
 sky130_fd_sc_hd__o21ai_1 _18832_ (.A1(_07091_),
    .A2(_07094_),
    .B1(_06479_),
    .Y(_07100_));
 sky130_fd_sc_hd__nor3_1 _18833_ (.A(net521),
    .B(net1133),
    .C(net1164),
    .Y(_07101_));
 sky130_fd_sc_hd__nand2_1 _18834_ (.A(_07100_),
    .B(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__xor2_1 _18835_ (.A(\hash.CA1.b[26] ),
    .B(_07102_),
    .X(_00707_));
 sky130_fd_sc_hd__a211o_1 _18836_ (.A1(_06479_),
    .A2(_07095_),
    .B1(net1133),
    .C1(net1164),
    .X(_07103_));
 sky130_fd_sc_hd__nand2_1 _18837_ (.A(\hash.CA1.b[26] ),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__xor2_1 _18838_ (.A(_06481_),
    .B(_07104_),
    .X(_00708_));
 sky130_fd_sc_hd__a21oi_1 _18839_ (.A1(\hash.CA1.b[26] ),
    .A2(_07102_),
    .B1(_06481_),
    .Y(_07105_));
 sky130_fd_sc_hd__xor2_1 _18840_ (.A(\hash.CA1.b[28] ),
    .B(_07105_),
    .X(_00709_));
 sky130_fd_sc_hd__or2_1 _18841_ (.A(net521),
    .B(_04756_),
    .X(\hash.CA1.b[29] ));
 sky130_fd_sc_hd__or2_0 _18842_ (.A(_04736_),
    .B(_06481_),
    .X(_07106_));
 sky130_fd_sc_hd__a21oi_1 _18843_ (.A1(\hash.CA1.b[26] ),
    .A2(_07103_),
    .B1(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__xor2_1 _18844_ (.A(\hash.CA1.b[29] ),
    .B(_07107_),
    .X(_00710_));
 sky130_fd_sc_hd__a2111oi_1 _18845_ (.A1(_04694_),
    .A2(_07102_),
    .B1(_06481_),
    .C1(_04756_),
    .D1(_04736_),
    .Y(_07108_));
 sky130_fd_sc_hd__xnor2_1 _18846_ (.A(\hash.CA1.b[30] ),
    .B(_07108_),
    .Y(_00712_));
 sky130_fd_sc_hd__nand2_1 _18847_ (.A(net519),
    .B(_04805_),
    .Y(_07109_));
 sky130_fd_sc_hd__nor2_1 _18848_ (.A(_04756_),
    .B(_07106_),
    .Y(_07110_));
 sky130_fd_sc_hd__o21ai_0 _18849_ (.A1(_04652_),
    .A2(net1165),
    .B1(\hash.CA1.b[26] ),
    .Y(_07111_));
 sky130_fd_sc_hd__nand3_1 _18850_ (.A(_06479_),
    .B(\hash.CA1.b[26] ),
    .C(_07095_),
    .Y(_07112_));
 sky130_fd_sc_hd__a31oi_2 _18851_ (.A1(_07110_),
    .A2(_07111_),
    .A3(_07112_),
    .B1(net1118),
    .Y(_07113_));
 sky130_fd_sc_hd__mux2i_1 _18852_ (.A0(\hash.CA1.b[31] ),
    .A1(_07109_),
    .S(_07113_),
    .Y(_00713_));
 sky130_fd_sc_hd__xnor2_1 _18853_ (.A(\hash.CA1.S1.X[6] ),
    .B(\hash.CA1.S1.X[11] ),
    .Y(_07114_));
 sky130_fd_sc_hd__xnor2_4 _18854_ (.A(_07114_),
    .B(\hash.CA1.S1.X[25] ),
    .Y(_14030_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1124 ();
 sky130_fd_sc_hd__nor2b_1 _18856_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[0] ),
    .Y(\hash.CA1.f[0] ));
 sky130_fd_sc_hd__xnor2_1 _18857_ (.A(_06722_),
    .B(\hash.CA1.S1.X[12] ),
    .Y(_07116_));
 sky130_fd_sc_hd__xnor2_2 _18858_ (.A(_06886_),
    .B(_07116_),
    .Y(_14035_));
 sky130_fd_sc_hd__inv_1 _18859_ (.A(_14035_),
    .Y(_12673_));
 sky130_fd_sc_hd__nor2b_1 _18860_ (.A(\hash.reset ),
    .B_N(\hash.CA2.S1.X[1] ),
    .Y(\hash.CA1.f[1] ));
 sky130_fd_sc_hd__mux2i_1 _18861_ (.A0(\hash.CA2.S1.X[1] ),
    .A1(\hash.CA2.e_dash[1] ),
    .S(_12536_),
    .Y(_07117_));
 sky130_fd_sc_hd__nor2_1 _18862_ (.A(\hash.reset ),
    .B(_07117_),
    .Y(_14034_));
 sky130_fd_sc_hd__inv_1 _18863_ (.A(_14034_),
    .Y(_12672_));
 sky130_fd_sc_hd__xor2_1 _18864_ (.A(_12669_),
    .B(_14039_),
    .X(_12680_));
 sky130_fd_sc_hd__inv_1 _18865_ (.A(_12680_),
    .Y(_12836_));
 sky130_fd_sc_hd__xnor2_2 _18866_ (.A(_12674_),
    .B(_14043_),
    .Y(_12679_));
 sky130_fd_sc_hd__inv_1 _18867_ (.A(_12679_),
    .Y(_12842_));
 sky130_fd_sc_hd__a21oi_1 _18868_ (.A1(_12668_),
    .A2(_14033_),
    .B1(_14032_),
    .Y(_07118_));
 sky130_fd_sc_hd__nor2b_1 _18869_ (.A(_07118_),
    .B_N(_14039_),
    .Y(_07119_));
 sky130_fd_sc_hd__nor2_1 _18870_ (.A(_14038_),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__xor2_2 _18871_ (.A(_14047_),
    .B(_07120_),
    .X(_12685_));
 sky130_fd_sc_hd__a21o_1 _18872_ (.A1(_14031_),
    .A2(_14037_),
    .B1(_14036_),
    .X(_07121_));
 sky130_fd_sc_hd__a21oi_1 _18873_ (.A1(_14043_),
    .A2(_07121_),
    .B1(_14042_),
    .Y(_07122_));
 sky130_fd_sc_hd__xor2_2 _18874_ (.A(_14051_),
    .B(_07122_),
    .X(_12684_));
 sky130_fd_sc_hd__inv_1 _18875_ (.A(_14056_),
    .Y(_07123_));
 sky130_fd_sc_hd__a21o_1 _18876_ (.A1(_12669_),
    .A2(_14039_),
    .B1(_14038_),
    .X(_07124_));
 sky130_fd_sc_hd__a21oi_2 _18877_ (.A1(_14047_),
    .A2(_07124_),
    .B1(_14046_),
    .Y(_07125_));
 sky130_fd_sc_hd__xnor2_2 _18878_ (.A(_07123_),
    .B(_07125_),
    .Y(_12690_));
 sky130_fd_sc_hd__inv_1 _18879_ (.A(_14050_),
    .Y(_07126_));
 sky130_fd_sc_hd__nor2b_1 _18880_ (.A(_12674_),
    .B_N(_14043_),
    .Y(_07127_));
 sky130_fd_sc_hd__o21ai_1 _18881_ (.A1(_14042_),
    .A2(_07127_),
    .B1(_14051_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand2_1 _18882_ (.A(_07126_),
    .B(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__xnor2_2 _18883_ (.A(_14060_),
    .B(_07129_),
    .Y(_12689_));
 sky130_fd_sc_hd__a211oi_2 _18884_ (.A1(_14031_),
    .A2(_14037_),
    .B1(_14036_),
    .C1(_14042_),
    .Y(_07130_));
 sky130_fd_sc_hd__o211ai_2 _18885_ (.A1(_14043_),
    .A2(_14042_),
    .B1(_14060_),
    .C1(_14051_),
    .Y(_07131_));
 sky130_fd_sc_hd__a21oi_4 _18886_ (.A1(_14060_),
    .A2(_14050_),
    .B1(_14059_),
    .Y(_07132_));
 sky130_fd_sc_hd__o21ai_4 _18887_ (.A1(_07131_),
    .A2(_07130_),
    .B1(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__xor2_2 _18888_ (.A(_14070_),
    .B(_07133_),
    .X(_12694_));
 sky130_fd_sc_hd__inv_1 _18889_ (.A(_12694_),
    .Y(_12859_));
 sky130_fd_sc_hd__o21bai_1 _18890_ (.A1(_07123_),
    .A2(_07125_),
    .B1_N(_14055_),
    .Y(_07134_));
 sky130_fd_sc_hd__a21oi_2 _18891_ (.A1(_14066_),
    .A2(_07134_),
    .B1(_14065_),
    .Y(_07135_));
 sky130_fd_sc_hd__xnor2_2 _18892_ (.A(_14075_),
    .B(_07135_),
    .Y(_12700_));
 sky130_fd_sc_hd__inv_1 _18893_ (.A(_12700_),
    .Y(_12862_));
 sky130_fd_sc_hd__a21boi_1 _18894_ (.A1(_07128_),
    .A2(_07126_),
    .B1_N(_14060_),
    .Y(_07136_));
 sky130_fd_sc_hd__o21ai_2 _18895_ (.A1(_07136_),
    .A2(_14059_),
    .B1(_14070_),
    .Y(_07137_));
 sky130_fd_sc_hd__nand2b_1 _18896_ (.A_N(_14069_),
    .B(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__xor2_2 _18897_ (.A(_14079_),
    .B(_07138_),
    .X(_12699_));
 sky130_fd_sc_hd__inv_1 _18898_ (.A(_12699_),
    .Y(_12868_));
 sky130_fd_sc_hd__inv_1 _18899_ (.A(_14065_),
    .Y(_07139_));
 sky130_fd_sc_hd__o21ai_0 _18900_ (.A1(_14056_),
    .A2(_14055_),
    .B1(_14066_),
    .Y(_07140_));
 sky130_fd_sc_hd__nand2_1 _18901_ (.A(_14039_),
    .B(_14047_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand2_1 _18902_ (.A(_14047_),
    .B(_14038_),
    .Y(_07142_));
 sky130_fd_sc_hd__inv_1 _18903_ (.A(_14046_),
    .Y(_07143_));
 sky130_fd_sc_hd__o211ai_2 _18904_ (.A1(_07118_),
    .A2(_07141_),
    .B1(_07142_),
    .C1(_07143_),
    .Y(_07144_));
 sky130_fd_sc_hd__nor3_1 _18905_ (.A(_14055_),
    .B(_14065_),
    .C(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__a21oi_1 _18906_ (.A1(_07139_),
    .A2(_07140_),
    .B1(_07145_),
    .Y(_07146_));
 sky130_fd_sc_hd__a21oi_2 _18907_ (.A1(_14075_),
    .A2(_07146_),
    .B1(_14074_),
    .Y(_07147_));
 sky130_fd_sc_hd__xnor2_4 _18908_ (.A(_14083_),
    .B(_07147_),
    .Y(_12705_));
 sky130_fd_sc_hd__inv_1 _18909_ (.A(_12705_),
    .Y(_12871_));
 sky130_fd_sc_hd__nor3_2 _18910_ (.A(_14070_),
    .B(_14069_),
    .C(_14078_),
    .Y(_07148_));
 sky130_fd_sc_hd__nor2_2 _18911_ (.A(_14079_),
    .B(_14078_),
    .Y(_07149_));
 sky130_fd_sc_hd__nor2_2 _18912_ (.A(_07148_),
    .B(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__o31ai_4 _18913_ (.A1(_14069_),
    .A2(_14078_),
    .A3(_07133_),
    .B1(_07150_),
    .Y(_07151_));
 sky130_fd_sc_hd__xnor2_1 _18914_ (.A(_14087_),
    .B(_07151_),
    .Y(_12704_));
 sky130_fd_sc_hd__inv_1 _18915_ (.A(_12704_),
    .Y(_12876_));
 sky130_fd_sc_hd__nand2_1 _18916_ (.A(_14075_),
    .B(_14083_),
    .Y(_07152_));
 sky130_fd_sc_hd__a21oi_2 _18917_ (.A1(_14083_),
    .A2(_14074_),
    .B1(_14082_),
    .Y(_07153_));
 sky130_fd_sc_hd__o21ai_2 _18918_ (.A1(_07135_),
    .A2(_07152_),
    .B1(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__xnor2_4 _18919_ (.A(_14091_),
    .B(_07154_),
    .Y(_12710_));
 sky130_fd_sc_hd__nor3_2 _18920_ (.A(_14069_),
    .B(_14078_),
    .C(_14086_),
    .Y(_07155_));
 sky130_fd_sc_hd__inv_1 _18921_ (.A(_14087_),
    .Y(_07156_));
 sky130_fd_sc_hd__nor2_1 _18922_ (.A(_07156_),
    .B(_07149_),
    .Y(_07157_));
 sky130_fd_sc_hd__nor2_1 _18923_ (.A(_14086_),
    .B(_07157_),
    .Y(_07158_));
 sky130_fd_sc_hd__a21oi_1 _18924_ (.A1(_07137_),
    .A2(_07155_),
    .B1(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__xnor2_2 _18925_ (.A(_14095_),
    .B(_07159_),
    .Y(_12709_));
 sky130_fd_sc_hd__nand3_1 _18926_ (.A(_14075_),
    .B(_14083_),
    .C(_07146_),
    .Y(_07160_));
 sky130_fd_sc_hd__nand2_1 _18927_ (.A(_07153_),
    .B(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__a21oi_2 _18928_ (.A1(_14091_),
    .A2(_07161_),
    .B1(_14090_),
    .Y(_07162_));
 sky130_fd_sc_hd__xnor2_4 _18929_ (.A(_14100_),
    .B(_07162_),
    .Y(_12715_));
 sky130_fd_sc_hd__inv_1 _18930_ (.A(_12715_),
    .Y(_12884_));
 sky130_fd_sc_hd__nor2_1 _18931_ (.A(_14065_),
    .B(_14090_),
    .Y(_07163_));
 sky130_fd_sc_hd__nand2_1 _18932_ (.A(_07153_),
    .B(_07163_),
    .Y(_07164_));
 sky130_fd_sc_hd__a21oi_1 _18933_ (.A1(_14066_),
    .A2(_07134_),
    .B1(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__a21boi_0 _18934_ (.A1(_07153_),
    .A2(_07152_),
    .B1_N(_14091_),
    .Y(_07166_));
 sky130_fd_sc_hd__o21ai_1 _18935_ (.A1(_14090_),
    .A2(_07166_),
    .B1(_14100_),
    .Y(_07167_));
 sky130_fd_sc_hd__o21bai_2 _18936_ (.A1(_07165_),
    .A2(_07167_),
    .B1_N(_14099_),
    .Y(_07168_));
 sky130_fd_sc_hd__xnor2_4 _18937_ (.A(_14109_),
    .B(_07168_),
    .Y(_12720_));
 sky130_fd_sc_hd__inv_1 _18938_ (.A(_14095_),
    .Y(_07169_));
 sky130_fd_sc_hd__a211oi_4 _18939_ (.A1(_07137_),
    .A2(_07155_),
    .B1(_07158_),
    .C1(_07169_),
    .Y(_07170_));
 sky130_fd_sc_hd__o21ai_1 _18940_ (.A1(_14094_),
    .A2(_07170_),
    .B1(_14104_),
    .Y(_07171_));
 sky130_fd_sc_hd__nand2b_1 _18941_ (.A_N(_14103_),
    .B(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__xor2_2 _18942_ (.A(_14113_),
    .B(_07172_),
    .X(_12899_));
 sky130_fd_sc_hd__inv_1 _18943_ (.A(_12899_),
    .Y(_12719_));
 sky130_fd_sc_hd__nand2_1 _18944_ (.A(_14091_),
    .B(_14100_),
    .Y(_07173_));
 sky130_fd_sc_hd__a211oi_1 _18945_ (.A1(_07139_),
    .A2(_07140_),
    .B1(_07152_),
    .C1(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__o31a_1 _18946_ (.A1(_14055_),
    .A2(_14065_),
    .A3(_07144_),
    .B1(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__nand2_1 _18947_ (.A(_14100_),
    .B(_14090_),
    .Y(_07176_));
 sky130_fd_sc_hd__o21ai_1 _18948_ (.A1(_07153_),
    .A2(_07173_),
    .B1(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__o31ai_1 _18949_ (.A1(_14099_),
    .A2(_07175_),
    .A3(_07177_),
    .B1(_14109_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2b_1 _18950_ (.A_N(_14108_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__xor2_4 _18951_ (.A(_14118_),
    .B(_07179_),
    .X(_12902_));
 sky130_fd_sc_hd__inv_1 _18952_ (.A(_12902_),
    .Y(_12725_));
 sky130_fd_sc_hd__nand3_1 _18953_ (.A(_14087_),
    .B(_14095_),
    .C(_14104_),
    .Y(_07180_));
 sky130_fd_sc_hd__a21o_1 _18954_ (.A1(_14095_),
    .A2(_14086_),
    .B1(_14094_),
    .X(_07181_));
 sky130_fd_sc_hd__nand2_1 _18955_ (.A(_14104_),
    .B(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__o21ai_4 _18956_ (.A1(_07151_),
    .A2(_07180_),
    .B1(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__o21ai_0 _18957_ (.A1(_14103_),
    .A2(_07183_),
    .B1(_14113_),
    .Y(_07184_));
 sky130_fd_sc_hd__nand2b_1 _18958_ (.A_N(_14112_),
    .B(_07184_),
    .Y(_07185_));
 sky130_fd_sc_hd__xor2_2 _18959_ (.A(_14122_),
    .B(_07185_),
    .X(_12908_));
 sky130_fd_sc_hd__inv_1 _18960_ (.A(_12908_),
    .Y(_12724_));
 sky130_fd_sc_hd__and2_0 _18961_ (.A(_14109_),
    .B(_14118_),
    .X(_07186_));
 sky130_fd_sc_hd__nor3b_2 _18962_ (.A(_07165_),
    .B(_07167_),
    .C_N(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__a22oi_1 _18963_ (.A1(_14118_),
    .A2(_14108_),
    .B1(_07186_),
    .B2(_14099_),
    .Y(_07188_));
 sky130_fd_sc_hd__nand2b_1 _18964_ (.A_N(_14117_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__o21ai_0 _18965_ (.A1(_07187_),
    .A2(_07189_),
    .B1(_14128_),
    .Y(_07190_));
 sky130_fd_sc_hd__nand2b_1 _18966_ (.A_N(_14127_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__a21oi_2 _18967_ (.A1(_14137_),
    .A2(_07191_),
    .B1(_14136_),
    .Y(_07192_));
 sky130_fd_sc_hd__xor2_4 _18968_ (.A(_14145_),
    .B(_07192_),
    .X(_12740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1123 ();
 sky130_fd_sc_hd__or4_1 _18970_ (.A(_14094_),
    .B(_14103_),
    .C(_14112_),
    .D(_14121_),
    .X(_07194_));
 sky130_fd_sc_hd__o21a_1 _18971_ (.A1(_14104_),
    .A2(_14103_),
    .B1(_14113_),
    .X(_07195_));
 sky130_fd_sc_hd__o21ai_0 _18972_ (.A1(_14112_),
    .A2(_07195_),
    .B1(_14122_),
    .Y(_07196_));
 sky130_fd_sc_hd__nand2b_1 _18973_ (.A_N(_14121_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__o21a_2 _18974_ (.A1(_07170_),
    .A2(_07194_),
    .B1(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__a21o_1 _18975_ (.A1(_07198_),
    .A2(_14132_),
    .B1(_14131_),
    .X(_07199_));
 sky130_fd_sc_hd__a21o_1 _18976_ (.A1(_07199_),
    .A2(_14141_),
    .B1(_14140_),
    .X(_07200_));
 sky130_fd_sc_hd__xor2_2 _18977_ (.A(_14149_),
    .B(_07200_),
    .X(_12927_));
 sky130_fd_sc_hd__inv_2 _18978_ (.A(_12927_),
    .Y(_12739_));
 sky130_fd_sc_hd__o211ai_1 _18979_ (.A1(_07175_),
    .A2(_07177_),
    .B1(_07186_),
    .C1(_14128_),
    .Y(_07201_));
 sky130_fd_sc_hd__a21oi_1 _18980_ (.A1(_14128_),
    .A2(_07189_),
    .B1(_14127_),
    .Y(_07202_));
 sky130_fd_sc_hd__a21boi_0 _18981_ (.A1(_07201_),
    .A2(_07202_),
    .B1_N(_14137_),
    .Y(_07203_));
 sky130_fd_sc_hd__or2_0 _18982_ (.A(_14136_),
    .B(_07203_),
    .X(_07204_));
 sky130_fd_sc_hd__a21oi_2 _18983_ (.A1(_14145_),
    .A2(_07204_),
    .B1(_14144_),
    .Y(_07205_));
 sky130_fd_sc_hd__xor2_4 _18984_ (.A(_14154_),
    .B(_07205_),
    .X(_12745_));
 sky130_fd_sc_hd__inv_1 _18985_ (.A(_14158_),
    .Y(_07206_));
 sky130_fd_sc_hd__inv_1 _18986_ (.A(_14132_),
    .Y(_07207_));
 sky130_fd_sc_hd__a21o_1 _18987_ (.A1(_14113_),
    .A2(_14103_),
    .B1(_14112_),
    .X(_07208_));
 sky130_fd_sc_hd__a21oi_1 _18988_ (.A1(_14122_),
    .A2(_07208_),
    .B1(_14121_),
    .Y(_07209_));
 sky130_fd_sc_hd__o21bai_1 _18989_ (.A1(_07207_),
    .A2(_07209_),
    .B1_N(_14131_),
    .Y(_07210_));
 sky130_fd_sc_hd__a41oi_4 _18990_ (.A1(_14122_),
    .A2(_07183_),
    .A3(_14132_),
    .A4(_14113_),
    .B1(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__nor2b_1 _18991_ (.A(_07211_),
    .B_N(_14141_),
    .Y(_07212_));
 sky130_fd_sc_hd__o21ai_1 _18992_ (.A1(_14140_),
    .A2(_07212_),
    .B1(_14149_),
    .Y(_07213_));
 sky130_fd_sc_hd__nand2b_1 _18993_ (.A_N(_14148_),
    .B(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__xnor2_1 _18994_ (.A(_07206_),
    .B(_07214_),
    .Y(_12935_));
 sky130_fd_sc_hd__inv_1 _18995_ (.A(_12935_),
    .Y(_12744_));
 sky130_fd_sc_hd__inv_1 _18996_ (.A(_07188_),
    .Y(_07215_));
 sky130_fd_sc_hd__and4_1 _18997_ (.A(_14128_),
    .B(_14137_),
    .C(_14145_),
    .D(_14154_),
    .X(_07216_));
 sky130_fd_sc_hd__o21ai_2 _18998_ (.A1(_07187_),
    .A2(_07215_),
    .B1(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__a21o_1 _18999_ (.A1(_14137_),
    .A2(_14127_),
    .B1(_14136_),
    .X(_07218_));
 sky130_fd_sc_hd__a21oi_1 _19000_ (.A1(_14145_),
    .A2(_07218_),
    .B1(_14144_),
    .Y(_07219_));
 sky130_fd_sc_hd__nor2b_1 _19001_ (.A(_07219_),
    .B_N(_14154_),
    .Y(_07220_));
 sky130_fd_sc_hd__a21oi_2 _19002_ (.A1(_14117_),
    .A2(_07216_),
    .B1(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__nor3_1 _19003_ (.A(_14153_),
    .B(_14163_),
    .C(_14172_),
    .Y(_07222_));
 sky130_fd_sc_hd__or2_0 _19004_ (.A(_14164_),
    .B(_14163_),
    .X(_07223_));
 sky130_fd_sc_hd__a21oi_1 _19005_ (.A1(_14173_),
    .A2(_07223_),
    .B1(_14172_),
    .Y(_07224_));
 sky130_fd_sc_hd__a31oi_4 _19006_ (.A1(_07217_),
    .A2(_07221_),
    .A3(_07222_),
    .B1(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__a21o_1 _19007_ (.A1(_14181_),
    .A2(_07225_),
    .B1(_14180_),
    .X(_07226_));
 sky130_fd_sc_hd__a21oi_4 _19008_ (.A1(_14189_),
    .A2(_07226_),
    .B1(_14188_),
    .Y(_07227_));
 sky130_fd_sc_hd__xnor2_4 _19009_ (.A(_14197_),
    .B(_07227_),
    .Y(_12770_));
 sky130_fd_sc_hd__inv_1 _19010_ (.A(_12770_),
    .Y(_12963_));
 sky130_fd_sc_hd__a211o_1 _19011_ (.A1(_14164_),
    .A2(_14153_),
    .B1(_14163_),
    .C1(_14144_),
    .X(_07228_));
 sky130_fd_sc_hd__o21a_1 _19012_ (.A1(_14145_),
    .A2(_14144_),
    .B1(_14154_),
    .X(_07229_));
 sky130_fd_sc_hd__o21ai_0 _19013_ (.A1(_14153_),
    .A2(_07229_),
    .B1(_14164_),
    .Y(_07230_));
 sky130_fd_sc_hd__nand2b_1 _19014_ (.A_N(_14163_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__a21oi_1 _19015_ (.A1(_14173_),
    .A2(_07231_),
    .B1(_14172_),
    .Y(_07232_));
 sky130_fd_sc_hd__nor2b_1 _19016_ (.A(_07232_),
    .B_N(_14181_),
    .Y(_07233_));
 sky130_fd_sc_hd__o41a_2 _19017_ (.A1(_14136_),
    .A2(_14172_),
    .A3(_07203_),
    .A4(_07228_),
    .B1(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__o21ai_0 _19018_ (.A1(_14180_),
    .A2(_07234_),
    .B1(_14189_),
    .Y(_07235_));
 sky130_fd_sc_hd__nand2b_1 _19019_ (.A_N(_14188_),
    .B(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__a21oi_2 _19020_ (.A1(_14197_),
    .A2(_07236_),
    .B1(_14196_),
    .Y(_07237_));
 sky130_fd_sc_hd__xnor2_4 _19021_ (.A(_14205_),
    .B(_07237_),
    .Y(_12972_));
 sky130_fd_sc_hd__inv_1 _19022_ (.A(_12972_),
    .Y(_12775_));
 sky130_fd_sc_hd__nand3_1 _19023_ (.A(_14141_),
    .B(_14149_),
    .C(_14158_),
    .Y(_07238_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1120 ();
 sky130_fd_sc_hd__nand4_1 _19027_ (.A(_14168_),
    .B(_14177_),
    .C(_14185_),
    .D(_14193_),
    .Y(_07242_));
 sky130_fd_sc_hd__a21oi_1 _19028_ (.A1(_14149_),
    .A2(_14140_),
    .B1(_14148_),
    .Y(_07243_));
 sky130_fd_sc_hd__o21bai_1 _19029_ (.A1(_07206_),
    .A2(_07243_),
    .B1_N(_14157_),
    .Y(_07244_));
 sky130_fd_sc_hd__a21oi_1 _19030_ (.A1(_14168_),
    .A2(_07244_),
    .B1(_14167_),
    .Y(_07245_));
 sky130_fd_sc_hd__nand2_1 _19031_ (.A(_14177_),
    .B(_14185_),
    .Y(_07246_));
 sky130_fd_sc_hd__a21oi_1 _19032_ (.A1(_14185_),
    .A2(_14176_),
    .B1(_14184_),
    .Y(_07247_));
 sky130_fd_sc_hd__o21ai_0 _19033_ (.A1(_07245_),
    .A2(_07246_),
    .B1(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__a21oi_2 _19034_ (.A1(_14193_),
    .A2(_07248_),
    .B1(_14192_),
    .Y(_07249_));
 sky130_fd_sc_hd__o31ai_4 _19035_ (.A1(net1112),
    .A2(_07238_),
    .A3(_07242_),
    .B1(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__a21oi_2 _19036_ (.A1(_07250_),
    .A2(_14201_),
    .B1(_14200_),
    .Y(_07251_));
 sky130_fd_sc_hd__xnor2_2 _19037_ (.A(_14209_),
    .B(_07251_),
    .Y(_12978_));
 sky130_fd_sc_hd__inv_1 _19038_ (.A(_12978_),
    .Y(_12774_));
 sky130_fd_sc_hd__inv_1 _19039_ (.A(_14197_),
    .Y(_07252_));
 sky130_fd_sc_hd__o21bai_1 _19040_ (.A1(_07252_),
    .A2(_07227_),
    .B1_N(_14196_),
    .Y(_07253_));
 sky130_fd_sc_hd__a21oi_2 _19041_ (.A1(_14205_),
    .A2(_07253_),
    .B1(_14204_),
    .Y(_07254_));
 sky130_fd_sc_hd__xor2_4 _19042_ (.A(_14214_),
    .B(_07254_),
    .X(_12780_));
 sky130_fd_sc_hd__nand2_1 _19043_ (.A(_14141_),
    .B(_14149_),
    .Y(_07255_));
 sky130_fd_sc_hd__nor3_1 _19044_ (.A(_07207_),
    .B(_07206_),
    .C(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__o211ai_2 _19045_ (.A1(_07170_),
    .A2(_07194_),
    .B1(_07197_),
    .C1(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__nor2_1 _19046_ (.A(_07206_),
    .B(_07243_),
    .Y(_07258_));
 sky130_fd_sc_hd__a41oi_2 _19047_ (.A1(_14141_),
    .A2(_14149_),
    .A3(_14158_),
    .A4(_14131_),
    .B1(_07258_),
    .Y(_07259_));
 sky130_fd_sc_hd__a21o_1 _19048_ (.A1(_14177_),
    .A2(_14167_),
    .B1(_14176_),
    .X(_07260_));
 sky130_fd_sc_hd__a211oi_1 _19049_ (.A1(_14185_),
    .A2(_07260_),
    .B1(_14184_),
    .C1(_14157_),
    .Y(_07261_));
 sky130_fd_sc_hd__o21a_1 _19050_ (.A1(_14168_),
    .A2(_14167_),
    .B1(_14177_),
    .X(_07262_));
 sky130_fd_sc_hd__o21a_1 _19051_ (.A1(_14176_),
    .A2(_07262_),
    .B1(_14185_),
    .X(_07263_));
 sky130_fd_sc_hd__o21ai_0 _19052_ (.A1(_14184_),
    .A2(_07263_),
    .B1(_14193_),
    .Y(_07264_));
 sky130_fd_sc_hd__a31oi_2 _19053_ (.A1(_07257_),
    .A2(_07259_),
    .A3(_07261_),
    .B1(_07264_),
    .Y(_07265_));
 sky130_fd_sc_hd__inv_1 _19054_ (.A(_14209_),
    .Y(_07266_));
 sky130_fd_sc_hd__nor2_1 _19055_ (.A(_14201_),
    .B(_14200_),
    .Y(_07267_));
 sky130_fd_sc_hd__o21bai_1 _19056_ (.A1(_07266_),
    .A2(_07267_),
    .B1_N(_14208_),
    .Y(_07268_));
 sky130_fd_sc_hd__o41a_2 _19057_ (.A1(_14192_),
    .A2(_14200_),
    .A3(_14208_),
    .A4(_07265_),
    .B1(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__xor2_1 _19058_ (.A(_14218_),
    .B(_07269_),
    .X(_12985_));
 sky130_fd_sc_hd__inv_1 _19059_ (.A(_12985_),
    .Y(_12779_));
 sky130_fd_sc_hd__and3_1 _19060_ (.A(_14197_),
    .B(_14205_),
    .C(_14214_),
    .X(_07270_));
 sky130_fd_sc_hd__a21oi_1 _19061_ (.A1(_14197_),
    .A2(_14188_),
    .B1(_14196_),
    .Y(_07271_));
 sky130_fd_sc_hd__nor2b_1 _19062_ (.A(_07271_),
    .B_N(_14205_),
    .Y(_07272_));
 sky130_fd_sc_hd__o21ai_0 _19063_ (.A1(_14204_),
    .A2(_07272_),
    .B1(_14214_),
    .Y(_07273_));
 sky130_fd_sc_hd__a31oi_1 _19064_ (.A1(_14189_),
    .A2(_14180_),
    .A3(_07270_),
    .B1(_14213_),
    .Y(_07274_));
 sky130_fd_sc_hd__nand2_1 _19065_ (.A(_07273_),
    .B(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__a31oi_4 _19066_ (.A1(_14189_),
    .A2(_07234_),
    .A3(_07270_),
    .B1(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__xnor2_4 _19067_ (.A(_14224_),
    .B(_07276_),
    .Y(_12988_));
 sky130_fd_sc_hd__inv_1 _19068_ (.A(_12988_),
    .Y(_12785_));
 sky130_fd_sc_hd__nor2_1 _19069_ (.A(_07251_),
    .B(_07266_),
    .Y(_07277_));
 sky130_fd_sc_hd__o21ai_1 _19070_ (.A1(_07277_),
    .A2(_14208_),
    .B1(_14218_),
    .Y(_07278_));
 sky130_fd_sc_hd__nand2b_1 _19071_ (.A_N(_14217_),
    .B(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__xor2_2 _19072_ (.A(_14228_),
    .B(_07279_),
    .X(_12994_));
 sky130_fd_sc_hd__inv_1 _19073_ (.A(_12994_),
    .Y(_12784_));
 sky130_fd_sc_hd__nand2_1 _19074_ (.A(_14224_),
    .B(_07270_),
    .Y(_07280_));
 sky130_fd_sc_hd__a21o_1 _19075_ (.A1(_14205_),
    .A2(_14196_),
    .B1(_14204_),
    .X(_07281_));
 sky130_fd_sc_hd__a21o_1 _19076_ (.A1(_14214_),
    .A2(_07281_),
    .B1(_14213_),
    .X(_07282_));
 sky130_fd_sc_hd__a21oi_1 _19077_ (.A1(_14224_),
    .A2(_07282_),
    .B1(_14223_),
    .Y(_07283_));
 sky130_fd_sc_hd__o21ai_2 _19078_ (.A1(_07227_),
    .A2(_07280_),
    .B1(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__xnor2_4 _19079_ (.A(_14234_),
    .B(_07284_),
    .Y(_12790_));
 sky130_fd_sc_hd__and2_0 _19080_ (.A(_14218_),
    .B(_14228_),
    .X(_07285_));
 sky130_fd_sc_hd__a221oi_4 _19081_ (.A1(_14228_),
    .A2(_14217_),
    .B1(_07269_),
    .B2(_07285_),
    .C1(_14227_),
    .Y(_07286_));
 sky130_fd_sc_hd__xnor2_1 _19082_ (.A(_14238_),
    .B(_07286_),
    .Y(_13001_));
 sky130_fd_sc_hd__inv_1 _19083_ (.A(_13001_),
    .Y(_12789_));
 sky130_fd_sc_hd__nand2_1 _19084_ (.A(_14224_),
    .B(_14234_),
    .Y(_07287_));
 sky130_fd_sc_hd__a21oi_1 _19085_ (.A1(_14234_),
    .A2(_14223_),
    .B1(_14233_),
    .Y(_07288_));
 sky130_fd_sc_hd__o21ai_2 _19086_ (.A1(_07276_),
    .A2(_07287_),
    .B1(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__xor2_4 _19087_ (.A(_14244_),
    .B(_07289_),
    .X(_13004_));
 sky130_fd_sc_hd__inv_1 _19088_ (.A(_13004_),
    .Y(_12795_));
 sky130_fd_sc_hd__nor2_2 _19089_ (.A(_07238_),
    .B(_07242_),
    .Y(_07290_));
 sky130_fd_sc_hd__and3_1 _19090_ (.A(_14113_),
    .B(_14122_),
    .C(_14132_),
    .X(_07291_));
 sky130_fd_sc_hd__nand2_1 _19091_ (.A(_14132_),
    .B(_07290_),
    .Y(_07292_));
 sky130_fd_sc_hd__nand2_1 _19092_ (.A(_14131_),
    .B(_07290_),
    .Y(_07293_));
 sky130_fd_sc_hd__o21ai_1 _19093_ (.A1(_07209_),
    .A2(_07292_),
    .B1(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__a311oi_4 _19094_ (.A1(_07183_),
    .A2(_07290_),
    .A3(_07291_),
    .B1(_07294_),
    .C1(_14200_),
    .Y(_07295_));
 sky130_fd_sc_hd__nand2_1 _19095_ (.A(_14238_),
    .B(_07285_),
    .Y(_07296_));
 sky130_fd_sc_hd__a2111oi_2 _19096_ (.A1(_07249_),
    .A2(_07295_),
    .B1(_07267_),
    .C1(_07296_),
    .D1(_07266_),
    .Y(_07297_));
 sky130_fd_sc_hd__inv_1 _19097_ (.A(_14238_),
    .Y(_07298_));
 sky130_fd_sc_hd__a21o_1 _19098_ (.A1(_14218_),
    .A2(_14208_),
    .B1(_14217_),
    .X(_07299_));
 sky130_fd_sc_hd__a21oi_1 _19099_ (.A1(_14228_),
    .A2(_07299_),
    .B1(_14227_),
    .Y(_07300_));
 sky130_fd_sc_hd__nor2_1 _19100_ (.A(_07298_),
    .B(_07300_),
    .Y(_07301_));
 sky130_fd_sc_hd__nor3_2 _19101_ (.A(_14237_),
    .B(_07297_),
    .C(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__xnor2_1 _19102_ (.A(_14248_),
    .B(_07302_),
    .Y(_13010_));
 sky130_fd_sc_hd__inv_1 _19103_ (.A(_13010_),
    .Y(_12794_));
 sky130_fd_sc_hd__nand2_2 _19104_ (.A(_14244_),
    .B(_14254_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand2_1 _19105_ (.A(_14254_),
    .B(_14243_),
    .Y(_07304_));
 sky130_fd_sc_hd__o21a_1 _19106_ (.A1(_07288_),
    .A2(_07303_),
    .B1(_07304_),
    .X(_07305_));
 sky130_fd_sc_hd__o31ai_4 _19107_ (.A1(_07276_),
    .A2(_07287_),
    .A3(_07303_),
    .B1(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__nor2_2 _19108_ (.A(_14253_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__xnor2_4 _19109_ (.A(_14263_),
    .B(_07307_),
    .Y(_13019_));
 sky130_fd_sc_hd__inv_1 _19110_ (.A(_13019_),
    .Y(_12805_));
 sky130_fd_sc_hd__nor2b_1 _19111_ (.A(_07302_),
    .B_N(_14248_),
    .Y(_07308_));
 sky130_fd_sc_hd__o21ai_0 _19112_ (.A1(_14247_),
    .A2(_07308_),
    .B1(_14258_),
    .Y(_07309_));
 sky130_fd_sc_hd__nand2b_1 _19113_ (.A_N(_14257_),
    .B(_07309_),
    .Y(_07310_));
 sky130_fd_sc_hd__xor2_1 _19114_ (.A(_14267_),
    .B(_07310_),
    .X(_13024_));
 sky130_fd_sc_hd__inv_1 _19115_ (.A(_13024_),
    .Y(_12804_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1119 ();
 sky130_fd_sc_hd__inv_1 _19117_ (.A(_14263_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand3_1 _19118_ (.A(_14224_),
    .B(_14234_),
    .C(_07270_),
    .Y(_07313_));
 sky130_fd_sc_hd__nor3_2 _19119_ (.A(_07227_),
    .B(_07303_),
    .C(_07313_),
    .Y(_07314_));
 sky130_fd_sc_hd__nor2b_1 _19120_ (.A(_07283_),
    .B_N(_14234_),
    .Y(_07315_));
 sky130_fd_sc_hd__nor2_1 _19121_ (.A(_14233_),
    .B(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__o21ai_2 _19122_ (.A1(_07303_),
    .A2(_07316_),
    .B1(_07304_),
    .Y(_07317_));
 sky130_fd_sc_hd__nor3_1 _19123_ (.A(_14253_),
    .B(_07314_),
    .C(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__o21bai_4 _19124_ (.A1(_07312_),
    .A2(_07318_),
    .B1_N(_14262_),
    .Y(_07319_));
 sky130_fd_sc_hd__xnor2_4 _19125_ (.A(_14272_),
    .B(_07319_),
    .Y(_12810_));
 sky130_fd_sc_hd__o21bai_2 _19126_ (.A1(_07298_),
    .A2(_07286_),
    .B1_N(_14237_),
    .Y(_07320_));
 sky130_fd_sc_hd__nand2_1 _19127_ (.A(_14248_),
    .B(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__nor3_1 _19128_ (.A(_14247_),
    .B(_14257_),
    .C(_14266_),
    .Y(_07322_));
 sky130_fd_sc_hd__or2_0 _19129_ (.A(_14258_),
    .B(_14257_),
    .X(_07323_));
 sky130_fd_sc_hd__a21oi_1 _19130_ (.A1(_14267_),
    .A2(_07323_),
    .B1(_14266_),
    .Y(_07324_));
 sky130_fd_sc_hd__a21oi_2 _19131_ (.A1(_07321_),
    .A2(_07322_),
    .B1(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__xnor2_1 _19132_ (.A(_14276_),
    .B(_07325_),
    .Y(_12809_));
 sky130_fd_sc_hd__o2111ai_2 _19133_ (.A1(_07314_),
    .A2(_07317_),
    .B1(_14263_),
    .C1(_14272_),
    .D1(_14282_),
    .Y(_07326_));
 sky130_fd_sc_hd__a21o_1 _19134_ (.A1(_14263_),
    .A2(_14253_),
    .B1(_14262_),
    .X(_07327_));
 sky130_fd_sc_hd__a21o_1 _19135_ (.A1(_14272_),
    .A2(_07327_),
    .B1(_14271_),
    .X(_07328_));
 sky130_fd_sc_hd__a21oi_1 _19136_ (.A1(_14282_),
    .A2(_07328_),
    .B1(_14281_),
    .Y(_07329_));
 sky130_fd_sc_hd__nand2_4 _19137_ (.A(_07326_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__xnor2_4 _19138_ (.A(_14291_),
    .B(_07330_),
    .Y(_12820_));
 sky130_fd_sc_hd__nand2_1 _19139_ (.A(_14276_),
    .B(_14286_),
    .Y(_07331_));
 sky130_fd_sc_hd__nand3_1 _19140_ (.A(_14248_),
    .B(_14258_),
    .C(_14267_),
    .Y(_07332_));
 sky130_fd_sc_hd__nor2_1 _19141_ (.A(_07331_),
    .B(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__nand3_1 _19142_ (.A(_14258_),
    .B(_14267_),
    .C(_14247_),
    .Y(_07334_));
 sky130_fd_sc_hd__a21oi_1 _19143_ (.A1(_14267_),
    .A2(_14257_),
    .B1(_14266_),
    .Y(_07335_));
 sky130_fd_sc_hd__a21boi_0 _19144_ (.A1(_07334_),
    .A2(_07335_),
    .B1_N(_14276_),
    .Y(_07336_));
 sky130_fd_sc_hd__o21ai_0 _19145_ (.A1(_14275_),
    .A2(_07336_),
    .B1(_14286_),
    .Y(_07337_));
 sky130_fd_sc_hd__nand2b_1 _19146_ (.A_N(_14285_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__a21oi_1 _19147_ (.A1(_07320_),
    .A2(_07333_),
    .B1(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__xor2_2 _19148_ (.A(_14295_),
    .B(_07339_),
    .X(_12819_));
 sky130_fd_sc_hd__nor2_1 _19149_ (.A(_07156_),
    .B(_07151_),
    .Y(_07340_));
 sky130_fd_sc_hd__o21ai_0 _19150_ (.A1(_14086_),
    .A2(_07340_),
    .B1(_14095_),
    .Y(_07341_));
 sky130_fd_sc_hd__nor2_1 _19151_ (.A(_14104_),
    .B(_14094_),
    .Y(_07342_));
 sky130_fd_sc_hd__a21oi_1 _19152_ (.A1(_07341_),
    .A2(_07342_),
    .B1(_07183_),
    .Y(_12891_));
 sky130_fd_sc_hd__xnor2_2 _19153_ (.A(_07207_),
    .B(_07198_),
    .Y(_12914_));
 sky130_fd_sc_hd__xnor2_1 _19154_ (.A(_14141_),
    .B(_07211_),
    .Y(_12920_));
 sky130_fd_sc_hd__nor2b_4 _19155_ (.A(_07238_),
    .B_N(_07199_),
    .Y(_07343_));
 sky130_fd_sc_hd__nor2_1 _19156_ (.A(_07244_),
    .B(_07343_),
    .Y(_07344_));
 sky130_fd_sc_hd__xnor2_1 _19157_ (.A(_14168_),
    .B(_07344_),
    .Y(_12942_));
 sky130_fd_sc_hd__a21o_1 _19158_ (.A1(_14158_),
    .A2(_07214_),
    .B1(_14157_),
    .X(_07345_));
 sky130_fd_sc_hd__a21oi_4 _19159_ (.A1(_07345_),
    .A2(_14168_),
    .B1(_14167_),
    .Y(_07346_));
 sky130_fd_sc_hd__xnor2_1 _19160_ (.A(_14177_),
    .B(_07346_),
    .Y(_12948_));
 sky130_fd_sc_hd__o21ai_1 _19161_ (.A1(_07244_),
    .A2(_07343_),
    .B1(_14168_),
    .Y(_07347_));
 sky130_fd_sc_hd__nand2b_1 _19162_ (.A_N(_14167_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__a21oi_2 _19163_ (.A1(_07348_),
    .A2(_14177_),
    .B1(_14176_),
    .Y(_07349_));
 sky130_fd_sc_hd__xnor2_2 _19164_ (.A(_14185_),
    .B(_07349_),
    .Y(_12954_));
 sky130_fd_sc_hd__o21a_2 _19165_ (.A1(_07246_),
    .A2(_07346_),
    .B1(_07247_),
    .X(_07350_));
 sky130_fd_sc_hd__xnor2_2 _19166_ (.A(_14193_),
    .B(_07350_),
    .Y(_12960_));
 sky130_fd_sc_hd__nor2_1 _19167_ (.A(_14192_),
    .B(_07265_),
    .Y(_07351_));
 sky130_fd_sc_hd__xnor2_1 _19168_ (.A(_14201_),
    .B(_07351_),
    .Y(_12969_));
 sky130_fd_sc_hd__a21oi_2 _19169_ (.A1(_14248_),
    .A2(_07320_),
    .B1(_14247_),
    .Y(_07352_));
 sky130_fd_sc_hd__xnor2_1 _19170_ (.A(_14258_),
    .B(_07352_),
    .Y(_13016_));
 sky130_fd_sc_hd__xor2_1 _19171_ (.A(_14276_),
    .B(_07325_),
    .X(_13032_));
 sky130_fd_sc_hd__a21o_1 _19172_ (.A1(_14267_),
    .A2(_07310_),
    .B1(_14266_),
    .X(_07353_));
 sky130_fd_sc_hd__a21oi_2 _19173_ (.A1(_14276_),
    .A2(_07353_),
    .B1(_14275_),
    .Y(_07354_));
 sky130_fd_sc_hd__xnor2_1 _19174_ (.A(_14286_),
    .B(_07354_),
    .Y(_13038_));
 sky130_fd_sc_hd__clkinv_16 _19175_ (.A(net1019),
    .Y(_00906_));
 sky130_fd_sc_hd__inv_1 _19176_ (.A(_13156_),
    .Y(_11771_));
 sky130_fd_sc_hd__inv_1 _19177_ (.A(_13279_),
    .Y(_12019_));
 sky130_fd_sc_hd__inv_2 _19178_ (.A(_13399_),
    .Y(_12254_));
 sky130_fd_sc_hd__inv_1 _19179_ (.A(_13408_),
    .Y(_12277_));
 sky130_fd_sc_hd__inv_1 _19180_ (.A(\hash.CA1.k_i2[1] ),
    .Y(_12537_));
 sky130_fd_sc_hd__inv_1 _19181_ (.A(\hash.CA1.k_i2[0] ),
    .Y(_12542_));
 sky130_fd_sc_hd__inv_1 _19182_ (.A(\hash.CA1.k_i2[3] ),
    .Y(_12552_));
 sky130_fd_sc_hd__inv_1 _19183_ (.A(\hash.CA1.k_i2[5] ),
    .Y(_12560_));
 sky130_fd_sc_hd__inv_1 _19184_ (.A(\hash.CA1.k_i2[7] ),
    .Y(_12568_));
 sky130_fd_sc_hd__inv_1 _19185_ (.A(\hash.CA1.k_i2[8] ),
    .Y(_12573_));
 sky130_fd_sc_hd__inv_1 _19186_ (.A(\hash.CA1.k_i2[11] ),
    .Y(_12584_));
 sky130_fd_sc_hd__inv_1 _19187_ (.A(\hash.CA1.k_i2[12] ),
    .Y(_12589_));
 sky130_fd_sc_hd__inv_1 _19188_ (.A(\hash.CA1.k_i2[14] ),
    .Y(_12597_));
 sky130_fd_sc_hd__inv_1 _19189_ (.A(\hash.CA1.k_i2[15] ),
    .Y(_12602_));
 sky130_fd_sc_hd__inv_1 _19190_ (.A(\hash.CA1.k_i2[16] ),
    .Y(_12607_));
 sky130_fd_sc_hd__inv_1 _19191_ (.A(\hash.CA1.k_i2[17] ),
    .Y(_12612_));
 sky130_fd_sc_hd__inv_1 _19192_ (.A(\hash.CA1.k_i2[23] ),
    .Y(_12632_));
 sky130_fd_sc_hd__inv_1 _19193_ (.A(\hash.CA1.k_i2[24] ),
    .Y(_12637_));
 sky130_fd_sc_hd__inv_1 _19194_ (.A(\hash.CA1.k_i2[25] ),
    .Y(_12642_));
 sky130_fd_sc_hd__inv_1 _19195_ (.A(\hash.CA1.k_i2[26] ),
    .Y(_12647_));
 sky130_fd_sc_hd__inv_1 _19196_ (.A(\hash.CA1.k_i2[27] ),
    .Y(_12652_));
 sky130_fd_sc_hd__clkinv_2 _19197_ (.A(\hash.CA1.k_i2[28] ),
    .Y(_12657_));
 sky130_fd_sc_hd__inv_2 _19198_ (.A(_14031_),
    .Y(_12671_));
 sky130_fd_sc_hd__inv_1 _19199_ (.A(_14375_),
    .Y(_13050_));
 sky130_fd_sc_hd__inv_1 _19200_ (.A(_14378_),
    .Y(_13054_));
 sky130_fd_sc_hd__inv_1 _19201_ (.A(_14379_),
    .Y(_13059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1115 ();
 sky130_fd_sc_hd__mux4_1 _19206_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[1] ),
    .X(_07359_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1111 ();
 sky130_fd_sc_hd__mux4_1 _19211_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[1] ),
    .X(_07364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1109 ();
 sky130_fd_sc_hd__mux4_1 _19214_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[1] ),
    .X(_07367_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1106 ();
 sky130_fd_sc_hd__mux4_1 _19218_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07371_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1102 ();
 sky130_fd_sc_hd__mux4_4 _19223_ (.A0(_07359_),
    .A1(_07364_),
    .A2(_07367_),
    .A3(_07371_),
    .S0(net579),
    .S1(net575),
    .X(_07376_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1100 ();
 sky130_fd_sc_hd__mux4_1 _19226_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07379_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1098 ();
 sky130_fd_sc_hd__mux4_1 _19229_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07382_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1096 ();
 sky130_fd_sc_hd__mux4_1 _19232_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07385_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1094 ();
 sky130_fd_sc_hd__mux4_1 _19235_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1092 ();
 sky130_fd_sc_hd__mux4_1 _19238_ (.A0(_07379_),
    .A1(_07382_),
    .A2(_07385_),
    .A3(_07388_),
    .S0(net579),
    .S1(net575),
    .X(_07391_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1091 ();
 sky130_fd_sc_hd__mux2i_4 _19240_ (.A0(_07376_),
    .A1(_07391_),
    .S(net573),
    .Y(_11751_));
 sky130_fd_sc_hd__mux4_1 _19241_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(\count7_1[2] ),
    .S1(net591),
    .X(_07393_));
 sky130_fd_sc_hd__mux4_1 _19242_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[1] ),
    .X(_07394_));
 sky130_fd_sc_hd__mux4_1 _19243_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[1] ),
    .X(_07395_));
 sky130_fd_sc_hd__mux4_1 _19244_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[1] ),
    .X(_07396_));
 sky130_fd_sc_hd__mux4_4 _19245_ (.A0(_07393_),
    .A1(_07394_),
    .A2(_07395_),
    .A3(_07396_),
    .S0(net579),
    .S1(net575),
    .X(_07397_));
 sky130_fd_sc_hd__mux4_1 _19246_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net583),
    .S1(net590),
    .X(_07398_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1090 ();
 sky130_fd_sc_hd__mux4_1 _19248_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net583),
    .S1(net590),
    .X(_07400_));
 sky130_fd_sc_hd__mux4_1 _19249_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net583),
    .S1(net590),
    .X(_07401_));
 sky130_fd_sc_hd__mux4_1 _19250_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net583),
    .S1(net590),
    .X(_07402_));
 sky130_fd_sc_hd__mux4_1 _19251_ (.A0(_07398_),
    .A1(_07400_),
    .A2(_07401_),
    .A3(_07402_),
    .S0(net577),
    .S1(net575),
    .X(_07403_));
 sky130_fd_sc_hd__mux2i_4 _19252_ (.A0(_07397_),
    .A1(_07403_),
    .S(net573),
    .Y(_11756_));
 sky130_fd_sc_hd__mux4_1 _19253_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07404_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1089 ();
 sky130_fd_sc_hd__mux4_1 _19255_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07406_));
 sky130_fd_sc_hd__mux4_1 _19256_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07407_));
 sky130_fd_sc_hd__mux4_1 _19257_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07408_));
 sky130_fd_sc_hd__mux4_4 _19258_ (.A0(_07404_),
    .A1(_07406_),
    .A2(_07407_),
    .A3(_07408_),
    .S0(net577),
    .S1(net575),
    .X(_07409_));
 sky130_fd_sc_hd__mux4_1 _19259_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07410_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1088 ();
 sky130_fd_sc_hd__mux4_1 _19261_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07412_));
 sky130_fd_sc_hd__mux4_1 _19262_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07413_));
 sky130_fd_sc_hd__mux4_1 _19263_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net581),
    .S1(net589),
    .X(_07414_));
 sky130_fd_sc_hd__mux4_1 _19264_ (.A0(_07410_),
    .A1(_07412_),
    .A2(_07413_),
    .A3(_07414_),
    .S0(net577),
    .S1(net575),
    .X(_07415_));
 sky130_fd_sc_hd__mux2i_4 _19265_ (.A0(_07409_),
    .A1(_07415_),
    .S(\count7_1[5] ),
    .Y(_11764_));
 sky130_fd_sc_hd__mux4_1 _19266_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(\count7_1[2] ),
    .S1(net591),
    .X(_07416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1087 ();
 sky130_fd_sc_hd__mux4_1 _19268_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(\count7_1[2] ),
    .S1(\count7_1[1] ),
    .X(_07418_));
 sky130_fd_sc_hd__mux4_1 _19269_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(\count7_1[2] ),
    .S1(net591),
    .X(_07419_));
 sky130_fd_sc_hd__mux4_1 _19270_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(\count7_1[2] ),
    .S1(net591),
    .X(_07420_));
 sky130_fd_sc_hd__mux4_4 _19271_ (.A0(_07416_),
    .A1(_07418_),
    .A2(_07419_),
    .A3(_07420_),
    .S0(net579),
    .S1(net575),
    .X(_07421_));
 sky130_fd_sc_hd__mux4_1 _19272_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net583),
    .S1(net588),
    .X(_07422_));
 sky130_fd_sc_hd__mux4_1 _19273_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net582),
    .S1(net588),
    .X(_07423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1086 ();
 sky130_fd_sc_hd__mux4_1 _19275_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net583),
    .S1(net588),
    .X(_07425_));
 sky130_fd_sc_hd__mux4_1 _19276_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net583),
    .S1(net588),
    .X(_07426_));
 sky130_fd_sc_hd__mux4_1 _19277_ (.A0(_07422_),
    .A1(_07423_),
    .A2(_07425_),
    .A3(_07426_),
    .S0(net577),
    .S1(net575),
    .X(_07427_));
 sky130_fd_sc_hd__mux2i_4 _19278_ (.A0(_07421_),
    .A1(_07427_),
    .S(\count7_1[5] ),
    .Y(_11775_));
 sky130_fd_sc_hd__mux4_1 _19279_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07428_));
 sky130_fd_sc_hd__mux4_1 _19280_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07429_));
 sky130_fd_sc_hd__mux4_1 _19281_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07430_));
 sky130_fd_sc_hd__mux4_1 _19282_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07431_));
 sky130_fd_sc_hd__mux4_4 _19283_ (.A0(_07428_),
    .A1(_07429_),
    .A2(_07430_),
    .A3(_07431_),
    .S0(net579),
    .S1(net575),
    .X(_07432_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1085 ();
 sky130_fd_sc_hd__mux4_1 _19285_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07434_));
 sky130_fd_sc_hd__mux4_1 _19286_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net583),
    .S1(net590),
    .X(_07435_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1084 ();
 sky130_fd_sc_hd__mux4_1 _19288_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07437_));
 sky130_fd_sc_hd__mux4_1 _19289_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07438_));
 sky130_fd_sc_hd__mux4_1 _19290_ (.A0(_07434_),
    .A1(_07435_),
    .A2(_07437_),
    .A3(_07438_),
    .S0(net577),
    .S1(net575),
    .X(_07439_));
 sky130_fd_sc_hd__mux2i_4 _19291_ (.A0(_07432_),
    .A1(_07439_),
    .S(net573),
    .Y(_11783_));
 sky130_fd_sc_hd__mux4_1 _19292_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net580),
    .S1(net591),
    .X(_07440_));
 sky130_fd_sc_hd__mux4_1 _19293_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net580),
    .S1(\count7_1[1] ),
    .X(_07441_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1083 ();
 sky130_fd_sc_hd__mux4_1 _19295_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net580),
    .S1(net591),
    .X(_07443_));
 sky130_fd_sc_hd__mux4_1 _19296_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net580),
    .S1(net591),
    .X(_07444_));
 sky130_fd_sc_hd__mux4_4 _19297_ (.A0(_07440_),
    .A1(_07441_),
    .A2(_07443_),
    .A3(_07444_),
    .S0(net579),
    .S1(net575),
    .X(_07445_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1082 ();
 sky130_fd_sc_hd__mux4_1 _19299_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net583),
    .S1(net589),
    .X(_07447_));
 sky130_fd_sc_hd__mux4_1 _19300_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net583),
    .S1(net589),
    .X(_07448_));
 sky130_fd_sc_hd__mux4_1 _19301_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net580),
    .S1(net589),
    .X(_07449_));
 sky130_fd_sc_hd__mux4_1 _19302_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net583),
    .S1(net589),
    .X(_07450_));
 sky130_fd_sc_hd__mux4_1 _19303_ (.A0(_07447_),
    .A1(_07448_),
    .A2(_07449_),
    .A3(_07450_),
    .S0(net577),
    .S1(net575),
    .X(_07451_));
 sky130_fd_sc_hd__mux2i_4 _19304_ (.A0(_07445_),
    .A1(_07451_),
    .S(net573),
    .Y(_11791_));
 sky130_fd_sc_hd__mux4_1 _19305_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net585),
    .S1(net587),
    .X(_07452_));
 sky130_fd_sc_hd__mux4_1 _19306_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net585),
    .S1(net587),
    .X(_07453_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1081 ();
 sky130_fd_sc_hd__mux4_1 _19308_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net585),
    .S1(net587),
    .X(_07455_));
 sky130_fd_sc_hd__mux4_1 _19309_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net585),
    .S1(net587),
    .X(_07456_));
 sky130_fd_sc_hd__mux4_4 _19310_ (.A0(_07452_),
    .A1(_07453_),
    .A2(_07455_),
    .A3(_07456_),
    .S0(net578),
    .S1(net576),
    .X(_07457_));
 sky130_fd_sc_hd__mux4_1 _19311_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net582),
    .S1(net588),
    .X(_07458_));
 sky130_fd_sc_hd__mux4_1 _19312_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net582),
    .S1(net588),
    .X(_07459_));
 sky130_fd_sc_hd__mux4_1 _19313_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net582),
    .S1(net588),
    .X(_07460_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1080 ();
 sky130_fd_sc_hd__mux4_1 _19315_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net582),
    .S1(net588),
    .X(_07462_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1079 ();
 sky130_fd_sc_hd__mux4_1 _19317_ (.A0(_07458_),
    .A1(_07459_),
    .A2(_07460_),
    .A3(_07462_),
    .S0(net578),
    .S1(net576),
    .X(_07464_));
 sky130_fd_sc_hd__mux2i_4 _19318_ (.A0(_07457_),
    .A1(_07464_),
    .S(net574),
    .Y(_11799_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1078 ();
 sky130_fd_sc_hd__mux4_1 _19320_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net580),
    .S1(net591),
    .X(_07466_));
 sky130_fd_sc_hd__mux4_1 _19321_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net580),
    .S1(\count7_1[1] ),
    .X(_07467_));
 sky130_fd_sc_hd__mux4_1 _19322_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net580),
    .S1(net591),
    .X(_07468_));
 sky130_fd_sc_hd__mux4_1 _19323_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net580),
    .S1(net591),
    .X(_07469_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1077 ();
 sky130_fd_sc_hd__mux4_4 _19325_ (.A0(_07466_),
    .A1(_07467_),
    .A2(_07468_),
    .A3(_07469_),
    .S0(net579),
    .S1(net575),
    .X(_07471_));
 sky130_fd_sc_hd__mux4_1 _19326_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net581),
    .S1(net589),
    .X(_07472_));
 sky130_fd_sc_hd__mux4_1 _19327_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net581),
    .S1(net589),
    .X(_07473_));
 sky130_fd_sc_hd__mux4_1 _19328_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net581),
    .S1(net589),
    .X(_07474_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1076 ();
 sky130_fd_sc_hd__mux4_1 _19330_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net581),
    .S1(net589),
    .X(_07476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1075 ();
 sky130_fd_sc_hd__mux4_1 _19332_ (.A0(_07472_),
    .A1(_07473_),
    .A2(_07474_),
    .A3(_07476_),
    .S0(net577),
    .S1(net575),
    .X(_07478_));
 sky130_fd_sc_hd__mux2i_4 _19333_ (.A0(_07471_),
    .A1(_07478_),
    .S(\count7_1[5] ),
    .Y(_11807_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1074 ();
 sky130_fd_sc_hd__mux4_1 _19335_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net581),
    .S1(net591),
    .X(_07480_));
 sky130_fd_sc_hd__mux4_1 _19336_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net581),
    .S1(net591),
    .X(_07481_));
 sky130_fd_sc_hd__mux4_1 _19337_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net581),
    .S1(net591),
    .X(_07482_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1073 ();
 sky130_fd_sc_hd__mux4_1 _19339_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net581),
    .S1(net591),
    .X(_07484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1072 ();
 sky130_fd_sc_hd__mux4_4 _19341_ (.A0(_07480_),
    .A1(_07481_),
    .A2(_07482_),
    .A3(_07484_),
    .S0(net577),
    .S1(net576),
    .X(_07486_));
 sky130_fd_sc_hd__mux4_1 _19342_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net582),
    .S1(net588),
    .X(_07487_));
 sky130_fd_sc_hd__mux4_1 _19343_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net582),
    .S1(net588),
    .X(_07488_));
 sky130_fd_sc_hd__mux4_1 _19344_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net582),
    .S1(net588),
    .X(_07489_));
 sky130_fd_sc_hd__mux4_1 _19345_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net582),
    .S1(net588),
    .X(_07490_));
 sky130_fd_sc_hd__mux4_1 _19346_ (.A0(_07487_),
    .A1(_07488_),
    .A2(_07489_),
    .A3(_07490_),
    .S0(net577),
    .S1(net575),
    .X(_07491_));
 sky130_fd_sc_hd__mux2i_4 _19347_ (.A0(_07486_),
    .A1(_07491_),
    .S(\count7_1[5] ),
    .Y(_11815_));
 sky130_fd_sc_hd__mux4_1 _19348_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net584),
    .S1(net588),
    .X(_07492_));
 sky130_fd_sc_hd__mux4_1 _19349_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net584),
    .S1(net588),
    .X(_07493_));
 sky130_fd_sc_hd__mux4_1 _19350_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net584),
    .S1(net588),
    .X(_07494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1071 ();
 sky130_fd_sc_hd__mux4_1 _19352_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net584),
    .S1(net588),
    .X(_07496_));
 sky130_fd_sc_hd__mux4_4 _19353_ (.A0(_07492_),
    .A1(_07493_),
    .A2(_07494_),
    .A3(_07496_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07497_));
 sky130_fd_sc_hd__mux4_1 _19354_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net586),
    .S1(net590),
    .X(_07498_));
 sky130_fd_sc_hd__mux4_1 _19355_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net586),
    .S1(net590),
    .X(_07499_));
 sky130_fd_sc_hd__mux4_1 _19356_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net586),
    .S1(net590),
    .X(_07500_));
 sky130_fd_sc_hd__mux4_1 _19357_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net586),
    .S1(net590),
    .X(_07501_));
 sky130_fd_sc_hd__mux4_1 _19358_ (.A0(_07498_),
    .A1(_07499_),
    .A2(_07500_),
    .A3(_07501_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07502_));
 sky130_fd_sc_hd__mux2i_4 _19359_ (.A0(_07497_),
    .A1(_07502_),
    .S(net574),
    .Y(_11823_));
 sky130_fd_sc_hd__mux4_1 _19360_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net584),
    .S1(net588),
    .X(_07503_));
 sky130_fd_sc_hd__mux4_1 _19361_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net584),
    .S1(net588),
    .X(_07504_));
 sky130_fd_sc_hd__mux4_1 _19362_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net584),
    .S1(net588),
    .X(_07505_));
 sky130_fd_sc_hd__mux4_1 _19363_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net584),
    .S1(net588),
    .X(_07506_));
 sky130_fd_sc_hd__mux4_4 _19364_ (.A0(_07503_),
    .A1(_07504_),
    .A2(_07505_),
    .A3(_07506_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07507_));
 sky130_fd_sc_hd__mux4_1 _19365_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net586),
    .S1(net588),
    .X(_07508_));
 sky130_fd_sc_hd__mux4_1 _19366_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net586),
    .S1(net588),
    .X(_07509_));
 sky130_fd_sc_hd__mux4_1 _19367_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net586),
    .S1(net588),
    .X(_07510_));
 sky130_fd_sc_hd__mux4_1 _19368_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net586),
    .S1(net588),
    .X(_07511_));
 sky130_fd_sc_hd__mux4_1 _19369_ (.A0(_07508_),
    .A1(_07509_),
    .A2(_07510_),
    .A3(_07511_),
    .S0(net578),
    .S1(net576),
    .X(_07512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1070 ();
 sky130_fd_sc_hd__mux2i_4 _19371_ (.A0(_07507_),
    .A1(_07512_),
    .S(net574),
    .Y(_11831_));
 sky130_fd_sc_hd__mux4_1 _19372_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net584),
    .S1(net588),
    .X(_07514_));
 sky130_fd_sc_hd__mux4_1 _19373_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net584),
    .S1(net588),
    .X(_07515_));
 sky130_fd_sc_hd__mux4_1 _19374_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net584),
    .S1(net588),
    .X(_07516_));
 sky130_fd_sc_hd__mux4_1 _19375_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net584),
    .S1(net588),
    .X(_07517_));
 sky130_fd_sc_hd__mux4_4 _19376_ (.A0(_07514_),
    .A1(_07515_),
    .A2(_07516_),
    .A3(_07517_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07518_));
 sky130_fd_sc_hd__mux4_1 _19377_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net586),
    .S1(net590),
    .X(_07519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1069 ();
 sky130_fd_sc_hd__mux4_1 _19379_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net586),
    .S1(net590),
    .X(_07521_));
 sky130_fd_sc_hd__mux4_1 _19380_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net586),
    .S1(net590),
    .X(_07522_));
 sky130_fd_sc_hd__mux4_1 _19381_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net586),
    .S1(net590),
    .X(_07523_));
 sky130_fd_sc_hd__mux4_2 _19382_ (.A0(_07519_),
    .A1(_07521_),
    .A2(_07522_),
    .A3(_07523_),
    .S0(net578),
    .S1(net576),
    .X(_07524_));
 sky130_fd_sc_hd__mux2i_4 _19383_ (.A0(_07518_),
    .A1(_07524_),
    .S(net574),
    .Y(_11839_));
 sky130_fd_sc_hd__mux4_1 _19384_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net580),
    .S1(net591),
    .X(_07525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1068 ();
 sky130_fd_sc_hd__mux4_1 _19386_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net580),
    .S1(\count7_1[1] ),
    .X(_07527_));
 sky130_fd_sc_hd__mux4_1 _19387_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net580),
    .S1(net591),
    .X(_07528_));
 sky130_fd_sc_hd__mux4_1 _19388_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net580),
    .S1(net591),
    .X(_07529_));
 sky130_fd_sc_hd__mux4_4 _19389_ (.A0(_07525_),
    .A1(_07527_),
    .A2(_07528_),
    .A3(_07529_),
    .S0(net579),
    .S1(net575),
    .X(_07530_));
 sky130_fd_sc_hd__mux4_1 _19390_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net582),
    .S1(net588),
    .X(_07531_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1067 ();
 sky130_fd_sc_hd__mux4_1 _19392_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net581),
    .S1(net588),
    .X(_07533_));
 sky130_fd_sc_hd__mux4_1 _19393_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net581),
    .S1(net588),
    .X(_07534_));
 sky130_fd_sc_hd__mux4_1 _19394_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net583),
    .S1(net588),
    .X(_07535_));
 sky130_fd_sc_hd__mux4_2 _19395_ (.A0(_07531_),
    .A1(_07533_),
    .A2(_07534_),
    .A3(_07535_),
    .S0(net577),
    .S1(net575),
    .X(_07536_));
 sky130_fd_sc_hd__mux2i_4 _19396_ (.A0(_07530_),
    .A1(_07536_),
    .S(\count7_1[5] ),
    .Y(_11847_));
 sky130_fd_sc_hd__mux4_1 _19397_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net584),
    .S1(net588),
    .X(_07537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1066 ();
 sky130_fd_sc_hd__mux4_1 _19399_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net584),
    .S1(net588),
    .X(_07539_));
 sky130_fd_sc_hd__mux4_1 _19400_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net584),
    .S1(net588),
    .X(_07540_));
 sky130_fd_sc_hd__mux4_1 _19401_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net584),
    .S1(net588),
    .X(_07541_));
 sky130_fd_sc_hd__mux4_4 _19402_ (.A0(_07537_),
    .A1(_07539_),
    .A2(_07540_),
    .A3(_07541_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07542_));
 sky130_fd_sc_hd__mux4_1 _19403_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net586),
    .S1(net590),
    .X(_07543_));
 sky130_fd_sc_hd__mux4_1 _19404_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net584),
    .S1(net590),
    .X(_07544_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1065 ();
 sky130_fd_sc_hd__mux4_1 _19406_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net586),
    .S1(net590),
    .X(_07546_));
 sky130_fd_sc_hd__mux4_1 _19407_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net586),
    .S1(net590),
    .X(_07547_));
 sky130_fd_sc_hd__mux4_1 _19408_ (.A0(_07543_),
    .A1(_07544_),
    .A2(_07546_),
    .A3(_07547_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07548_));
 sky130_fd_sc_hd__mux2i_4 _19409_ (.A0(_07542_),
    .A1(_07548_),
    .S(net574),
    .Y(_11855_));
 sky130_fd_sc_hd__mux4_1 _19410_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net580),
    .S1(net591),
    .X(_07549_));
 sky130_fd_sc_hd__mux4_1 _19411_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net580),
    .S1(net591),
    .X(_07550_));
 sky130_fd_sc_hd__mux4_1 _19412_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net580),
    .S1(net591),
    .X(_07551_));
 sky130_fd_sc_hd__mux4_1 _19413_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net580),
    .S1(net591),
    .X(_07552_));
 sky130_fd_sc_hd__mux4_4 _19414_ (.A0(_07549_),
    .A1(_07550_),
    .A2(_07551_),
    .A3(_07552_),
    .S0(net579),
    .S1(net575),
    .X(_07553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1064 ();
 sky130_fd_sc_hd__mux4_1 _19416_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net583),
    .S1(net589),
    .X(_07555_));
 sky130_fd_sc_hd__mux4_1 _19417_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net583),
    .S1(net589),
    .X(_07556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1063 ();
 sky130_fd_sc_hd__mux4_1 _19419_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net583),
    .S1(net589),
    .X(_07558_));
 sky130_fd_sc_hd__mux4_1 _19420_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net583),
    .S1(net589),
    .X(_07559_));
 sky130_fd_sc_hd__mux4_1 _19421_ (.A0(_07555_),
    .A1(_07556_),
    .A2(_07558_),
    .A3(_07559_),
    .S0(net577),
    .S1(net575),
    .X(_07560_));
 sky130_fd_sc_hd__mux2i_4 _19422_ (.A0(_07553_),
    .A1(_07560_),
    .S(net573),
    .Y(_11863_));
 sky130_fd_sc_hd__mux4_1 _19423_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net580),
    .S1(net591),
    .X(_07561_));
 sky130_fd_sc_hd__mux4_1 _19424_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net580),
    .S1(\count7_1[1] ),
    .X(_07562_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1062 ();
 sky130_fd_sc_hd__mux4_1 _19426_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net580),
    .S1(net591),
    .X(_07564_));
 sky130_fd_sc_hd__mux4_1 _19427_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net580),
    .S1(net591),
    .X(_07565_));
 sky130_fd_sc_hd__mux4_4 _19428_ (.A0(_07561_),
    .A1(_07562_),
    .A2(_07564_),
    .A3(_07565_),
    .S0(net579),
    .S1(net575),
    .X(_07566_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1061 ();
 sky130_fd_sc_hd__mux4_1 _19430_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net583),
    .S1(net589),
    .X(_07568_));
 sky130_fd_sc_hd__mux4_1 _19431_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net583),
    .S1(net589),
    .X(_07569_));
 sky130_fd_sc_hd__mux4_1 _19432_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net583),
    .S1(net589),
    .X(_07570_));
 sky130_fd_sc_hd__mux4_1 _19433_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net583),
    .S1(net589),
    .X(_07571_));
 sky130_fd_sc_hd__mux4_1 _19434_ (.A0(_07568_),
    .A1(_07569_),
    .A2(_07570_),
    .A3(_07571_),
    .S0(net577),
    .S1(net575),
    .X(_07572_));
 sky130_fd_sc_hd__mux2i_4 _19435_ (.A0(_07566_),
    .A1(_07572_),
    .S(net573),
    .Y(_11871_));
 sky130_fd_sc_hd__mux4_1 _19436_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net580),
    .S1(net591),
    .X(_07573_));
 sky130_fd_sc_hd__mux4_1 _19437_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net580),
    .S1(\count7_1[1] ),
    .X(_07574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1060 ();
 sky130_fd_sc_hd__mux4_1 _19439_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net580),
    .S1(net591),
    .X(_07576_));
 sky130_fd_sc_hd__mux4_1 _19440_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net580),
    .S1(net591),
    .X(_07577_));
 sky130_fd_sc_hd__mux4_2 _19441_ (.A0(_07573_),
    .A1(_07574_),
    .A2(_07576_),
    .A3(_07577_),
    .S0(net579),
    .S1(net575),
    .X(_07578_));
 sky130_fd_sc_hd__mux4_1 _19442_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net583),
    .S1(net589),
    .X(_07579_));
 sky130_fd_sc_hd__mux4_1 _19443_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net583),
    .S1(net589),
    .X(_07580_));
 sky130_fd_sc_hd__mux4_1 _19444_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net583),
    .S1(net589),
    .X(_07581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1059 ();
 sky130_fd_sc_hd__mux4_1 _19446_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net583),
    .S1(net589),
    .X(_07583_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1058 ();
 sky130_fd_sc_hd__mux4_1 _19448_ (.A0(_07579_),
    .A1(_07580_),
    .A2(_07581_),
    .A3(_07583_),
    .S0(net577),
    .S1(net575),
    .X(_07585_));
 sky130_fd_sc_hd__mux2i_4 _19449_ (.A0(_07578_),
    .A1(_07585_),
    .S(net573),
    .Y(_11879_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1057 ();
 sky130_fd_sc_hd__mux4_1 _19451_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net580),
    .S1(net591),
    .X(_07587_));
 sky130_fd_sc_hd__mux4_1 _19452_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net580),
    .S1(net591),
    .X(_07588_));
 sky130_fd_sc_hd__mux4_1 _19453_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net580),
    .S1(net591),
    .X(_07589_));
 sky130_fd_sc_hd__mux4_1 _19454_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net580),
    .S1(net591),
    .X(_07590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1056 ();
 sky130_fd_sc_hd__mux4_4 _19456_ (.A0(_07587_),
    .A1(_07588_),
    .A2(_07589_),
    .A3(_07590_),
    .S0(net579),
    .S1(net575),
    .X(_07592_));
 sky130_fd_sc_hd__mux4_1 _19457_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net583),
    .S1(net591),
    .X(_07593_));
 sky130_fd_sc_hd__mux4_1 _19458_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net583),
    .S1(net591),
    .X(_07594_));
 sky130_fd_sc_hd__mux4_1 _19459_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net583),
    .S1(net591),
    .X(_07595_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1055 ();
 sky130_fd_sc_hd__mux4_1 _19461_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net583),
    .S1(net591),
    .X(_07597_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1054 ();
 sky130_fd_sc_hd__mux4_1 _19463_ (.A0(_07593_),
    .A1(_07594_),
    .A2(_07595_),
    .A3(_07597_),
    .S0(net577),
    .S1(net575),
    .X(_07599_));
 sky130_fd_sc_hd__mux2i_4 _19464_ (.A0(_07592_),
    .A1(_07599_),
    .S(net573),
    .Y(_11887_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1053 ();
 sky130_fd_sc_hd__mux4_1 _19466_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net585),
    .S1(net587),
    .X(_07601_));
 sky130_fd_sc_hd__mux4_1 _19467_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net585),
    .S1(net587),
    .X(_07602_));
 sky130_fd_sc_hd__mux4_1 _19468_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net585),
    .S1(net587),
    .X(_07603_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1052 ();
 sky130_fd_sc_hd__mux4_1 _19470_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net585),
    .S1(net587),
    .X(_07605_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1051 ();
 sky130_fd_sc_hd__mux4_4 _19472_ (.A0(_07601_),
    .A1(_07602_),
    .A2(_07603_),
    .A3(_07605_),
    .S0(net578),
    .S1(net576),
    .X(_07607_));
 sky130_fd_sc_hd__mux4_1 _19473_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net585),
    .S1(net588),
    .X(_07608_));
 sky130_fd_sc_hd__mux4_1 _19474_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net585),
    .S1(net588),
    .X(_07609_));
 sky130_fd_sc_hd__mux4_1 _19475_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net585),
    .S1(net588),
    .X(_07610_));
 sky130_fd_sc_hd__mux4_1 _19476_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net585),
    .S1(net588),
    .X(_07611_));
 sky130_fd_sc_hd__mux4_1 _19477_ (.A0(_07608_),
    .A1(_07609_),
    .A2(_07610_),
    .A3(_07611_),
    .S0(net578),
    .S1(net576),
    .X(_07612_));
 sky130_fd_sc_hd__mux2i_4 _19478_ (.A0(_07607_),
    .A1(_07612_),
    .S(net574),
    .Y(_11895_));
 sky130_fd_sc_hd__mux4_1 _19479_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net586),
    .S1(net587),
    .X(_07613_));
 sky130_fd_sc_hd__mux4_1 _19480_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net586),
    .S1(net587),
    .X(_07614_));
 sky130_fd_sc_hd__mux4_1 _19481_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net586),
    .S1(net587),
    .X(_07615_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1050 ();
 sky130_fd_sc_hd__mux4_1 _19483_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net586),
    .S1(net587),
    .X(_07617_));
 sky130_fd_sc_hd__mux4_4 _19484_ (.A0(_07613_),
    .A1(_07614_),
    .A2(_07615_),
    .A3(_07617_),
    .S0(net578),
    .S1(net576),
    .X(_07618_));
 sky130_fd_sc_hd__mux4_1 _19485_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07619_));
 sky130_fd_sc_hd__mux4_1 _19486_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net586),
    .S1(net590),
    .X(_07620_));
 sky130_fd_sc_hd__mux4_1 _19487_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net586),
    .S1(net590),
    .X(_07621_));
 sky130_fd_sc_hd__mux4_1 _19488_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net586),
    .S1(net590),
    .X(_07622_));
 sky130_fd_sc_hd__mux4_1 _19489_ (.A0(_07619_),
    .A1(_07620_),
    .A2(_07621_),
    .A3(_07622_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07623_));
 sky130_fd_sc_hd__mux2i_4 _19490_ (.A0(_07618_),
    .A1(_07623_),
    .S(net574),
    .Y(_11903_));
 sky130_fd_sc_hd__mux4_1 _19491_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07624_));
 sky130_fd_sc_hd__mux4_1 _19492_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07625_));
 sky130_fd_sc_hd__mux4_1 _19493_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07626_));
 sky130_fd_sc_hd__mux4_1 _19494_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07627_));
 sky130_fd_sc_hd__mux4_2 _19495_ (.A0(_07624_),
    .A1(_07625_),
    .A2(_07626_),
    .A3(_07627_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07628_));
 sky130_fd_sc_hd__mux4_1 _19496_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07629_));
 sky130_fd_sc_hd__mux4_1 _19497_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07630_));
 sky130_fd_sc_hd__mux4_1 _19498_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07631_));
 sky130_fd_sc_hd__mux4_1 _19499_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(\count7_1[2] ),
    .S1(net590),
    .X(_07632_));
 sky130_fd_sc_hd__mux4_1 _19500_ (.A0(_07629_),
    .A1(_07630_),
    .A2(_07631_),
    .A3(_07632_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07633_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1049 ();
 sky130_fd_sc_hd__mux2i_4 _19502_ (.A0(_07628_),
    .A1(_07633_),
    .S(net574),
    .Y(_11911_));
 sky130_fd_sc_hd__mux4_1 _19503_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net586),
    .S1(net587),
    .X(_07635_));
 sky130_fd_sc_hd__mux4_1 _19504_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net586),
    .S1(net587),
    .X(_07636_));
 sky130_fd_sc_hd__mux4_1 _19505_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net586),
    .S1(net587),
    .X(_07637_));
 sky130_fd_sc_hd__mux4_1 _19506_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net586),
    .S1(net587),
    .X(_07638_));
 sky130_fd_sc_hd__mux4_4 _19507_ (.A0(_07635_),
    .A1(_07636_),
    .A2(_07637_),
    .A3(_07638_),
    .S0(net578),
    .S1(net576),
    .X(_07639_));
 sky130_fd_sc_hd__mux4_1 _19508_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net585),
    .S1(net590),
    .X(_07640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1048 ();
 sky130_fd_sc_hd__mux4_1 _19510_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net585),
    .S1(net590),
    .X(_07642_));
 sky130_fd_sc_hd__mux4_1 _19511_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net585),
    .S1(net590),
    .X(_07643_));
 sky130_fd_sc_hd__mux4_1 _19512_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net585),
    .S1(net590),
    .X(_07644_));
 sky130_fd_sc_hd__mux4_1 _19513_ (.A0(_07640_),
    .A1(_07642_),
    .A2(_07643_),
    .A3(_07644_),
    .S0(net578),
    .S1(net576),
    .X(_07645_));
 sky130_fd_sc_hd__mux2i_4 _19514_ (.A0(_07639_),
    .A1(_07645_),
    .S(net574),
    .Y(_11919_));
 sky130_fd_sc_hd__mux4_1 _19515_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net584),
    .S1(net588),
    .X(_07646_));
 sky130_fd_sc_hd__mux4_1 _19516_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net584),
    .S1(net588),
    .X(_07647_));
 sky130_fd_sc_hd__mux4_1 _19517_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net584),
    .S1(net588),
    .X(_07648_));
 sky130_fd_sc_hd__mux4_1 _19518_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net584),
    .S1(net588),
    .X(_07649_));
 sky130_fd_sc_hd__mux4_4 _19519_ (.A0(_07646_),
    .A1(_07647_),
    .A2(_07648_),
    .A3(_07649_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07650_));
 sky130_fd_sc_hd__mux4_1 _19520_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net586),
    .S1(net588),
    .X(_07651_));
 sky130_fd_sc_hd__mux4_1 _19521_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net586),
    .S1(net588),
    .X(_07652_));
 sky130_fd_sc_hd__mux4_1 _19522_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net586),
    .S1(net588),
    .X(_07653_));
 sky130_fd_sc_hd__mux4_1 _19523_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net586),
    .S1(net588),
    .X(_07654_));
 sky130_fd_sc_hd__mux4_1 _19524_ (.A0(_07651_),
    .A1(_07652_),
    .A2(_07653_),
    .A3(_07654_),
    .S0(net578),
    .S1(net576),
    .X(_07655_));
 sky130_fd_sc_hd__mux2i_4 _19525_ (.A0(_07650_),
    .A1(_07655_),
    .S(net574),
    .Y(_11927_));
 sky130_fd_sc_hd__mux4_1 _19526_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net582),
    .S1(net589),
    .X(_07656_));
 sky130_fd_sc_hd__mux4_1 _19527_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net581),
    .S1(net591),
    .X(_07657_));
 sky130_fd_sc_hd__mux4_1 _19528_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net582),
    .S1(net589),
    .X(_07658_));
 sky130_fd_sc_hd__mux4_1 _19529_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net582),
    .S1(net589),
    .X(_07659_));
 sky130_fd_sc_hd__mux4_4 _19530_ (.A0(_07656_),
    .A1(_07657_),
    .A2(_07658_),
    .A3(_07659_),
    .S0(net578),
    .S1(net576),
    .X(_07660_));
 sky130_fd_sc_hd__mux4_1 _19531_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net582),
    .S1(net587),
    .X(_07661_));
 sky130_fd_sc_hd__mux4_1 _19532_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net582),
    .S1(net587),
    .X(_07662_));
 sky130_fd_sc_hd__mux4_1 _19533_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net582),
    .S1(net587),
    .X(_07663_));
 sky130_fd_sc_hd__mux4_1 _19534_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net582),
    .S1(net587),
    .X(_07664_));
 sky130_fd_sc_hd__mux4_1 _19535_ (.A0(_07661_),
    .A1(_07662_),
    .A2(_07663_),
    .A3(_07664_),
    .S0(net578),
    .S1(net576),
    .X(_07665_));
 sky130_fd_sc_hd__mux2i_4 _19536_ (.A0(_07660_),
    .A1(_07665_),
    .S(net574),
    .Y(_11935_));
 sky130_fd_sc_hd__mux4_1 _19537_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net580),
    .S1(net591),
    .X(_07666_));
 sky130_fd_sc_hd__mux4_1 _19538_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net580),
    .S1(net591),
    .X(_07667_));
 sky130_fd_sc_hd__mux4_1 _19539_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net580),
    .S1(net591),
    .X(_07668_));
 sky130_fd_sc_hd__mux4_1 _19540_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net580),
    .S1(net591),
    .X(_07669_));
 sky130_fd_sc_hd__mux4_4 _19541_ (.A0(_07666_),
    .A1(_07667_),
    .A2(_07668_),
    .A3(_07669_),
    .S0(net577),
    .S1(net575),
    .X(_07670_));
 sky130_fd_sc_hd__mux4_1 _19542_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net581),
    .S1(net591),
    .X(_07671_));
 sky130_fd_sc_hd__mux4_1 _19543_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net581),
    .S1(net591),
    .X(_07672_));
 sky130_fd_sc_hd__mux4_1 _19544_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net581),
    .S1(net591),
    .X(_07673_));
 sky130_fd_sc_hd__mux4_1 _19545_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net581),
    .S1(net591),
    .X(_07674_));
 sky130_fd_sc_hd__mux4_1 _19546_ (.A0(_07671_),
    .A1(_07672_),
    .A2(_07673_),
    .A3(_07674_),
    .S0(net577),
    .S1(net575),
    .X(_07675_));
 sky130_fd_sc_hd__mux2i_4 _19547_ (.A0(_07670_),
    .A1(_07675_),
    .S(net573),
    .Y(_11943_));
 sky130_fd_sc_hd__mux4_1 _19548_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net581),
    .S1(net591),
    .X(_07676_));
 sky130_fd_sc_hd__mux4_1 _19549_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net581),
    .S1(net591),
    .X(_07677_));
 sky130_fd_sc_hd__mux4_1 _19550_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net581),
    .S1(net591),
    .X(_07678_));
 sky130_fd_sc_hd__mux4_1 _19551_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net581),
    .S1(net591),
    .X(_07679_));
 sky130_fd_sc_hd__mux4_4 _19552_ (.A0(_07676_),
    .A1(_07677_),
    .A2(_07678_),
    .A3(_07679_),
    .S0(net577),
    .S1(net575),
    .X(_07680_));
 sky130_fd_sc_hd__mux4_1 _19553_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net581),
    .S1(net589),
    .X(_07681_));
 sky130_fd_sc_hd__mux4_1 _19554_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net581),
    .S1(net589),
    .X(_07682_));
 sky130_fd_sc_hd__mux4_1 _19555_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net581),
    .S1(net589),
    .X(_07683_));
 sky130_fd_sc_hd__mux4_1 _19556_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net581),
    .S1(net589),
    .X(_07684_));
 sky130_fd_sc_hd__mux4_1 _19557_ (.A0(_07681_),
    .A1(_07682_),
    .A2(_07683_),
    .A3(_07684_),
    .S0(net577),
    .S1(net575),
    .X(_07685_));
 sky130_fd_sc_hd__mux2i_4 _19558_ (.A0(_07680_),
    .A1(_07685_),
    .S(\count7_1[5] ),
    .Y(_11951_));
 sky130_fd_sc_hd__mux4_1 _19559_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net581),
    .S1(net591),
    .X(_07686_));
 sky130_fd_sc_hd__mux4_1 _19560_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net581),
    .S1(net591),
    .X(_07687_));
 sky130_fd_sc_hd__mux4_1 _19561_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net581),
    .S1(net591),
    .X(_07688_));
 sky130_fd_sc_hd__mux4_1 _19562_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net581),
    .S1(net591),
    .X(_07689_));
 sky130_fd_sc_hd__mux4_4 _19563_ (.A0(_07686_),
    .A1(_07687_),
    .A2(_07688_),
    .A3(_07689_),
    .S0(net577),
    .S1(net576),
    .X(_07690_));
 sky130_fd_sc_hd__mux4_1 _19564_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net582),
    .S1(net589),
    .X(_07691_));
 sky130_fd_sc_hd__mux4_1 _19565_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net582),
    .S1(net589),
    .X(_07692_));
 sky130_fd_sc_hd__mux4_1 _19566_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net582),
    .S1(net589),
    .X(_07693_));
 sky130_fd_sc_hd__mux4_1 _19567_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net582),
    .S1(net589),
    .X(_07694_));
 sky130_fd_sc_hd__mux4_1 _19568_ (.A0(_07691_),
    .A1(_07692_),
    .A2(_07693_),
    .A3(_07694_),
    .S0(net577),
    .S1(net576),
    .X(_07695_));
 sky130_fd_sc_hd__mux2i_4 _19569_ (.A0(_07690_),
    .A1(_07695_),
    .S(\count7_1[5] ),
    .Y(_11959_));
 sky130_fd_sc_hd__mux4_1 _19570_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net581),
    .S1(net591),
    .X(_07696_));
 sky130_fd_sc_hd__mux4_1 _19571_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net581),
    .S1(net591),
    .X(_07697_));
 sky130_fd_sc_hd__mux4_1 _19572_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net581),
    .S1(net591),
    .X(_07698_));
 sky130_fd_sc_hd__mux4_1 _19573_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net581),
    .S1(net591),
    .X(_07699_));
 sky130_fd_sc_hd__mux4_4 _19574_ (.A0(_07696_),
    .A1(_07697_),
    .A2(_07698_),
    .A3(_07699_),
    .S0(net577),
    .S1(net576),
    .X(_07700_));
 sky130_fd_sc_hd__mux4_1 _19575_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net582),
    .S1(net589),
    .X(_07701_));
 sky130_fd_sc_hd__mux4_1 _19576_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net582),
    .S1(net589),
    .X(_07702_));
 sky130_fd_sc_hd__mux4_1 _19577_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net582),
    .S1(net589),
    .X(_07703_));
 sky130_fd_sc_hd__mux4_1 _19578_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net582),
    .S1(net589),
    .X(_07704_));
 sky130_fd_sc_hd__mux4_1 _19579_ (.A0(_07701_),
    .A1(_07702_),
    .A2(_07703_),
    .A3(_07704_),
    .S0(net577),
    .S1(net576),
    .X(_07705_));
 sky130_fd_sc_hd__mux2i_4 _19580_ (.A0(_07700_),
    .A1(_07705_),
    .S(\count7_1[5] ),
    .Y(_11967_));
 sky130_fd_sc_hd__mux4_1 _19581_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net585),
    .S1(net589),
    .X(_07706_));
 sky130_fd_sc_hd__mux4_1 _19582_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net585),
    .S1(net589),
    .X(_07707_));
 sky130_fd_sc_hd__mux4_1 _19583_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net585),
    .S1(net589),
    .X(_07708_));
 sky130_fd_sc_hd__mux4_1 _19584_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net585),
    .S1(net589),
    .X(_07709_));
 sky130_fd_sc_hd__mux4_4 _19585_ (.A0(_07706_),
    .A1(_07707_),
    .A2(_07708_),
    .A3(_07709_),
    .S0(net578),
    .S1(net576),
    .X(_07710_));
 sky130_fd_sc_hd__mux4_1 _19586_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net585),
    .S1(net587),
    .X(_07711_));
 sky130_fd_sc_hd__mux4_1 _19587_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net585),
    .S1(net587),
    .X(_07712_));
 sky130_fd_sc_hd__mux4_1 _19588_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net585),
    .S1(net587),
    .X(_07713_));
 sky130_fd_sc_hd__mux4_1 _19589_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net585),
    .S1(net587),
    .X(_07714_));
 sky130_fd_sc_hd__mux4_1 _19590_ (.A0(_07711_),
    .A1(_07712_),
    .A2(_07713_),
    .A3(_07714_),
    .S0(net578),
    .S1(net576),
    .X(_07715_));
 sky130_fd_sc_hd__mux2i_4 _19591_ (.A0(_07710_),
    .A1(_07715_),
    .S(net574),
    .Y(_11975_));
 sky130_fd_sc_hd__mux4_1 _19592_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net584),
    .S1(net588),
    .X(_07716_));
 sky130_fd_sc_hd__mux4_1 _19593_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net584),
    .S1(net588),
    .X(_07717_));
 sky130_fd_sc_hd__mux4_1 _19594_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net584),
    .S1(net588),
    .X(_07718_));
 sky130_fd_sc_hd__mux4_1 _19595_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net584),
    .S1(net588),
    .X(_07719_));
 sky130_fd_sc_hd__mux4_4 _19596_ (.A0(_07716_),
    .A1(_07717_),
    .A2(_07718_),
    .A3(_07719_),
    .S0(\count7_1[3] ),
    .S1(\count7_1[4] ),
    .X(_07720_));
 sky130_fd_sc_hd__mux4_1 _19597_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net586),
    .S1(net587),
    .X(_07721_));
 sky130_fd_sc_hd__mux4_1 _19598_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net586),
    .S1(net587),
    .X(_07722_));
 sky130_fd_sc_hd__mux4_1 _19599_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net586),
    .S1(net587),
    .X(_07723_));
 sky130_fd_sc_hd__mux4_1 _19600_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net586),
    .S1(net587),
    .X(_07724_));
 sky130_fd_sc_hd__mux4_1 _19601_ (.A0(_07721_),
    .A1(_07722_),
    .A2(_07723_),
    .A3(_07724_),
    .S0(net578),
    .S1(net576),
    .X(_07725_));
 sky130_fd_sc_hd__mux2i_4 _19602_ (.A0(_07720_),
    .A1(_07725_),
    .S(net574),
    .Y(_11983_));
 sky130_fd_sc_hd__mux4_1 _19603_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07726_));
 sky130_fd_sc_hd__mux4_1 _19604_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07727_));
 sky130_fd_sc_hd__mux4_1 _19605_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07728_));
 sky130_fd_sc_hd__mux4_1 _19606_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07729_));
 sky130_fd_sc_hd__mux4_2 _19607_ (.A0(_07726_),
    .A1(_07727_),
    .A2(_07728_),
    .A3(_07729_),
    .S0(net578),
    .S1(net576),
    .X(_07730_));
 sky130_fd_sc_hd__mux4_1 _19608_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07731_));
 sky130_fd_sc_hd__mux4_1 _19609_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07732_));
 sky130_fd_sc_hd__mux4_1 _19610_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07733_));
 sky130_fd_sc_hd__mux4_1 _19611_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net585),
    .S1(net587),
    .X(_07734_));
 sky130_fd_sc_hd__mux4_1 _19612_ (.A0(_07731_),
    .A1(_07732_),
    .A2(_07733_),
    .A3(_07734_),
    .S0(net578),
    .S1(net576),
    .X(_07735_));
 sky130_fd_sc_hd__mux2i_4 _19613_ (.A0(_07730_),
    .A1(_07735_),
    .S(net574),
    .Y(_11991_));
 sky130_fd_sc_hd__inv_1 _19614_ (.A(\hash.CA1.w_i2[1] ),
    .Y(_12538_));
 sky130_fd_sc_hd__inv_1 _19615_ (.A(\hash.CA1.w_i2[0] ),
    .Y(_12543_));
 sky130_fd_sc_hd__inv_1 _19616_ (.A(\hash.CA1.w_i2[3] ),
    .Y(_12553_));
 sky130_fd_sc_hd__inv_1 _19617_ (.A(\hash.CA1.w_i2[5] ),
    .Y(_12561_));
 sky130_fd_sc_hd__inv_1 _19618_ (.A(\hash.CA1.w_i2[7] ),
    .Y(_12569_));
 sky130_fd_sc_hd__inv_1 _19619_ (.A(\hash.CA1.w_i2[8] ),
    .Y(_12574_));
 sky130_fd_sc_hd__inv_1 _19620_ (.A(\hash.CA1.w_i2[11] ),
    .Y(_12585_));
 sky130_fd_sc_hd__inv_1 _19621_ (.A(\hash.CA1.w_i2[12] ),
    .Y(_12590_));
 sky130_fd_sc_hd__inv_1 _19622_ (.A(\hash.CA1.w_i2[14] ),
    .Y(_12598_));
 sky130_fd_sc_hd__inv_1 _19623_ (.A(\hash.CA1.w_i2[15] ),
    .Y(_12603_));
 sky130_fd_sc_hd__inv_1 _19624_ (.A(\hash.CA1.w_i2[16] ),
    .Y(_12608_));
 sky130_fd_sc_hd__inv_1 _19625_ (.A(\hash.CA1.w_i2[17] ),
    .Y(_12613_));
 sky130_fd_sc_hd__inv_1 _19626_ (.A(\hash.CA1.w_i2[23] ),
    .Y(_12633_));
 sky130_fd_sc_hd__inv_1 _19627_ (.A(\hash.CA1.w_i2[24] ),
    .Y(_12638_));
 sky130_fd_sc_hd__inv_1 _19628_ (.A(\hash.CA1.w_i2[25] ),
    .Y(_12643_));
 sky130_fd_sc_hd__inv_1 _19629_ (.A(\hash.CA1.w_i2[26] ),
    .Y(_12648_));
 sky130_fd_sc_hd__inv_1 _19630_ (.A(\hash.CA1.w_i2[27] ),
    .Y(_12653_));
 sky130_fd_sc_hd__inv_1 _19631_ (.A(\hash.CA1.w_i2[28] ),
    .Y(_12658_));
 sky130_fd_sc_hd__inv_1 _19632_ (.A(_13066_),
    .Y(_13063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1044 ();
 sky130_fd_sc_hd__mux4_1 _19637_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1040 ();
 sky130_fd_sc_hd__mux4_1 _19642_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07745_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1038 ();
 sky130_fd_sc_hd__mux4_1 _19645_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07748_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1035 ();
 sky130_fd_sc_hd__mux4_1 _19649_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07752_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1031 ();
 sky130_fd_sc_hd__mux4_4 _19654_ (.A0(_07740_),
    .A1(_07745_),
    .A2(_07748_),
    .A3(_07752_),
    .S0(net652),
    .S1(net650),
    .X(_07757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1029 ();
 sky130_fd_sc_hd__mux4_1 _19657_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1027 ();
 sky130_fd_sc_hd__mux4_1 _19660_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07763_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1025 ();
 sky130_fd_sc_hd__mux4_1 _19663_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1023 ();
 sky130_fd_sc_hd__mux4_1 _19666_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net656),
    .S1(net660),
    .X(_07769_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1021 ();
 sky130_fd_sc_hd__mux4_1 _19669_ (.A0(_07760_),
    .A1(_07763_),
    .A2(_07766_),
    .A3(_07769_),
    .S0(net652),
    .S1(net650),
    .X(_07772_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1020 ();
 sky130_fd_sc_hd__mux2i_4 _19671_ (.A0(_07757_),
    .A1(_07772_),
    .S(net649),
    .Y(_11752_));
 sky130_fd_sc_hd__mux4_1 _19672_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net656),
    .S1(net660),
    .X(_07774_));
 sky130_fd_sc_hd__mux4_1 _19673_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net656),
    .S1(net660),
    .X(_07775_));
 sky130_fd_sc_hd__mux4_1 _19674_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net656),
    .S1(net660),
    .X(_07776_));
 sky130_fd_sc_hd__mux4_1 _19675_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net656),
    .S1(net660),
    .X(_07777_));
 sky130_fd_sc_hd__mux4_4 _19676_ (.A0(_07774_),
    .A1(_07775_),
    .A2(_07776_),
    .A3(_07777_),
    .S0(net652),
    .S1(net650),
    .X(_07778_));
 sky130_fd_sc_hd__mux4_1 _19677_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net658),
    .S1(net662),
    .X(_07779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1019 ();
 sky130_fd_sc_hd__mux4_1 _19679_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net658),
    .S1(net662),
    .X(_07781_));
 sky130_fd_sc_hd__mux4_1 _19680_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net658),
    .S1(net662),
    .X(_07782_));
 sky130_fd_sc_hd__mux4_1 _19681_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net658),
    .S1(net662),
    .X(_07783_));
 sky130_fd_sc_hd__mux4_1 _19682_ (.A0(_07779_),
    .A1(_07781_),
    .A2(_07782_),
    .A3(_07783_),
    .S0(net652),
    .S1(net650),
    .X(_07784_));
 sky130_fd_sc_hd__mux2i_4 _19683_ (.A0(_07778_),
    .A1(_07784_),
    .S(net649),
    .Y(_11757_));
 sky130_fd_sc_hd__mux4_1 _19684_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net656),
    .S1(net660),
    .X(_07785_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1018 ();
 sky130_fd_sc_hd__mux4_1 _19686_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net656),
    .S1(net660),
    .X(_07787_));
 sky130_fd_sc_hd__mux4_1 _19687_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net656),
    .S1(net660),
    .X(_07788_));
 sky130_fd_sc_hd__mux4_1 _19688_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net656),
    .S1(net660),
    .X(_07789_));
 sky130_fd_sc_hd__mux4_4 _19689_ (.A0(_07785_),
    .A1(_07787_),
    .A2(_07788_),
    .A3(_07789_),
    .S0(net652),
    .S1(net650),
    .X(_07790_));
 sky130_fd_sc_hd__mux4_1 _19690_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net658),
    .S1(net661),
    .X(_07791_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1017 ();
 sky130_fd_sc_hd__mux4_1 _19692_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net658),
    .S1(net661),
    .X(_07793_));
 sky130_fd_sc_hd__mux4_1 _19693_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net658),
    .S1(net661),
    .X(_07794_));
 sky130_fd_sc_hd__mux4_1 _19694_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net658),
    .S1(net661),
    .X(_07795_));
 sky130_fd_sc_hd__mux4_1 _19695_ (.A0(_07791_),
    .A1(_07793_),
    .A2(_07794_),
    .A3(_07795_),
    .S0(net652),
    .S1(net650),
    .X(_07796_));
 sky130_fd_sc_hd__mux2i_4 _19696_ (.A0(_07790_),
    .A1(_07796_),
    .S(net649),
    .Y(_11765_));
 sky130_fd_sc_hd__mux4_1 _19697_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net656),
    .S1(net660),
    .X(_07797_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1016 ();
 sky130_fd_sc_hd__mux4_1 _19699_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net656),
    .S1(net660),
    .X(_07799_));
 sky130_fd_sc_hd__mux4_1 _19700_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net656),
    .S1(net660),
    .X(_07800_));
 sky130_fd_sc_hd__mux4_1 _19701_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net656),
    .S1(net660),
    .X(_07801_));
 sky130_fd_sc_hd__mux4_4 _19702_ (.A0(_07797_),
    .A1(_07799_),
    .A2(_07800_),
    .A3(_07801_),
    .S0(net652),
    .S1(net650),
    .X(_07802_));
 sky130_fd_sc_hd__mux4_1 _19703_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net657),
    .S1(net663),
    .X(_07803_));
 sky130_fd_sc_hd__mux4_1 _19704_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net657),
    .S1(net663),
    .X(_07804_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1015 ();
 sky130_fd_sc_hd__mux4_1 _19706_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net657),
    .S1(net663),
    .X(_07806_));
 sky130_fd_sc_hd__mux4_1 _19707_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net657),
    .S1(net663),
    .X(_07807_));
 sky130_fd_sc_hd__mux4_1 _19708_ (.A0(_07803_),
    .A1(_07804_),
    .A2(_07806_),
    .A3(_07807_),
    .S0(net652),
    .S1(net650),
    .X(_07808_));
 sky130_fd_sc_hd__mux2i_4 _19709_ (.A0(_07802_),
    .A1(_07808_),
    .S(net649),
    .Y(_11776_));
 sky130_fd_sc_hd__mux4_1 _19710_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net657),
    .S1(net660),
    .X(_07809_));
 sky130_fd_sc_hd__mux4_1 _19711_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net657),
    .S1(net660),
    .X(_07810_));
 sky130_fd_sc_hd__mux4_1 _19712_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net657),
    .S1(net660),
    .X(_07811_));
 sky130_fd_sc_hd__mux4_1 _19713_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net657),
    .S1(net660),
    .X(_07812_));
 sky130_fd_sc_hd__mux4_2 _19714_ (.A0(_07809_),
    .A1(_07810_),
    .A2(_07811_),
    .A3(_07812_),
    .S0(net652),
    .S1(net650),
    .X(_07813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1014 ();
 sky130_fd_sc_hd__mux4_1 _19716_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net657),
    .S1(net663),
    .X(_07815_));
 sky130_fd_sc_hd__mux4_1 _19717_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net657),
    .S1(net663),
    .X(_07816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1013 ();
 sky130_fd_sc_hd__mux4_1 _19719_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net657),
    .S1(net663),
    .X(_07818_));
 sky130_fd_sc_hd__mux4_1 _19720_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net657),
    .S1(net663),
    .X(_07819_));
 sky130_fd_sc_hd__mux4_1 _19721_ (.A0(_07815_),
    .A1(_07816_),
    .A2(_07818_),
    .A3(_07819_),
    .S0(net652),
    .S1(net650),
    .X(_07820_));
 sky130_fd_sc_hd__mux2i_4 _19722_ (.A0(_07813_),
    .A1(_07820_),
    .S(net649),
    .Y(_11784_));
 sky130_fd_sc_hd__mux4_1 _19723_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net659),
    .S1(net664),
    .X(_07821_));
 sky130_fd_sc_hd__mux4_1 _19724_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net659),
    .S1(net664),
    .X(_07822_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1012 ();
 sky130_fd_sc_hd__mux4_1 _19726_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net659),
    .S1(net664),
    .X(_07824_));
 sky130_fd_sc_hd__mux4_1 _19727_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net659),
    .S1(net664),
    .X(_07825_));
 sky130_fd_sc_hd__mux4_4 _19728_ (.A0(_07821_),
    .A1(_07822_),
    .A2(_07824_),
    .A3(_07825_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1011 ();
 sky130_fd_sc_hd__mux4_1 _19730_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07828_));
 sky130_fd_sc_hd__mux4_1 _19731_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07829_));
 sky130_fd_sc_hd__mux4_1 _19732_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07830_));
 sky130_fd_sc_hd__mux4_1 _19733_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07831_));
 sky130_fd_sc_hd__mux4_1 _19734_ (.A0(_07828_),
    .A1(_07829_),
    .A2(_07830_),
    .A3(_07831_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07832_));
 sky130_fd_sc_hd__mux2i_4 _19735_ (.A0(_07826_),
    .A1(_07832_),
    .S(\count16_1[5] ),
    .Y(_11792_));
 sky130_fd_sc_hd__mux4_1 _19736_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net659),
    .S1(net664),
    .X(_07833_));
 sky130_fd_sc_hd__mux4_1 _19737_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net659),
    .S1(net664),
    .X(_07834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1010 ();
 sky130_fd_sc_hd__mux4_1 _19739_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net659),
    .S1(net664),
    .X(_07836_));
 sky130_fd_sc_hd__mux4_1 _19740_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net659),
    .S1(net664),
    .X(_07837_));
 sky130_fd_sc_hd__mux4_4 _19741_ (.A0(_07833_),
    .A1(_07834_),
    .A2(_07836_),
    .A3(_07837_),
    .S0(\count16_1[3] ),
    .S1(net650),
    .X(_07838_));
 sky130_fd_sc_hd__mux4_1 _19742_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07839_));
 sky130_fd_sc_hd__mux4_1 _19743_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07840_));
 sky130_fd_sc_hd__mux4_1 _19744_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1009 ();
 sky130_fd_sc_hd__mux4_1 _19746_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1008 ();
 sky130_fd_sc_hd__mux4_1 _19748_ (.A0(_07839_),
    .A1(_07840_),
    .A2(_07841_),
    .A3(_07843_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07845_));
 sky130_fd_sc_hd__mux2i_4 _19749_ (.A0(_07838_),
    .A1(_07845_),
    .S(\count16_1[5] ),
    .Y(_11800_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1007 ();
 sky130_fd_sc_hd__mux4_1 _19751_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net658),
    .S1(net660),
    .X(_07847_));
 sky130_fd_sc_hd__mux4_1 _19752_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net658),
    .S1(net660),
    .X(_07848_));
 sky130_fd_sc_hd__mux4_1 _19753_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net658),
    .S1(net660),
    .X(_07849_));
 sky130_fd_sc_hd__mux4_1 _19754_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net658),
    .S1(net660),
    .X(_07850_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1006 ();
 sky130_fd_sc_hd__mux4_2 _19756_ (.A0(_07847_),
    .A1(_07848_),
    .A2(_07849_),
    .A3(_07850_),
    .S0(net652),
    .S1(net650),
    .X(_07852_));
 sky130_fd_sc_hd__mux4_1 _19757_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net658),
    .S1(net661),
    .X(_07853_));
 sky130_fd_sc_hd__mux4_1 _19758_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net654),
    .S1(net661),
    .X(_07854_));
 sky130_fd_sc_hd__mux4_1 _19759_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net658),
    .S1(net661),
    .X(_07855_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1005 ();
 sky130_fd_sc_hd__mux4_1 _19761_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net654),
    .S1(net661),
    .X(_07857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1004 ();
 sky130_fd_sc_hd__mux4_1 _19763_ (.A0(_07853_),
    .A1(_07854_),
    .A2(_07855_),
    .A3(_07857_),
    .S0(net653),
    .S1(net651),
    .X(_07859_));
 sky130_fd_sc_hd__mux2i_4 _19764_ (.A0(_07852_),
    .A1(_07859_),
    .S(net648),
    .Y(_11808_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1003 ();
 sky130_fd_sc_hd__mux4_1 _19766_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07861_));
 sky130_fd_sc_hd__mux4_1 _19767_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07862_));
 sky130_fd_sc_hd__mux4_1 _19768_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1002 ();
 sky130_fd_sc_hd__mux4_1 _19770_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1001 ();
 sky130_fd_sc_hd__mux4_4 _19772_ (.A0(_07861_),
    .A1(_07862_),
    .A2(_07863_),
    .A3(_07865_),
    .S0(net653),
    .S1(net651),
    .X(_07867_));
 sky130_fd_sc_hd__mux4_1 _19773_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07868_));
 sky130_fd_sc_hd__mux4_1 _19774_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07869_));
 sky130_fd_sc_hd__mux4_1 _19775_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07870_));
 sky130_fd_sc_hd__mux4_1 _19776_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net654),
    .S1(net661),
    .X(_07871_));
 sky130_fd_sc_hd__mux4_1 _19777_ (.A0(_07868_),
    .A1(_07869_),
    .A2(_07870_),
    .A3(_07871_),
    .S0(net653),
    .S1(net651),
    .X(_07872_));
 sky130_fd_sc_hd__mux2i_4 _19778_ (.A0(_07867_),
    .A1(_07872_),
    .S(net648),
    .Y(_11816_));
 sky130_fd_sc_hd__mux4_1 _19779_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07873_));
 sky130_fd_sc_hd__mux4_1 _19780_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07874_));
 sky130_fd_sc_hd__mux4_1 _19781_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1000 ();
 sky130_fd_sc_hd__mux4_1 _19783_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07877_));
 sky130_fd_sc_hd__mux4_4 _19784_ (.A0(_07873_),
    .A1(_07874_),
    .A2(_07875_),
    .A3(_07877_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07878_));
 sky130_fd_sc_hd__mux4_1 _19785_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07879_));
 sky130_fd_sc_hd__mux4_1 _19786_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07880_));
 sky130_fd_sc_hd__mux4_1 _19787_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07881_));
 sky130_fd_sc_hd__mux4_1 _19788_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07882_));
 sky130_fd_sc_hd__mux4_1 _19789_ (.A0(_07879_),
    .A1(_07880_),
    .A2(_07881_),
    .A3(_07882_),
    .S0(net653),
    .S1(\count16_1[4] ),
    .X(_07883_));
 sky130_fd_sc_hd__mux2i_4 _19790_ (.A0(_07878_),
    .A1(_07883_),
    .S(net648),
    .Y(_11824_));
 sky130_fd_sc_hd__mux4_1 _19791_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net654),
    .S1(net661),
    .X(_07884_));
 sky130_fd_sc_hd__mux4_1 _19792_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net654),
    .S1(net661),
    .X(_07885_));
 sky130_fd_sc_hd__mux4_1 _19793_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net655),
    .S1(net662),
    .X(_07886_));
 sky130_fd_sc_hd__mux4_1 _19794_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net655),
    .S1(net662),
    .X(_07887_));
 sky130_fd_sc_hd__mux4_4 _19795_ (.A0(_07884_),
    .A1(_07885_),
    .A2(_07886_),
    .A3(_07887_),
    .S0(net653),
    .S1(net651),
    .X(_07888_));
 sky130_fd_sc_hd__mux4_1 _19796_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net658),
    .S1(net662),
    .X(_07889_));
 sky130_fd_sc_hd__mux4_1 _19797_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net658),
    .S1(net662),
    .X(_07890_));
 sky130_fd_sc_hd__mux4_1 _19798_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net658),
    .S1(net662),
    .X(_07891_));
 sky130_fd_sc_hd__mux4_1 _19799_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net658),
    .S1(net662),
    .X(_07892_));
 sky130_fd_sc_hd__mux4_1 _19800_ (.A0(_07889_),
    .A1(_07890_),
    .A2(_07891_),
    .A3(_07892_),
    .S0(net653),
    .S1(net651),
    .X(_07893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_999 ();
 sky130_fd_sc_hd__mux2i_4 _19802_ (.A0(_07888_),
    .A1(_07893_),
    .S(net648),
    .Y(_11832_));
 sky130_fd_sc_hd__mux4_1 _19803_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net656),
    .S1(net660),
    .X(_07895_));
 sky130_fd_sc_hd__mux4_1 _19804_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net656),
    .S1(net660),
    .X(_07896_));
 sky130_fd_sc_hd__mux4_1 _19805_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net656),
    .S1(net660),
    .X(_07897_));
 sky130_fd_sc_hd__mux4_1 _19806_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net656),
    .S1(net660),
    .X(_07898_));
 sky130_fd_sc_hd__mux4_2 _19807_ (.A0(_07895_),
    .A1(_07896_),
    .A2(_07897_),
    .A3(_07898_),
    .S0(net652),
    .S1(net650),
    .X(_07899_));
 sky130_fd_sc_hd__mux4_1 _19808_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net657),
    .S1(net663),
    .X(_07900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_998 ();
 sky130_fd_sc_hd__mux4_1 _19810_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net657),
    .S1(net663),
    .X(_07902_));
 sky130_fd_sc_hd__mux4_1 _19811_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net657),
    .S1(net663),
    .X(_07903_));
 sky130_fd_sc_hd__mux4_1 _19812_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net657),
    .S1(net663),
    .X(_07904_));
 sky130_fd_sc_hd__mux4_1 _19813_ (.A0(_07900_),
    .A1(_07902_),
    .A2(_07903_),
    .A3(_07904_),
    .S0(net652),
    .S1(net650),
    .X(_07905_));
 sky130_fd_sc_hd__mux2i_4 _19814_ (.A0(_07899_),
    .A1(_07905_),
    .S(net649),
    .Y(_11840_));
 sky130_fd_sc_hd__mux4_1 _19815_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07906_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_997 ();
 sky130_fd_sc_hd__mux4_1 _19817_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07908_));
 sky130_fd_sc_hd__mux4_1 _19818_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07909_));
 sky130_fd_sc_hd__mux4_1 _19819_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07910_));
 sky130_fd_sc_hd__mux4_4 _19820_ (.A0(_07906_),
    .A1(_07908_),
    .A2(_07909_),
    .A3(_07910_),
    .S0(\count16_1[3] ),
    .S1(net650),
    .X(_07911_));
 sky130_fd_sc_hd__mux4_1 _19821_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net657),
    .S1(net663),
    .X(_07912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_996 ();
 sky130_fd_sc_hd__mux4_1 _19823_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07914_));
 sky130_fd_sc_hd__mux4_1 _19824_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07915_));
 sky130_fd_sc_hd__mux4_1 _19825_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07916_));
 sky130_fd_sc_hd__mux4_1 _19826_ (.A0(_07912_),
    .A1(_07914_),
    .A2(_07915_),
    .A3(_07916_),
    .S0(net652),
    .S1(net650),
    .X(_07917_));
 sky130_fd_sc_hd__mux2i_4 _19827_ (.A0(_07911_),
    .A1(_07917_),
    .S(net649),
    .Y(_11848_));
 sky130_fd_sc_hd__mux4_1 _19828_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07918_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_995 ();
 sky130_fd_sc_hd__mux4_1 _19830_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07920_));
 sky130_fd_sc_hd__mux4_1 _19831_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07921_));
 sky130_fd_sc_hd__mux4_1 _19832_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07922_));
 sky130_fd_sc_hd__mux4_2 _19833_ (.A0(_07918_),
    .A1(_07920_),
    .A2(_07921_),
    .A3(_07922_),
    .S0(net653),
    .S1(net651),
    .X(_07923_));
 sky130_fd_sc_hd__mux4_1 _19834_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07924_));
 sky130_fd_sc_hd__mux4_1 _19835_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07925_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_994 ();
 sky130_fd_sc_hd__mux4_1 _19837_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07927_));
 sky130_fd_sc_hd__mux4_1 _19838_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net654),
    .S1(net661),
    .X(_07928_));
 sky130_fd_sc_hd__mux4_1 _19839_ (.A0(_07924_),
    .A1(_07925_),
    .A2(_07927_),
    .A3(_07928_),
    .S0(net653),
    .S1(net651),
    .X(_07929_));
 sky130_fd_sc_hd__mux2i_4 _19840_ (.A0(_07923_),
    .A1(_07929_),
    .S(net648),
    .Y(_11856_));
 sky130_fd_sc_hd__mux4_1 _19841_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07930_));
 sky130_fd_sc_hd__mux4_1 _19842_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07931_));
 sky130_fd_sc_hd__mux4_1 _19843_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07932_));
 sky130_fd_sc_hd__mux4_1 _19844_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07933_));
 sky130_fd_sc_hd__mux4_2 _19845_ (.A0(_07930_),
    .A1(_07931_),
    .A2(_07932_),
    .A3(_07933_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07934_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_993 ();
 sky130_fd_sc_hd__mux4_1 _19847_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07936_));
 sky130_fd_sc_hd__mux4_1 _19848_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_992 ();
 sky130_fd_sc_hd__mux4_1 _19850_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count16_1[2] ),
    .S1(\count16_1[1] ),
    .X(_07939_));
 sky130_fd_sc_hd__mux4_1 _19851_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count16_1[2] ),
    .S1(net663),
    .X(_07940_));
 sky130_fd_sc_hd__mux4_1 _19852_ (.A0(_07936_),
    .A1(_07937_),
    .A2(_07939_),
    .A3(_07940_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07941_));
 sky130_fd_sc_hd__mux2i_4 _19853_ (.A0(_07934_),
    .A1(_07941_),
    .S(\count16_1[5] ),
    .Y(_11864_));
 sky130_fd_sc_hd__mux4_1 _19854_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net659),
    .S1(net664),
    .X(_07942_));
 sky130_fd_sc_hd__mux4_1 _19855_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net659),
    .S1(net664),
    .X(_07943_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_991 ();
 sky130_fd_sc_hd__mux4_1 _19857_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07945_));
 sky130_fd_sc_hd__mux4_1 _19858_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07946_));
 sky130_fd_sc_hd__mux4_2 _19859_ (.A0(_07942_),
    .A1(_07943_),
    .A2(_07945_),
    .A3(_07946_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07947_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_990 ();
 sky130_fd_sc_hd__mux4_1 _19861_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net659),
    .S1(net664),
    .X(_07949_));
 sky130_fd_sc_hd__mux4_1 _19862_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net659),
    .S1(net664),
    .X(_07950_));
 sky130_fd_sc_hd__mux4_1 _19863_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net659),
    .S1(net664),
    .X(_07951_));
 sky130_fd_sc_hd__mux4_1 _19864_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net659),
    .S1(net664),
    .X(_07952_));
 sky130_fd_sc_hd__mux4_1 _19865_ (.A0(_07949_),
    .A1(_07950_),
    .A2(_07951_),
    .A3(_07952_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07953_));
 sky130_fd_sc_hd__mux2i_4 _19866_ (.A0(_07947_),
    .A1(_07953_),
    .S(\count16_1[5] ),
    .Y(_11872_));
 sky130_fd_sc_hd__mux4_1 _19867_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07954_));
 sky130_fd_sc_hd__mux4_1 _19868_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07955_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_989 ();
 sky130_fd_sc_hd__mux4_1 _19870_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07957_));
 sky130_fd_sc_hd__mux4_1 _19871_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07958_));
 sky130_fd_sc_hd__mux4_4 _19872_ (.A0(_07954_),
    .A1(_07955_),
    .A2(_07957_),
    .A3(_07958_),
    .S0(net652),
    .S1(net650),
    .X(_07959_));
 sky130_fd_sc_hd__mux4_1 _19873_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07960_));
 sky130_fd_sc_hd__mux4_1 _19874_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07961_));
 sky130_fd_sc_hd__mux4_1 _19875_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07962_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_988 ();
 sky130_fd_sc_hd__mux4_1 _19877_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net657),
    .S1(net663),
    .X(_07964_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_987 ();
 sky130_fd_sc_hd__mux4_1 _19879_ (.A0(_07960_),
    .A1(_07961_),
    .A2(_07962_),
    .A3(_07964_),
    .S0(net652),
    .S1(net650),
    .X(_07966_));
 sky130_fd_sc_hd__mux2i_4 _19880_ (.A0(_07959_),
    .A1(_07966_),
    .S(net649),
    .Y(_11880_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_986 ();
 sky130_fd_sc_hd__mux4_1 _19882_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net654),
    .S1(net661),
    .X(_07968_));
 sky130_fd_sc_hd__mux4_1 _19883_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net654),
    .S1(net661),
    .X(_07969_));
 sky130_fd_sc_hd__mux4_1 _19884_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net654),
    .S1(net661),
    .X(_07970_));
 sky130_fd_sc_hd__mux4_1 _19885_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net654),
    .S1(net661),
    .X(_07971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_985 ();
 sky130_fd_sc_hd__mux4_4 _19887_ (.A0(_07968_),
    .A1(_07969_),
    .A2(_07970_),
    .A3(_07971_),
    .S0(net653),
    .S1(net651),
    .X(_07973_));
 sky130_fd_sc_hd__mux4_1 _19888_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net658),
    .S1(net661),
    .X(_07974_));
 sky130_fd_sc_hd__mux4_1 _19889_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net658),
    .S1(net661),
    .X(_07975_));
 sky130_fd_sc_hd__mux4_1 _19890_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net658),
    .S1(net661),
    .X(_07976_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_984 ();
 sky130_fd_sc_hd__mux4_1 _19892_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net658),
    .S1(net661),
    .X(_07978_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_983 ();
 sky130_fd_sc_hd__mux4_1 _19894_ (.A0(_07974_),
    .A1(_07975_),
    .A2(_07976_),
    .A3(_07978_),
    .S0(net653),
    .S1(net651),
    .X(_07980_));
 sky130_fd_sc_hd__mux2i_4 _19895_ (.A0(_07973_),
    .A1(_07980_),
    .S(net649),
    .Y(_11888_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_982 ();
 sky130_fd_sc_hd__mux4_1 _19897_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07982_));
 sky130_fd_sc_hd__mux4_1 _19898_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07983_));
 sky130_fd_sc_hd__mux4_1 _19899_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_981 ();
 sky130_fd_sc_hd__mux4_1 _19901_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07986_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_980 ();
 sky130_fd_sc_hd__mux4_2 _19903_ (.A0(_07982_),
    .A1(_07983_),
    .A2(_07984_),
    .A3(_07986_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07988_));
 sky130_fd_sc_hd__mux4_1 _19904_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07989_));
 sky130_fd_sc_hd__mux4_1 _19905_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07990_));
 sky130_fd_sc_hd__mux4_1 _19906_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07991_));
 sky130_fd_sc_hd__mux4_1 _19907_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_07992_));
 sky130_fd_sc_hd__mux4_1 _19908_ (.A0(_07989_),
    .A1(_07990_),
    .A2(_07991_),
    .A3(_07992_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07993_));
 sky130_fd_sc_hd__mux2i_4 _19909_ (.A0(_07988_),
    .A1(_07993_),
    .S(\count16_1[5] ),
    .Y(_11896_));
 sky130_fd_sc_hd__mux4_1 _19910_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07994_));
 sky130_fd_sc_hd__mux4_1 _19911_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07995_));
 sky130_fd_sc_hd__mux4_1 _19912_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07996_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_979 ();
 sky130_fd_sc_hd__mux4_1 _19914_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_07998_));
 sky130_fd_sc_hd__mux4_4 _19915_ (.A0(_07994_),
    .A1(_07995_),
    .A2(_07996_),
    .A3(_07998_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07999_));
 sky130_fd_sc_hd__mux4_1 _19916_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net659),
    .S1(net664),
    .X(_08000_));
 sky130_fd_sc_hd__mux4_1 _19917_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net659),
    .S1(net664),
    .X(_08001_));
 sky130_fd_sc_hd__mux4_1 _19918_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net659),
    .S1(net664),
    .X(_08002_));
 sky130_fd_sc_hd__mux4_1 _19919_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net659),
    .S1(net664),
    .X(_08003_));
 sky130_fd_sc_hd__mux4_1 _19920_ (.A0(_08000_),
    .A1(_08001_),
    .A2(_08002_),
    .A3(_08003_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_08004_));
 sky130_fd_sc_hd__mux2i_4 _19921_ (.A0(_07999_),
    .A1(_08004_),
    .S(\count16_1[5] ),
    .Y(_11904_));
 sky130_fd_sc_hd__mux4_1 _19922_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08005_));
 sky130_fd_sc_hd__mux4_1 _19923_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08006_));
 sky130_fd_sc_hd__mux4_1 _19924_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08007_));
 sky130_fd_sc_hd__mux4_1 _19925_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08008_));
 sky130_fd_sc_hd__mux4_4 _19926_ (.A0(_08005_),
    .A1(_08006_),
    .A2(_08007_),
    .A3(_08008_),
    .S0(net653),
    .S1(net651),
    .X(_08009_));
 sky130_fd_sc_hd__mux4_1 _19927_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08010_));
 sky130_fd_sc_hd__mux4_1 _19928_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08011_));
 sky130_fd_sc_hd__mux4_1 _19929_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08012_));
 sky130_fd_sc_hd__mux4_1 _19930_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net654),
    .S1(net661),
    .X(_08013_));
 sky130_fd_sc_hd__mux4_1 _19931_ (.A0(_08010_),
    .A1(_08011_),
    .A2(_08012_),
    .A3(_08013_),
    .S0(net653),
    .S1(net651),
    .X(_08014_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_978 ();
 sky130_fd_sc_hd__mux2i_4 _19933_ (.A0(_08009_),
    .A1(_08014_),
    .S(net648),
    .Y(_11912_));
 sky130_fd_sc_hd__mux4_1 _19934_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net656),
    .S1(net660),
    .X(_08016_));
 sky130_fd_sc_hd__mux4_1 _19935_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net656),
    .S1(net660),
    .X(_08017_));
 sky130_fd_sc_hd__mux4_1 _19936_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net656),
    .S1(net660),
    .X(_08018_));
 sky130_fd_sc_hd__mux4_1 _19937_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net656),
    .S1(net660),
    .X(_08019_));
 sky130_fd_sc_hd__mux4_4 _19938_ (.A0(_08016_),
    .A1(_08017_),
    .A2(_08018_),
    .A3(_08019_),
    .S0(net652),
    .S1(net650),
    .X(_08020_));
 sky130_fd_sc_hd__mux4_1 _19939_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net657),
    .S1(net663),
    .X(_08021_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_977 ();
 sky130_fd_sc_hd__mux4_1 _19941_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net657),
    .S1(net663),
    .X(_08023_));
 sky130_fd_sc_hd__mux4_1 _19942_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net657),
    .S1(net663),
    .X(_08024_));
 sky130_fd_sc_hd__mux4_1 _19943_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net657),
    .S1(net663),
    .X(_08025_));
 sky130_fd_sc_hd__mux4_1 _19944_ (.A0(_08021_),
    .A1(_08023_),
    .A2(_08024_),
    .A3(_08025_),
    .S0(net652),
    .S1(net650),
    .X(_08026_));
 sky130_fd_sc_hd__mux2i_4 _19945_ (.A0(_08020_),
    .A1(_08026_),
    .S(net649),
    .Y(_11920_));
 sky130_fd_sc_hd__mux4_1 _19946_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net657),
    .S1(net660),
    .X(_08027_));
 sky130_fd_sc_hd__mux4_1 _19947_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net657),
    .S1(net660),
    .X(_08028_));
 sky130_fd_sc_hd__mux4_1 _19948_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net657),
    .S1(net660),
    .X(_08029_));
 sky130_fd_sc_hd__mux4_1 _19949_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net657),
    .S1(net660),
    .X(_08030_));
 sky130_fd_sc_hd__mux4_4 _19950_ (.A0(_08027_),
    .A1(_08028_),
    .A2(_08029_),
    .A3(_08030_),
    .S0(net652),
    .S1(net650),
    .X(_08031_));
 sky130_fd_sc_hd__mux4_1 _19951_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net656),
    .S1(net660),
    .X(_08032_));
 sky130_fd_sc_hd__mux4_1 _19952_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net656),
    .S1(net660),
    .X(_08033_));
 sky130_fd_sc_hd__mux4_1 _19953_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net656),
    .S1(net660),
    .X(_08034_));
 sky130_fd_sc_hd__mux4_1 _19954_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net656),
    .S1(net660),
    .X(_08035_));
 sky130_fd_sc_hd__mux4_1 _19955_ (.A0(_08032_),
    .A1(_08033_),
    .A2(_08034_),
    .A3(_08035_),
    .S0(net652),
    .S1(net650),
    .X(_08036_));
 sky130_fd_sc_hd__mux2i_4 _19956_ (.A0(_08031_),
    .A1(_08036_),
    .S(net649),
    .Y(_11928_));
 sky130_fd_sc_hd__mux4_1 _19957_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08037_));
 sky130_fd_sc_hd__mux4_1 _19958_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08038_));
 sky130_fd_sc_hd__mux4_1 _19959_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08039_));
 sky130_fd_sc_hd__mux4_1 _19960_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08040_));
 sky130_fd_sc_hd__mux4_4 _19961_ (.A0(_08037_),
    .A1(_08038_),
    .A2(_08039_),
    .A3(_08040_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_08041_));
 sky130_fd_sc_hd__mux4_1 _19962_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net658),
    .S1(net662),
    .X(_08042_));
 sky130_fd_sc_hd__mux4_1 _19963_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net658),
    .S1(net662),
    .X(_08043_));
 sky130_fd_sc_hd__mux4_1 _19964_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net658),
    .S1(net662),
    .X(_08044_));
 sky130_fd_sc_hd__mux4_1 _19965_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net658),
    .S1(net662),
    .X(_08045_));
 sky130_fd_sc_hd__mux4_1 _19966_ (.A0(_08042_),
    .A1(_08043_),
    .A2(_08044_),
    .A3(_08045_),
    .S0(net653),
    .S1(net651),
    .X(_08046_));
 sky130_fd_sc_hd__mux2i_2 _19967_ (.A0(_08041_),
    .A1(_08046_),
    .S(net648),
    .Y(_11936_));
 sky130_fd_sc_hd__mux4_1 _19968_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08047_));
 sky130_fd_sc_hd__mux4_1 _19969_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08048_));
 sky130_fd_sc_hd__mux4_1 _19970_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08049_));
 sky130_fd_sc_hd__mux4_1 _19971_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08050_));
 sky130_fd_sc_hd__mux4_4 _19972_ (.A0(_08047_),
    .A1(_08048_),
    .A2(_08049_),
    .A3(_08050_),
    .S0(net653),
    .S1(net651),
    .X(_08051_));
 sky130_fd_sc_hd__mux4_1 _19973_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08052_));
 sky130_fd_sc_hd__mux4_1 _19974_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08053_));
 sky130_fd_sc_hd__mux4_1 _19975_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08054_));
 sky130_fd_sc_hd__mux4_1 _19976_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net655),
    .S1(net662),
    .X(_08055_));
 sky130_fd_sc_hd__mux4_1 _19977_ (.A0(_08052_),
    .A1(_08053_),
    .A2(_08054_),
    .A3(_08055_),
    .S0(net653),
    .S1(net651),
    .X(_08056_));
 sky130_fd_sc_hd__mux2i_4 _19978_ (.A0(_08051_),
    .A1(_08056_),
    .S(net648),
    .Y(_11944_));
 sky130_fd_sc_hd__mux4_1 _19979_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net656),
    .S1(net660),
    .X(_08057_));
 sky130_fd_sc_hd__mux4_1 _19980_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net656),
    .S1(net660),
    .X(_08058_));
 sky130_fd_sc_hd__mux4_1 _19981_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net656),
    .S1(net660),
    .X(_08059_));
 sky130_fd_sc_hd__mux4_1 _19982_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net656),
    .S1(net660),
    .X(_08060_));
 sky130_fd_sc_hd__mux4_4 _19983_ (.A0(_08057_),
    .A1(_08058_),
    .A2(_08059_),
    .A3(_08060_),
    .S0(net652),
    .S1(net650),
    .X(_08061_));
 sky130_fd_sc_hd__mux4_1 _19984_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net658),
    .S1(net661),
    .X(_08062_));
 sky130_fd_sc_hd__mux4_1 _19985_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net658),
    .S1(net662),
    .X(_08063_));
 sky130_fd_sc_hd__mux4_1 _19986_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net658),
    .S1(net662),
    .X(_08064_));
 sky130_fd_sc_hd__mux4_1 _19987_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net658),
    .S1(net662),
    .X(_08065_));
 sky130_fd_sc_hd__mux4_1 _19988_ (.A0(_08062_),
    .A1(_08063_),
    .A2(_08064_),
    .A3(_08065_),
    .S0(net653),
    .S1(net651),
    .X(_08066_));
 sky130_fd_sc_hd__mux2i_4 _19989_ (.A0(_08061_),
    .A1(_08066_),
    .S(net648),
    .Y(_11952_));
 sky130_fd_sc_hd__mux4_1 _19990_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net657),
    .S1(net663),
    .X(_08067_));
 sky130_fd_sc_hd__mux4_1 _19991_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net657),
    .S1(net663),
    .X(_08068_));
 sky130_fd_sc_hd__mux4_1 _19992_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net657),
    .S1(net663),
    .X(_08069_));
 sky130_fd_sc_hd__mux4_1 _19993_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net657),
    .S1(net663),
    .X(_08070_));
 sky130_fd_sc_hd__mux4_4 _19994_ (.A0(_08067_),
    .A1(_08068_),
    .A2(_08069_),
    .A3(_08070_),
    .S0(net652),
    .S1(net650),
    .X(_08071_));
 sky130_fd_sc_hd__mux4_1 _19995_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net658),
    .S1(net662),
    .X(_08072_));
 sky130_fd_sc_hd__mux4_1 _19996_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net658),
    .S1(net662),
    .X(_08073_));
 sky130_fd_sc_hd__mux4_1 _19997_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net658),
    .S1(net662),
    .X(_08074_));
 sky130_fd_sc_hd__mux4_1 _19998_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net658),
    .S1(net662),
    .X(_08075_));
 sky130_fd_sc_hd__mux4_1 _19999_ (.A0(_08072_),
    .A1(_08073_),
    .A2(_08074_),
    .A3(_08075_),
    .S0(net653),
    .S1(net651),
    .X(_08076_));
 sky130_fd_sc_hd__mux2i_4 _20000_ (.A0(_08071_),
    .A1(_08076_),
    .S(net648),
    .Y(_11960_));
 sky130_fd_sc_hd__mux4_1 _20001_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08077_));
 sky130_fd_sc_hd__mux4_1 _20002_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08078_));
 sky130_fd_sc_hd__mux4_1 _20003_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08079_));
 sky130_fd_sc_hd__mux4_1 _20004_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08080_));
 sky130_fd_sc_hd__mux4_4 _20005_ (.A0(_08077_),
    .A1(_08078_),
    .A2(_08079_),
    .A3(_08080_),
    .S0(net653),
    .S1(net651),
    .X(_08081_));
 sky130_fd_sc_hd__mux4_1 _20006_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08082_));
 sky130_fd_sc_hd__mux4_1 _20007_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08083_));
 sky130_fd_sc_hd__mux4_1 _20008_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08084_));
 sky130_fd_sc_hd__mux4_1 _20009_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net655),
    .S1(net662),
    .X(_08085_));
 sky130_fd_sc_hd__mux4_1 _20010_ (.A0(_08082_),
    .A1(_08083_),
    .A2(_08084_),
    .A3(_08085_),
    .S0(net653),
    .S1(net651),
    .X(_08086_));
 sky130_fd_sc_hd__mux2i_4 _20011_ (.A0(_08081_),
    .A1(_08086_),
    .S(net648),
    .Y(_11968_));
 sky130_fd_sc_hd__mux4_1 _20012_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08087_));
 sky130_fd_sc_hd__mux4_1 _20013_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08088_));
 sky130_fd_sc_hd__mux4_1 _20014_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08089_));
 sky130_fd_sc_hd__mux4_1 _20015_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08090_));
 sky130_fd_sc_hd__mux4_4 _20016_ (.A0(_08087_),
    .A1(_08088_),
    .A2(_08089_),
    .A3(_08090_),
    .S0(net653),
    .S1(net651),
    .X(_08091_));
 sky130_fd_sc_hd__mux4_1 _20017_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08092_));
 sky130_fd_sc_hd__mux4_1 _20018_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08093_));
 sky130_fd_sc_hd__mux4_1 _20019_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08094_));
 sky130_fd_sc_hd__mux4_1 _20020_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net655),
    .S1(net662),
    .X(_08095_));
 sky130_fd_sc_hd__mux4_1 _20021_ (.A0(_08092_),
    .A1(_08093_),
    .A2(_08094_),
    .A3(_08095_),
    .S0(net653),
    .S1(net651),
    .X(_08096_));
 sky130_fd_sc_hd__mux2i_4 _20022_ (.A0(_08091_),
    .A1(_08096_),
    .S(net648),
    .Y(_11976_));
 sky130_fd_sc_hd__mux4_1 _20023_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net656),
    .S1(net660),
    .X(_08097_));
 sky130_fd_sc_hd__mux4_1 _20024_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net656),
    .S1(net660),
    .X(_08098_));
 sky130_fd_sc_hd__mux4_1 _20025_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net656),
    .S1(net660),
    .X(_08099_));
 sky130_fd_sc_hd__mux4_1 _20026_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net656),
    .S1(net660),
    .X(_08100_));
 sky130_fd_sc_hd__mux4_4 _20027_ (.A0(_08097_),
    .A1(_08098_),
    .A2(_08099_),
    .A3(_08100_),
    .S0(net652),
    .S1(net650),
    .X(_08101_));
 sky130_fd_sc_hd__mux4_1 _20028_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net657),
    .S1(net663),
    .X(_08102_));
 sky130_fd_sc_hd__mux4_1 _20029_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net657),
    .S1(net663),
    .X(_08103_));
 sky130_fd_sc_hd__mux4_1 _20030_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net657),
    .S1(net663),
    .X(_08104_));
 sky130_fd_sc_hd__mux4_1 _20031_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net657),
    .S1(net663),
    .X(_08105_));
 sky130_fd_sc_hd__mux4_1 _20032_ (.A0(_08102_),
    .A1(_08103_),
    .A2(_08104_),
    .A3(_08105_),
    .S0(net652),
    .S1(net650),
    .X(_08106_));
 sky130_fd_sc_hd__mux2i_4 _20033_ (.A0(_08101_),
    .A1(_08106_),
    .S(net649),
    .Y(_11984_));
 sky130_fd_sc_hd__mux4_1 _20034_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08107_));
 sky130_fd_sc_hd__mux4_1 _20035_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08108_));
 sky130_fd_sc_hd__mux4_1 _20036_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08109_));
 sky130_fd_sc_hd__mux4_1 _20037_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count16_1[2] ),
    .S1(net664),
    .X(_08110_));
 sky130_fd_sc_hd__mux4_4 _20038_ (.A0(_08107_),
    .A1(_08108_),
    .A2(_08109_),
    .A3(_08110_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_08111_));
 sky130_fd_sc_hd__mux4_1 _20039_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_08112_));
 sky130_fd_sc_hd__mux4_1 _20040_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_08113_));
 sky130_fd_sc_hd__mux4_1 _20041_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_08114_));
 sky130_fd_sc_hd__mux4_1 _20042_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net659),
    .S1(\count16_1[1] ),
    .X(_08115_));
 sky130_fd_sc_hd__mux4_1 _20043_ (.A0(_08112_),
    .A1(_08113_),
    .A2(_08114_),
    .A3(_08115_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_08116_));
 sky130_fd_sc_hd__mux2i_4 _20044_ (.A0(_08111_),
    .A1(_08116_),
    .S(net649),
    .Y(_11992_));
 sky130_fd_sc_hd__inv_1 _20045_ (.A(_12258_),
    .Y(_12260_));
 sky130_fd_sc_hd__inv_1 _20046_ (.A(_12276_),
    .Y(_12279_));
 sky130_fd_sc_hd__inv_1 _20047_ (.A(_12675_),
    .Y(_12833_));
 sky130_fd_sc_hd__inv_1 _20048_ (.A(_12683_),
    .Y(_13061_));
 sky130_fd_sc_hd__inv_1 _20049_ (.A(_12830_),
    .Y(_12832_));
 sky130_fd_sc_hd__inv_1 _20050_ (.A(_12857_),
    .Y(_12858_));
 sky130_fd_sc_hd__inv_1 _20051_ (.A(_13045_),
    .Y(_13047_));
 sky130_fd_sc_hd__inv_1 _20052_ (.A(_13058_),
    .Y(\hash.CA1.p3[0] ));
 sky130_fd_sc_hd__inv_1 _20053_ (.A(_12266_),
    .Y(_12278_));
 sky130_fd_sc_hd__inv_1 _20054_ (.A(_12677_),
    .Y(_13060_));
 sky130_fd_sc_hd__inv_1 _20055_ (.A(_12826_),
    .Y(_12831_));
 sky130_fd_sc_hd__inv_1 _20056_ (.A(_12829_),
    .Y(_12841_));
 sky130_fd_sc_hd__inv_1 _20057_ (.A(_12856_),
    .Y(_12867_));
 sky130_fd_sc_hd__inv_1 _20058_ (.A(_13036_),
    .Y(_13046_));
 sky130_fd_sc_hd__clkinvlp_4 _20059_ (.A(\count_hash2[1] ),
    .Y(_00656_));
 sky130_fd_sc_hd__clkinv_2 _20060_ (.A(\count_hash1[1] ),
    .Y(_00642_));
 sky130_fd_sc_hd__xor2_1 _20061_ (.A(_11689_),
    .B(_02871_),
    .X(_08117_));
 sky130_fd_sc_hd__xnor2_1 _20062_ (.A(_11397_),
    .B(_08117_),
    .Y(_13151_));
 sky130_fd_sc_hd__inv_1 _20063_ (.A(_11761_),
    .Y(_13158_));
 sky130_fd_sc_hd__inv_1 _20064_ (.A(_11769_),
    .Y(_13162_));
 sky130_fd_sc_hd__inv_1 _20065_ (.A(_11780_),
    .Y(_13166_));
 sky130_fd_sc_hd__inv_1 _20066_ (.A(_11788_),
    .Y(_13170_));
 sky130_fd_sc_hd__inv_1 _20067_ (.A(_11796_),
    .Y(_13174_));
 sky130_fd_sc_hd__inv_1 _20068_ (.A(_11804_),
    .Y(_13178_));
 sky130_fd_sc_hd__inv_1 _20069_ (.A(_11812_),
    .Y(_13182_));
 sky130_fd_sc_hd__inv_1 _20070_ (.A(_11820_),
    .Y(_13186_));
 sky130_fd_sc_hd__inv_1 _20071_ (.A(_11828_),
    .Y(_13190_));
 sky130_fd_sc_hd__inv_1 _20072_ (.A(_11836_),
    .Y(_13194_));
 sky130_fd_sc_hd__inv_1 _20073_ (.A(_11844_),
    .Y(_13198_));
 sky130_fd_sc_hd__inv_1 _20074_ (.A(_11852_),
    .Y(_13202_));
 sky130_fd_sc_hd__inv_1 _20075_ (.A(_11860_),
    .Y(_13206_));
 sky130_fd_sc_hd__inv_1 _20076_ (.A(_11868_),
    .Y(_13210_));
 sky130_fd_sc_hd__inv_1 _20077_ (.A(_11876_),
    .Y(_13214_));
 sky130_fd_sc_hd__inv_1 _20078_ (.A(_11884_),
    .Y(_13218_));
 sky130_fd_sc_hd__inv_1 _20079_ (.A(_11892_),
    .Y(_13222_));
 sky130_fd_sc_hd__inv_1 _20080_ (.A(_11900_),
    .Y(_13226_));
 sky130_fd_sc_hd__inv_1 _20081_ (.A(_11908_),
    .Y(_13230_));
 sky130_fd_sc_hd__inv_1 _20082_ (.A(_11916_),
    .Y(_13234_));
 sky130_fd_sc_hd__inv_1 _20083_ (.A(_11924_),
    .Y(_13238_));
 sky130_fd_sc_hd__inv_1 _20084_ (.A(_11932_),
    .Y(_13242_));
 sky130_fd_sc_hd__inv_1 _20085_ (.A(_11940_),
    .Y(_13246_));
 sky130_fd_sc_hd__inv_1 _20086_ (.A(_11948_),
    .Y(_13250_));
 sky130_fd_sc_hd__inv_1 _20087_ (.A(_11956_),
    .Y(_13254_));
 sky130_fd_sc_hd__inv_1 _20088_ (.A(_11964_),
    .Y(_13258_));
 sky130_fd_sc_hd__inv_1 _20089_ (.A(_11972_),
    .Y(_13262_));
 sky130_fd_sc_hd__inv_1 _20090_ (.A(_11980_),
    .Y(_13266_));
 sky130_fd_sc_hd__inv_1 _20091_ (.A(_11988_),
    .Y(_13270_));
 sky130_fd_sc_hd__mux4_1 _20092_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net641),
    .S1(\count16_2[1] ),
    .X(_08118_));
 sky130_fd_sc_hd__mux4_1 _20093_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net641),
    .S1(\count16_2[1] ),
    .X(_08119_));
 sky130_fd_sc_hd__mux4_1 _20094_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net641),
    .S1(\count16_2[1] ),
    .X(_08120_));
 sky130_fd_sc_hd__mux4_1 _20095_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net641),
    .S1(\count16_2[1] ),
    .X(_08121_));
 sky130_fd_sc_hd__mux4_2 _20096_ (.A0(_08118_),
    .A1(_08119_),
    .A2(_08120_),
    .A3(_08121_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_08122_));
 sky130_fd_sc_hd__mux4_1 _20097_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net641),
    .S1(net642),
    .X(_08123_));
 sky130_fd_sc_hd__mux4_1 _20098_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net641),
    .S1(net642),
    .X(_08124_));
 sky130_fd_sc_hd__mux4_1 _20099_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net641),
    .S1(net642),
    .X(_08125_));
 sky130_fd_sc_hd__mux4_1 _20100_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net641),
    .S1(net642),
    .X(_08126_));
 sky130_fd_sc_hd__mux4_1 _20101_ (.A0(_08123_),
    .A1(_08124_),
    .A2(_08125_),
    .A3(_08126_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_08127_));
 sky130_fd_sc_hd__mux2_1 _20102_ (.A0(_08122_),
    .A1(_08127_),
    .S(\count16_2[5] ),
    .X(_13274_));
 sky130_fd_sc_hd__inv_1 _20103_ (.A(_12009_),
    .Y(_13281_));
 sky130_fd_sc_hd__inv_1 _20104_ (.A(_12017_),
    .Y(_13285_));
 sky130_fd_sc_hd__inv_1 _20105_ (.A(_12028_),
    .Y(_13289_));
 sky130_fd_sc_hd__inv_1 _20106_ (.A(_12036_),
    .Y(_13293_));
 sky130_fd_sc_hd__inv_1 _20107_ (.A(_12044_),
    .Y(_13297_));
 sky130_fd_sc_hd__inv_1 _20108_ (.A(_12052_),
    .Y(_13301_));
 sky130_fd_sc_hd__inv_1 _20109_ (.A(_12060_),
    .Y(_13305_));
 sky130_fd_sc_hd__inv_1 _20110_ (.A(_12068_),
    .Y(_13309_));
 sky130_fd_sc_hd__inv_1 _20111_ (.A(_12076_),
    .Y(_13313_));
 sky130_fd_sc_hd__inv_1 _20112_ (.A(_12084_),
    .Y(_13317_));
 sky130_fd_sc_hd__inv_1 _20113_ (.A(_12092_),
    .Y(_13321_));
 sky130_fd_sc_hd__inv_1 _20114_ (.A(_12100_),
    .Y(_13325_));
 sky130_fd_sc_hd__inv_1 _20115_ (.A(_12108_),
    .Y(_13329_));
 sky130_fd_sc_hd__inv_1 _20116_ (.A(_12116_),
    .Y(_13333_));
 sky130_fd_sc_hd__inv_1 _20117_ (.A(_12124_),
    .Y(_13337_));
 sky130_fd_sc_hd__inv_1 _20118_ (.A(_12132_),
    .Y(_13341_));
 sky130_fd_sc_hd__inv_1 _20119_ (.A(_12140_),
    .Y(_13345_));
 sky130_fd_sc_hd__inv_1 _20120_ (.A(_12148_),
    .Y(_13349_));
 sky130_fd_sc_hd__inv_1 _20121_ (.A(_12156_),
    .Y(_13353_));
 sky130_fd_sc_hd__inv_1 _20122_ (.A(_12164_),
    .Y(_13357_));
 sky130_fd_sc_hd__inv_1 _20123_ (.A(_12172_),
    .Y(_13361_));
 sky130_fd_sc_hd__inv_1 _20124_ (.A(_12180_),
    .Y(_13365_));
 sky130_fd_sc_hd__inv_1 _20125_ (.A(_12188_),
    .Y(_13369_));
 sky130_fd_sc_hd__inv_1 _20126_ (.A(_12196_),
    .Y(_13373_));
 sky130_fd_sc_hd__inv_1 _20127_ (.A(_12204_),
    .Y(_13377_));
 sky130_fd_sc_hd__inv_1 _20128_ (.A(_12212_),
    .Y(_13381_));
 sky130_fd_sc_hd__inv_1 _20129_ (.A(_12220_),
    .Y(_13385_));
 sky130_fd_sc_hd__inv_1 _20130_ (.A(_12228_),
    .Y(_13389_));
 sky130_fd_sc_hd__inv_1 _20131_ (.A(_12236_),
    .Y(_13393_));
 sky130_fd_sc_hd__mux2_1 _20132_ (.A0(\hash.CA2.f_dash[0] ),
    .A1(\hash.CA2.e_dash[0] ),
    .S(\hash.CA2.S1.X[0] ),
    .X(_13397_));
 sky130_fd_sc_hd__inv_1 _20133_ (.A(_12249_),
    .Y(_12264_));
 sky130_fd_sc_hd__mux2_1 _20134_ (.A0(\hash.CA2.f_dash[2] ),
    .A1(\hash.CA2.e_dash[2] ),
    .S(\hash.CA2.S1.X[2] ),
    .X(_13410_));
 sky130_fd_sc_hd__inv_1 _20135_ (.A(_12262_),
    .Y(_12273_));
 sky130_fd_sc_hd__mux2_1 _20136_ (.A0(\hash.CA2.f_dash[3] ),
    .A1(\hash.CA2.e_dash[3] ),
    .S(\hash.CA2.S1.X[3] ),
    .X(_13417_));
 sky130_fd_sc_hd__inv_1 _20137_ (.A(_12271_),
    .Y(_12287_));
 sky130_fd_sc_hd__mux2_1 _20138_ (.A0(\hash.CA2.f_dash[4] ),
    .A1(\hash.CA2.e_dash[4] ),
    .S(\hash.CA2.S1.X[4] ),
    .X(_13424_));
 sky130_fd_sc_hd__inv_1 _20139_ (.A(_12285_),
    .Y(_12296_));
 sky130_fd_sc_hd__mux2_1 _20140_ (.A0(\hash.CA2.f_dash[5] ),
    .A1(\hash.CA2.e_dash[5] ),
    .S(\hash.CA2.S1.X[5] ),
    .X(_13431_));
 sky130_fd_sc_hd__inv_1 _20141_ (.A(_12294_),
    .Y(_12305_));
 sky130_fd_sc_hd__mux2_1 _20142_ (.A0(\hash.CA2.f_dash[6] ),
    .A1(\hash.CA2.e_dash[6] ),
    .S(\hash.CA2.S1.X[6] ),
    .X(_13438_));
 sky130_fd_sc_hd__inv_1 _20143_ (.A(_12303_),
    .Y(_12314_));
 sky130_fd_sc_hd__mux2_1 _20144_ (.A0(\hash.CA2.f_dash[7] ),
    .A1(\hash.CA2.e_dash[7] ),
    .S(\hash.CA2.S1.X[7] ),
    .X(_13445_));
 sky130_fd_sc_hd__inv_1 _20145_ (.A(_12312_),
    .Y(_12323_));
 sky130_fd_sc_hd__mux2_1 _20146_ (.A0(\hash.CA2.f_dash[8] ),
    .A1(\hash.CA2.e_dash[8] ),
    .S(\hash.CA2.S1.X[8] ),
    .X(_13452_));
 sky130_fd_sc_hd__inv_1 _20147_ (.A(_12321_),
    .Y(_12332_));
 sky130_fd_sc_hd__mux2_1 _20148_ (.A0(\hash.CA2.f_dash[9] ),
    .A1(\hash.CA2.e_dash[9] ),
    .S(\hash.CA2.S1.X[9] ),
    .X(_13459_));
 sky130_fd_sc_hd__inv_1 _20149_ (.A(_12330_),
    .Y(_12341_));
 sky130_fd_sc_hd__mux2_1 _20150_ (.A0(\hash.CA2.f_dash[10] ),
    .A1(\hash.CA2.e_dash[10] ),
    .S(\hash.CA2.S1.X[10] ),
    .X(_13466_));
 sky130_fd_sc_hd__inv_1 _20151_ (.A(_12339_),
    .Y(_12350_));
 sky130_fd_sc_hd__mux2_1 _20152_ (.A0(\hash.CA2.f_dash[11] ),
    .A1(\hash.CA2.e_dash[11] ),
    .S(\hash.CA2.S1.X[11] ),
    .X(_13473_));
 sky130_fd_sc_hd__inv_1 _20153_ (.A(_12348_),
    .Y(_12359_));
 sky130_fd_sc_hd__mux2_1 _20154_ (.A0(\hash.CA2.f_dash[12] ),
    .A1(\hash.CA2.e_dash[12] ),
    .S(\hash.CA2.S1.X[12] ),
    .X(_13480_));
 sky130_fd_sc_hd__inv_1 _20155_ (.A(_12357_),
    .Y(_12368_));
 sky130_fd_sc_hd__mux2_1 _20156_ (.A0(\hash.CA2.f_dash[13] ),
    .A1(\hash.CA2.e_dash[13] ),
    .S(\hash.CA2.S1.X[13] ),
    .X(_13487_));
 sky130_fd_sc_hd__inv_1 _20157_ (.A(_12366_),
    .Y(_12377_));
 sky130_fd_sc_hd__mux2_1 _20158_ (.A0(\hash.CA2.f_dash[14] ),
    .A1(\hash.CA2.e_dash[14] ),
    .S(\hash.CA2.S1.X[14] ),
    .X(_13494_));
 sky130_fd_sc_hd__inv_1 _20159_ (.A(_12375_),
    .Y(_12386_));
 sky130_fd_sc_hd__mux2_1 _20160_ (.A0(\hash.CA2.f_dash[15] ),
    .A1(\hash.CA2.e_dash[15] ),
    .S(\hash.CA2.S1.X[15] ),
    .X(_13501_));
 sky130_fd_sc_hd__inv_1 _20161_ (.A(_12384_),
    .Y(_12395_));
 sky130_fd_sc_hd__mux2_1 _20162_ (.A0(\hash.CA2.f_dash[16] ),
    .A1(\hash.CA2.e_dash[16] ),
    .S(\hash.CA2.S1.X[16] ),
    .X(_13508_));
 sky130_fd_sc_hd__inv_1 _20163_ (.A(_12393_),
    .Y(_12404_));
 sky130_fd_sc_hd__mux2_1 _20164_ (.A0(\hash.CA2.f_dash[17] ),
    .A1(\hash.CA2.e_dash[17] ),
    .S(\hash.CA2.S1.X[17] ),
    .X(_13515_));
 sky130_fd_sc_hd__inv_1 _20165_ (.A(_12402_),
    .Y(_12413_));
 sky130_fd_sc_hd__mux2_1 _20166_ (.A0(\hash.CA2.f_dash[18] ),
    .A1(\hash.CA2.e_dash[18] ),
    .S(\hash.CA2.S1.X[18] ),
    .X(_13522_));
 sky130_fd_sc_hd__inv_1 _20167_ (.A(_12411_),
    .Y(_12422_));
 sky130_fd_sc_hd__mux2_1 _20168_ (.A0(\hash.CA2.f_dash[19] ),
    .A1(\hash.CA2.e_dash[19] ),
    .S(\hash.CA2.S1.X[19] ),
    .X(_13529_));
 sky130_fd_sc_hd__inv_1 _20169_ (.A(_12420_),
    .Y(_12431_));
 sky130_fd_sc_hd__mux2_1 _20170_ (.A0(\hash.CA2.f_dash[20] ),
    .A1(\hash.CA2.e_dash[20] ),
    .S(\hash.CA2.S1.X[20] ),
    .X(_13536_));
 sky130_fd_sc_hd__inv_1 _20171_ (.A(_12429_),
    .Y(_12440_));
 sky130_fd_sc_hd__mux2_1 _20172_ (.A0(\hash.CA2.f_dash[21] ),
    .A1(\hash.CA2.e_dash[21] ),
    .S(\hash.CA2.S1.X[21] ),
    .X(_13543_));
 sky130_fd_sc_hd__inv_1 _20173_ (.A(_12438_),
    .Y(_12449_));
 sky130_fd_sc_hd__mux2_1 _20174_ (.A0(\hash.CA2.f_dash[22] ),
    .A1(\hash.CA2.e_dash[22] ),
    .S(\hash.CA2.S1.X[22] ),
    .X(_13550_));
 sky130_fd_sc_hd__inv_1 _20175_ (.A(_12447_),
    .Y(_12458_));
 sky130_fd_sc_hd__mux2_1 _20176_ (.A0(\hash.CA2.f_dash[23] ),
    .A1(\hash.CA2.e_dash[23] ),
    .S(\hash.CA2.S1.X[23] ),
    .X(_13557_));
 sky130_fd_sc_hd__inv_1 _20177_ (.A(_12456_),
    .Y(_12467_));
 sky130_fd_sc_hd__mux2_1 _20178_ (.A0(\hash.CA2.f_dash[24] ),
    .A1(\hash.CA2.e_dash[24] ),
    .S(\hash.CA2.S1.X[24] ),
    .X(_13564_));
 sky130_fd_sc_hd__inv_1 _20179_ (.A(_12465_),
    .Y(_12476_));
 sky130_fd_sc_hd__mux2_1 _20180_ (.A0(\hash.CA2.f_dash[25] ),
    .A1(\hash.CA2.e_dash[25] ),
    .S(net1089),
    .X(_13571_));
 sky130_fd_sc_hd__inv_1 _20181_ (.A(_12474_),
    .Y(_12485_));
 sky130_fd_sc_hd__mux2_1 _20182_ (.A0(\hash.CA2.f_dash[26] ),
    .A1(\hash.CA2.e_dash[26] ),
    .S(\hash.CA2.S1.X[26] ),
    .X(_13578_));
 sky130_fd_sc_hd__inv_1 _20183_ (.A(_12483_),
    .Y(_12494_));
 sky130_fd_sc_hd__mux2_1 _20184_ (.A0(\hash.CA2.f_dash[27] ),
    .A1(\hash.CA2.e_dash[27] ),
    .S(\hash.CA2.S1.X[27] ),
    .X(_13585_));
 sky130_fd_sc_hd__inv_1 _20185_ (.A(_12492_),
    .Y(_12503_));
 sky130_fd_sc_hd__mux2_1 _20186_ (.A0(\hash.CA2.f_dash[28] ),
    .A1(\hash.CA2.e_dash[28] ),
    .S(\hash.CA2.S1.X[28] ),
    .X(_13592_));
 sky130_fd_sc_hd__inv_1 _20187_ (.A(_12501_),
    .Y(_12512_));
 sky130_fd_sc_hd__mux2_1 _20188_ (.A0(\hash.CA2.f_dash[29] ),
    .A1(\hash.CA2.e_dash[29] ),
    .S(\hash.CA2.S1.X[29] ),
    .X(_13599_));
 sky130_fd_sc_hd__inv_1 _20189_ (.A(_12510_),
    .Y(_12521_));
 sky130_fd_sc_hd__mux2_1 _20190_ (.A0(\hash.CA2.f_dash[30] ),
    .A1(\hash.CA2.e_dash[30] ),
    .S(\hash.CA2.S1.X[30] ),
    .X(_13606_));
 sky130_fd_sc_hd__inv_1 _20191_ (.A(_12519_),
    .Y(_12530_));
 sky130_fd_sc_hd__clkinvlp_4 _20192_ (.A(\count_1[1] ),
    .Y(_00651_));
 sky130_fd_sc_hd__clkinvlp_4 _20193_ (.A(\count_2[1] ),
    .Y(_00653_));
 sky130_fd_sc_hd__a21oi_1 _20194_ (.A1(\hash.CA2.a_dash[2] ),
    .A2(_12281_),
    .B1(_04592_),
    .Y(_08128_));
 sky130_fd_sc_hd__nor2_1 _20195_ (.A(\hash.CA2.a_dash[2] ),
    .B(_12281_),
    .Y(_08129_));
 sky130_fd_sc_hd__o21ai_0 _20196_ (.A1(_08128_),
    .A2(_08129_),
    .B1(net519),
    .Y(_13719_));
 sky130_fd_sc_hd__o21ai_0 _20197_ (.A1(\hash.CA1.S0.X[3] ),
    .A2(\hash.CA1.b[3] ),
    .B1(\hash.CA2.a_dash[3] ),
    .Y(_08130_));
 sky130_fd_sc_hd__o21ai_0 _20198_ (.A1(_04646_),
    .A2(_06179_),
    .B1(_08130_),
    .Y(_13723_));
 sky130_fd_sc_hd__o21bai_1 _20199_ (.A1(\hash.CA2.a_dash[4] ),
    .A2(_04654_),
    .B1_N(_06183_),
    .Y(_08131_));
 sky130_fd_sc_hd__a21oi_1 _20200_ (.A1(_04676_),
    .A2(_08131_),
    .B1(net520),
    .Y(_13727_));
 sky130_fd_sc_hd__o21ai_0 _20201_ (.A1(net520),
    .A2(_04674_),
    .B1(\hash.CA1.S0.X[5] ),
    .Y(_08132_));
 sky130_fd_sc_hd__o21ai_0 _20202_ (.A1(\hash.CA1.S0.X[5] ),
    .A2(\hash.CA1.b[5] ),
    .B1(\hash.CA2.a_dash[5] ),
    .Y(_08133_));
 sky130_fd_sc_hd__nand2_1 _20203_ (.A(_08132_),
    .B(_08133_),
    .Y(_13731_));
 sky130_fd_sc_hd__a21oi_1 _20204_ (.A1(_04701_),
    .A2(_06197_),
    .B1(net520),
    .Y(_08134_));
 sky130_fd_sc_hd__o21ai_0 _20205_ (.A1(\hash.CA1.S0.X[6] ),
    .A2(\hash.CA1.b[6] ),
    .B1(\hash.CA2.a_dash[6] ),
    .Y(_08135_));
 sky130_fd_sc_hd__nand2_1 _20206_ (.A(_08134_),
    .B(_08135_),
    .Y(_13735_));
 sky130_fd_sc_hd__a21o_1 _20207_ (.A1(net519),
    .A2(_04724_),
    .B1(\hash.CA1.S0.X[7] ),
    .X(_08136_));
 sky130_fd_sc_hd__a22o_1 _20208_ (.A1(\hash.CA1.S0.X[7] ),
    .A2(\hash.CA1.b[7] ),
    .B1(_08136_),
    .B2(\hash.CA2.a_dash[7] ),
    .X(_13739_));
 sky130_fd_sc_hd__maj3_1 _20209_ (.A(\hash.CA2.a_dash[8] ),
    .B(\hash.CA1.S0.X[8] ),
    .C(\hash.CA1.b[8] ),
    .X(_13743_));
 sky130_fd_sc_hd__maj3_1 _20210_ (.A(\hash.CA2.a_dash[9] ),
    .B(\hash.CA1.S0.X[9] ),
    .C(\hash.CA1.b[9] ),
    .X(_13747_));
 sky130_fd_sc_hd__maj3_1 _20211_ (.A(\hash.CA2.a_dash[10] ),
    .B(\hash.CA1.S0.X[10] ),
    .C(\hash.CA1.b[10] ),
    .X(_13751_));
 sky130_fd_sc_hd__a21oi_1 _20212_ (.A1(_04813_),
    .A2(_06244_),
    .B1(net520),
    .Y(_08137_));
 sky130_fd_sc_hd__a22o_1 _20213_ (.A1(\hash.CA1.S0.X[11] ),
    .A2(\hash.CA1.b[11] ),
    .B1(_08137_),
    .B2(\hash.CA2.a_dash[11] ),
    .X(_13755_));
 sky130_fd_sc_hd__maj3_1 _20214_ (.A(\hash.CA2.a_dash[12] ),
    .B(\hash.CA1.S0.X[12] ),
    .C(\hash.CA1.b[12] ),
    .X(_13759_));
 sky130_fd_sc_hd__a21oi_1 _20215_ (.A1(\hash.CA2.a_dash[13] ),
    .A2(_04842_),
    .B1(_06258_),
    .Y(_08138_));
 sky130_fd_sc_hd__o21ai_0 _20216_ (.A1(_04843_),
    .A2(_08138_),
    .B1(net519),
    .Y(_13763_));
 sky130_fd_sc_hd__a21oi_1 _20217_ (.A1(\hash.CA2.a_dash[14] ),
    .A2(_04627_),
    .B1(_06273_),
    .Y(_08139_));
 sky130_fd_sc_hd__o21ai_0 _20218_ (.A1(_04850_),
    .A2(_08139_),
    .B1(net519),
    .Y(_13767_));
 sky130_fd_sc_hd__maj3_1 _20219_ (.A(\hash.CA2.a_dash[15] ),
    .B(\hash.CA1.S0.X[15] ),
    .C(\hash.CA1.b[15] ),
    .X(_13771_));
 sky130_fd_sc_hd__maj3_1 _20220_ (.A(\hash.CA2.a_dash[16] ),
    .B(\hash.CA1.S0.X[16] ),
    .C(\hash.CA1.b[16] ),
    .X(_13775_));
 sky130_fd_sc_hd__a21oi_1 _20221_ (.A1(\hash.CA2.a_dash[17] ),
    .A2(_04699_),
    .B1(\hash.CA1.S0.X[17] ),
    .Y(_08140_));
 sky130_fd_sc_hd__o21ai_0 _20222_ (.A1(_04872_),
    .A2(_08140_),
    .B1(net519),
    .Y(_13779_));
 sky130_fd_sc_hd__a22oi_1 _20223_ (.A1(\hash.CA2.a_dash[18] ),
    .A2(_04721_),
    .B1(_06310_),
    .B2(_06311_),
    .Y(_08141_));
 sky130_fd_sc_hd__o21ai_1 _20224_ (.A1(_04880_),
    .A2(_08141_),
    .B1(net519),
    .Y(_13783_));
 sky130_fd_sc_hd__nor2_1 _20225_ (.A(net524),
    .B(_04878_),
    .Y(_08142_));
 sky130_fd_sc_hd__o21ai_0 _20226_ (.A1(\hash.CA1.S0.X[19] ),
    .A2(\hash.CA1.b[19] ),
    .B1(\hash.CA2.a_dash[19] ),
    .Y(_08143_));
 sky130_fd_sc_hd__o21ai_0 _20227_ (.A1(_06321_),
    .A2(_08142_),
    .B1(_08143_),
    .Y(_13787_));
 sky130_fd_sc_hd__maj3_1 _20228_ (.A(\hash.CA2.a_dash[20] ),
    .B(\hash.CA1.S0.X[20] ),
    .C(\hash.CA1.b[20] ),
    .X(_13791_));
 sky130_fd_sc_hd__nor2_1 _20229_ (.A(\hash.CA2.a_dash[21] ),
    .B(_04786_),
    .Y(_08144_));
 sky130_fd_sc_hd__a21oi_1 _20230_ (.A1(\hash.CA2.a_dash[21] ),
    .A2(_04786_),
    .B1(_06337_),
    .Y(_08145_));
 sky130_fd_sc_hd__o21ai_0 _20231_ (.A1(_08144_),
    .A2(_08145_),
    .B1(net519),
    .Y(_13795_));
 sky130_fd_sc_hd__a21oi_1 _20232_ (.A1(\hash.CA2.a_dash[22] ),
    .A2(net1124),
    .B1(_06349_),
    .Y(_08146_));
 sky130_fd_sc_hd__o21ai_0 _20233_ (.A1(_04910_),
    .A2(_08146_),
    .B1(net519),
    .Y(_13799_));
 sky130_fd_sc_hd__maj3_1 _20234_ (.A(\hash.CA2.a_dash[23] ),
    .B(\hash.CA1.S0.X[23] ),
    .C(_06479_),
    .X(_13803_));
 sky130_fd_sc_hd__o21ai_0 _20235_ (.A1(\hash.CA2.a_dash[24] ),
    .A2(_04652_),
    .B1(_06378_),
    .Y(_08147_));
 sky130_fd_sc_hd__a21oi_1 _20236_ (.A1(_04932_),
    .A2(_08147_),
    .B1(net521),
    .Y(_13807_));
 sky130_fd_sc_hd__maj3_1 _20237_ (.A(\hash.CA2.a_dash[25] ),
    .B(\hash.CA1.S0.X[25] ),
    .C(\hash.CA1.b[25] ),
    .X(_13811_));
 sky130_fd_sc_hd__maj3_1 _20238_ (.A(\hash.CA2.a_dash[26] ),
    .B(\hash.CA1.S0.X[26] ),
    .C(\hash.CA1.b[26] ),
    .X(_13815_));
 sky130_fd_sc_hd__nand2_1 _20239_ (.A(_04954_),
    .B(_06402_),
    .Y(_08148_));
 sky130_fd_sc_hd__o21ai_0 _20240_ (.A1(\hash.CA2.a_dash[27] ),
    .A2(_04716_),
    .B1(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand2_1 _20241_ (.A(net519),
    .B(_08149_),
    .Y(_13819_));
 sky130_fd_sc_hd__a21oi_1 _20242_ (.A1(\hash.CA2.a_dash[28] ),
    .A2(_04736_),
    .B1(_06411_),
    .Y(_08150_));
 sky130_fd_sc_hd__o21ai_0 _20243_ (.A1(_04960_),
    .A2(_08150_),
    .B1(net519),
    .Y(_13823_));
 sky130_fd_sc_hd__maj3_1 _20244_ (.A(\hash.CA2.a_dash[29] ),
    .B(\hash.CA1.S0.X[29] ),
    .C(\hash.CA1.b[29] ),
    .X(_13827_));
 sky130_fd_sc_hd__a21oi_1 _20245_ (.A1(_04977_),
    .A2(\hash.CA1.S0.X[30] ),
    .B1(_04978_),
    .Y(_08151_));
 sky130_fd_sc_hd__nor2_1 _20246_ (.A(net521),
    .B(_08151_),
    .Y(_13831_));
 sky130_fd_sc_hd__inv_1 _20247_ (.A(_12544_),
    .Y(_13835_));
 sky130_fd_sc_hd__inv_1 _20248_ (.A(_12540_),
    .Y(_12550_));
 sky130_fd_sc_hd__xor2_4 _20249_ (.A(_13846_),
    .B(_12551_),
    .X(\hash.CA1.p4[3] ));
 sky130_fd_sc_hd__inv_1 _20250_ (.A(_12555_),
    .Y(_13850_));
 sky130_fd_sc_hd__a21o_1 _20251_ (.A1(_12549_),
    .A2(_13840_),
    .B1(_13839_),
    .X(_08152_));
 sky130_fd_sc_hd__a21oi_2 _20252_ (.A1(_13846_),
    .A2(_08152_),
    .B1(_13845_),
    .Y(_08153_));
 sky130_fd_sc_hd__xnor2_4 _20253_ (.A(_13852_),
    .B(_08153_),
    .Y(\hash.CA1.p4[4] ));
 sky130_fd_sc_hd__a21o_1 _20254_ (.A1(_13846_),
    .A2(_12551_),
    .B1(_13845_),
    .X(_08154_));
 sky130_fd_sc_hd__a21oi_4 _20255_ (.A1(_13852_),
    .A2(_08154_),
    .B1(_13851_),
    .Y(_08155_));
 sky130_fd_sc_hd__xnor2_4 _20256_ (.A(_13858_),
    .B(_08155_),
    .Y(\hash.CA1.p4[5] ));
 sky130_fd_sc_hd__inv_1 _20257_ (.A(_12563_),
    .Y(_13862_));
 sky130_fd_sc_hd__inv_1 _20258_ (.A(_13852_),
    .Y(_08156_));
 sky130_fd_sc_hd__o21bai_1 _20259_ (.A1(_08156_),
    .A2(_08153_),
    .B1_N(_13851_),
    .Y(_08157_));
 sky130_fd_sc_hd__a21oi_2 _20260_ (.A1(_13858_),
    .A2(_08157_),
    .B1(_13857_),
    .Y(_08158_));
 sky130_fd_sc_hd__xnor2_4 _20261_ (.A(_13864_),
    .B(_08158_),
    .Y(\hash.CA1.p4[6] ));
 sky130_fd_sc_hd__inv_1 _20262_ (.A(_13858_),
    .Y(_08159_));
 sky130_fd_sc_hd__o21bai_1 _20263_ (.A1(_08159_),
    .A2(_08155_),
    .B1_N(_13857_),
    .Y(_08160_));
 sky130_fd_sc_hd__a21oi_2 _20264_ (.A1(_13864_),
    .A2(_08160_),
    .B1(_13863_),
    .Y(_08161_));
 sky130_fd_sc_hd__xnor2_4 _20265_ (.A(_13870_),
    .B(_08161_),
    .Y(\hash.CA1.p4[7] ));
 sky130_fd_sc_hd__inv_1 _20266_ (.A(_12571_),
    .Y(_13874_));
 sky130_fd_sc_hd__clkinvlp_4 _20267_ (.A(_13877_),
    .Y(_08162_));
 sky130_fd_sc_hd__o21a_1 _20268_ (.A1(_13864_),
    .A2(_13863_),
    .B1(_13870_),
    .X(_08163_));
 sky130_fd_sc_hd__nor2_1 _20269_ (.A(_13869_),
    .B(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__nor3_1 _20270_ (.A(_13857_),
    .B(_13863_),
    .C(_13869_),
    .Y(_08165_));
 sky130_fd_sc_hd__a21boi_1 _20271_ (.A1(_13858_),
    .A2(_08157_),
    .B1_N(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__nor2_1 _20272_ (.A(_08164_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__xnor2_4 _20273_ (.A(_08162_),
    .B(_08167_),
    .Y(\hash.CA1.p4[8] ));
 sky130_fd_sc_hd__inv_1 _20274_ (.A(_12576_),
    .Y(_13881_));
 sky130_fd_sc_hd__o21ai_1 _20275_ (.A1(_08159_),
    .A2(_08155_),
    .B1(_08165_),
    .Y(_08168_));
 sky130_fd_sc_hd__nor2_1 _20276_ (.A(_08162_),
    .B(_08164_),
    .Y(_08169_));
 sky130_fd_sc_hd__a21oi_4 _20277_ (.A1(_08168_),
    .A2(_08169_),
    .B1(_13876_),
    .Y(_08170_));
 sky130_fd_sc_hd__xnor2_2 _20278_ (.A(_13883_),
    .B(_08170_),
    .Y(\hash.CA1.p4[9] ));
 sky130_fd_sc_hd__inv_1 _20279_ (.A(_13876_),
    .Y(_08171_));
 sky130_fd_sc_hd__o31ai_2 _20280_ (.A1(_08162_),
    .A2(_08164_),
    .A3(_08166_),
    .B1(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__a21oi_4 _20281_ (.A1(_13883_),
    .A2(_08172_),
    .B1(_13882_),
    .Y(_08173_));
 sky130_fd_sc_hd__xnor2_4 _20282_ (.A(_13888_),
    .B(_08173_),
    .Y(\hash.CA1.p4[10] ));
 sky130_fd_sc_hd__inv_1 _20283_ (.A(_13883_),
    .Y(_08174_));
 sky130_fd_sc_hd__inv_1 _20284_ (.A(_13882_),
    .Y(_08175_));
 sky130_fd_sc_hd__o21ai_0 _20285_ (.A1(_08174_),
    .A2(_08170_),
    .B1(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__a21oi_1 _20286_ (.A1(_13888_),
    .A2(_08176_),
    .B1(_13887_),
    .Y(_08177_));
 sky130_fd_sc_hd__xnor2_2 _20287_ (.A(_13894_),
    .B(_08177_),
    .Y(\hash.CA1.p4[11] ));
 sky130_fd_sc_hd__inv_1 _20288_ (.A(_12587_),
    .Y(_13898_));
 sky130_fd_sc_hd__inv_1 _20289_ (.A(_13901_),
    .Y(_08178_));
 sky130_fd_sc_hd__nand2_1 _20290_ (.A(_13888_),
    .B(_13894_),
    .Y(_08179_));
 sky130_fd_sc_hd__a21oi_1 _20291_ (.A1(_13894_),
    .A2(_13887_),
    .B1(_13893_),
    .Y(_08180_));
 sky130_fd_sc_hd__o21ai_1 _20292_ (.A1(_08173_),
    .A2(_08179_),
    .B1(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__xnor2_2 _20293_ (.A(_08178_),
    .B(_08181_),
    .Y(\hash.CA1.p4[12] ));
 sky130_fd_sc_hd__inv_1 _20294_ (.A(_12592_),
    .Y(_13905_));
 sky130_fd_sc_hd__inv_1 _20295_ (.A(_13894_),
    .Y(_08182_));
 sky130_fd_sc_hd__o21bai_1 _20296_ (.A1(_08182_),
    .A2(_08177_),
    .B1_N(_13893_),
    .Y(_08183_));
 sky130_fd_sc_hd__a21oi_2 _20297_ (.A1(_13901_),
    .A2(_08183_),
    .B1(_13900_),
    .Y(_08184_));
 sky130_fd_sc_hd__xnor2_4 _20298_ (.A(_13907_),
    .B(_08184_),
    .Y(\hash.CA1.p4[13] ));
 sky130_fd_sc_hd__nand4_4 _20299_ (.A(_13888_),
    .B(_13894_),
    .C(_13901_),
    .D(_13907_),
    .Y(_08185_));
 sky130_fd_sc_hd__o21bai_1 _20300_ (.A1(_08178_),
    .A2(_08180_),
    .B1_N(_13900_),
    .Y(_08186_));
 sky130_fd_sc_hd__a21oi_4 _20301_ (.A1(_13907_),
    .A2(_08186_),
    .B1(_13906_),
    .Y(_08187_));
 sky130_fd_sc_hd__o21ai_4 _20302_ (.A1(_08173_),
    .A2(_08185_),
    .B1(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__xor2_4 _20303_ (.A(_13913_),
    .B(_08188_),
    .X(\hash.CA1.p4[14] ));
 sky130_fd_sc_hd__inv_1 _20304_ (.A(_12600_),
    .Y(_13917_));
 sky130_fd_sc_hd__or2_0 _20305_ (.A(_08175_),
    .B(_08185_),
    .X(_08189_));
 sky130_fd_sc_hd__o31ai_4 _20306_ (.A1(_08174_),
    .A2(_08170_),
    .A3(_08185_),
    .B1(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__nand2b_1 _20307_ (.A_N(_08190_),
    .B(_08187_),
    .Y(_08191_));
 sky130_fd_sc_hd__a21oi_4 _20308_ (.A1(_13913_),
    .A2(_08191_),
    .B1(_13912_),
    .Y(_08192_));
 sky130_fd_sc_hd__xnor2_4 _20309_ (.A(_13920_),
    .B(_08192_),
    .Y(\hash.CA1.p4[15] ));
 sky130_fd_sc_hd__inv_1 _20310_ (.A(_12605_),
    .Y(_13924_));
 sky130_fd_sc_hd__a21o_1 _20311_ (.A1(_13913_),
    .A2(_08188_),
    .B1(_13912_),
    .X(_08193_));
 sky130_fd_sc_hd__a21oi_2 _20312_ (.A1(_13920_),
    .A2(_08193_),
    .B1(_13919_),
    .Y(_08194_));
 sky130_fd_sc_hd__xnor2_4 _20313_ (.A(_13927_),
    .B(_08194_),
    .Y(\hash.CA1.p4[16] ));
 sky130_fd_sc_hd__inv_1 _20314_ (.A(_12610_),
    .Y(_13931_));
 sky130_fd_sc_hd__nand2_1 _20315_ (.A(_13920_),
    .B(_13927_),
    .Y(_08195_));
 sky130_fd_sc_hd__a21oi_1 _20316_ (.A1(_13927_),
    .A2(_13919_),
    .B1(_13926_),
    .Y(_08196_));
 sky130_fd_sc_hd__o21ai_2 _20317_ (.A1(_08192_),
    .A2(_08195_),
    .B1(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__xor2_4 _20318_ (.A(_13934_),
    .B(_08197_),
    .X(\hash.CA1.p4[17] ));
 sky130_fd_sc_hd__inv_1 _20319_ (.A(_12615_),
    .Y(_13938_));
 sky130_fd_sc_hd__a21o_1 _20320_ (.A1(_13920_),
    .A2(_13912_),
    .B1(_13919_),
    .X(_08198_));
 sky130_fd_sc_hd__a21o_1 _20321_ (.A1(_13927_),
    .A2(_08198_),
    .B1(_13926_),
    .X(_08199_));
 sky130_fd_sc_hd__a21oi_1 _20322_ (.A1(_13934_),
    .A2(_08199_),
    .B1(_13933_),
    .Y(_08200_));
 sky130_fd_sc_hd__and3_1 _20323_ (.A(_13920_),
    .B(_13927_),
    .C(_13934_),
    .X(_08201_));
 sky130_fd_sc_hd__nand3_1 _20324_ (.A(_13913_),
    .B(_08188_),
    .C(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_1 _20325_ (.A(_08200_),
    .B(_08202_),
    .Y(_08203_));
 sky130_fd_sc_hd__xor2_4 _20326_ (.A(_13940_),
    .B(_08203_),
    .X(\hash.CA1.p4[18] ));
 sky130_fd_sc_hd__nand3_1 _20327_ (.A(_13920_),
    .B(_13927_),
    .C(_13934_),
    .Y(_08204_));
 sky130_fd_sc_hd__nor2b_1 _20328_ (.A(_08196_),
    .B_N(_13934_),
    .Y(_08205_));
 sky130_fd_sc_hd__nor2_1 _20329_ (.A(_13933_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__o21ai_1 _20330_ (.A1(_08192_),
    .A2(_08204_),
    .B1(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__a21oi_2 _20331_ (.A1(_13940_),
    .A2(_08207_),
    .B1(_13939_),
    .Y(_08208_));
 sky130_fd_sc_hd__xnor2_4 _20332_ (.A(_13945_),
    .B(_08208_),
    .Y(\hash.CA1.p4[19] ));
 sky130_fd_sc_hd__a21bo_1 _20333_ (.A1(_08200_),
    .A2(_08202_),
    .B1_N(_13940_),
    .X(_08209_));
 sky130_fd_sc_hd__nand2b_1 _20334_ (.A_N(_13939_),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__a21oi_2 _20335_ (.A1(_13945_),
    .A2(_08210_),
    .B1(_13944_),
    .Y(_08211_));
 sky130_fd_sc_hd__xnor2_4 _20336_ (.A(_13950_),
    .B(_08211_),
    .Y(\hash.CA1.p4[20] ));
 sky130_fd_sc_hd__nand3b_1 _20337_ (.A_N(_13912_),
    .B(_08187_),
    .C(_08206_),
    .Y(_08212_));
 sky130_fd_sc_hd__nor2_1 _20338_ (.A(_13913_),
    .B(_13912_),
    .Y(_08213_));
 sky130_fd_sc_hd__o21ai_0 _20339_ (.A1(_08204_),
    .A2(_08213_),
    .B1(_08206_),
    .Y(_08214_));
 sky130_fd_sc_hd__o21ai_1 _20340_ (.A1(_08190_),
    .A2(_08212_),
    .B1(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__nand3_1 _20341_ (.A(_13940_),
    .B(_13945_),
    .C(_13950_),
    .Y(_08216_));
 sky130_fd_sc_hd__nor2_1 _20342_ (.A(_08215_),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__and3_1 _20343_ (.A(_13945_),
    .B(_13950_),
    .C(_13939_),
    .X(_08218_));
 sky130_fd_sc_hd__a2111oi_4 _20344_ (.A1(_13950_),
    .A2(_13944_),
    .B1(_13949_),
    .C1(_08217_),
    .D1(_08218_),
    .Y(_08219_));
 sky130_fd_sc_hd__xnor2_4 _20345_ (.A(_13955_),
    .B(_08219_),
    .Y(\hash.CA1.p4[21] ));
 sky130_fd_sc_hd__nor3_1 _20346_ (.A(_13939_),
    .B(_13944_),
    .C(_13949_),
    .Y(_08220_));
 sky130_fd_sc_hd__or2_0 _20347_ (.A(_13945_),
    .B(_13944_),
    .X(_08221_));
 sky130_fd_sc_hd__a21oi_1 _20348_ (.A1(_13950_),
    .A2(_08221_),
    .B1(_13949_),
    .Y(_08222_));
 sky130_fd_sc_hd__a21oi_4 _20349_ (.A1(_08209_),
    .A2(_08220_),
    .B1(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__a21oi_2 _20350_ (.A1(_13955_),
    .A2(_08223_),
    .B1(_13954_),
    .Y(_08224_));
 sky130_fd_sc_hd__xnor2_4 _20351_ (.A(_13960_),
    .B(_08224_),
    .Y(\hash.CA1.p4[22] ));
 sky130_fd_sc_hd__inv_1 _20352_ (.A(_13955_),
    .Y(_08225_));
 sky130_fd_sc_hd__o21bai_1 _20353_ (.A1(_08225_),
    .A2(_08219_),
    .B1_N(_13954_),
    .Y(_08226_));
 sky130_fd_sc_hd__a21oi_2 _20354_ (.A1(_13960_),
    .A2(_08226_),
    .B1(_13959_),
    .Y(_08227_));
 sky130_fd_sc_hd__xnor2_4 _20355_ (.A(_13966_),
    .B(_08227_),
    .Y(\hash.CA1.p4[23] ));
 sky130_fd_sc_hd__inv_1 _20356_ (.A(_12635_),
    .Y(_13970_));
 sky130_fd_sc_hd__and2_1 _20357_ (.A(_13955_),
    .B(_13960_),
    .X(_08228_));
 sky130_fd_sc_hd__a221o_1 _20358_ (.A1(_13960_),
    .A2(_13954_),
    .B1(_08223_),
    .B2(_08228_),
    .C1(_13959_),
    .X(_08229_));
 sky130_fd_sc_hd__a21oi_2 _20359_ (.A1(_13966_),
    .A2(_08229_),
    .B1(_13965_),
    .Y(_08230_));
 sky130_fd_sc_hd__xnor2_4 _20360_ (.A(_13973_),
    .B(_08230_),
    .Y(\hash.CA1.p4[24] ));
 sky130_fd_sc_hd__inv_1 _20361_ (.A(_12640_),
    .Y(_13977_));
 sky130_fd_sc_hd__inv_1 _20362_ (.A(_13966_),
    .Y(_08231_));
 sky130_fd_sc_hd__o21bai_1 _20363_ (.A1(_08231_),
    .A2(_08227_),
    .B1_N(_13965_),
    .Y(_08232_));
 sky130_fd_sc_hd__a21oi_2 _20364_ (.A1(_13973_),
    .A2(_08232_),
    .B1(_13972_),
    .Y(_08233_));
 sky130_fd_sc_hd__xnor2_4 _20365_ (.A(_13980_),
    .B(_08233_),
    .Y(\hash.CA1.p4[25] ));
 sky130_fd_sc_hd__inv_1 _20366_ (.A(_12645_),
    .Y(_13984_));
 sky130_fd_sc_hd__and3_1 _20367_ (.A(_13966_),
    .B(_13973_),
    .C(_13980_),
    .X(_08234_));
 sky130_fd_sc_hd__and3_1 _20368_ (.A(_13960_),
    .B(_13954_),
    .C(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__a21o_1 _20369_ (.A1(_13959_),
    .A2(_08234_),
    .B1(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__a31oi_4 _20370_ (.A1(_08223_),
    .A2(_08228_),
    .A3(_08234_),
    .B1(_08236_),
    .Y(_08237_));
 sky130_fd_sc_hd__a21o_1 _20371_ (.A1(_13973_),
    .A2(_13965_),
    .B1(_13972_),
    .X(_08238_));
 sky130_fd_sc_hd__a21oi_4 _20372_ (.A1(_13980_),
    .A2(_08238_),
    .B1(_13979_),
    .Y(_08239_));
 sky130_fd_sc_hd__nand2_1 _20373_ (.A(_08237_),
    .B(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__xor2_4 _20374_ (.A(_13987_),
    .B(_08240_),
    .X(\hash.CA1.p4[26] ));
 sky130_fd_sc_hd__inv_1 _20375_ (.A(_12650_),
    .Y(_13991_));
 sky130_fd_sc_hd__nand2_1 _20376_ (.A(_08228_),
    .B(_08234_),
    .Y(_08241_));
 sky130_fd_sc_hd__a22o_1 _20377_ (.A1(_13959_),
    .A2(_08234_),
    .B1(_08238_),
    .B2(_13980_),
    .X(_08242_));
 sky130_fd_sc_hd__nor3_1 _20378_ (.A(_13979_),
    .B(_08235_),
    .C(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__o21ai_0 _20379_ (.A1(_08219_),
    .A2(_08241_),
    .B1(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__a21oi_2 _20380_ (.A1(_13987_),
    .A2(_08244_),
    .B1(_13986_),
    .Y(_08245_));
 sky130_fd_sc_hd__xnor2_4 _20381_ (.A(_13994_),
    .B(_08245_),
    .Y(\hash.CA1.p4[27] ));
 sky130_fd_sc_hd__inv_1 _20382_ (.A(_12655_),
    .Y(_13998_));
 sky130_fd_sc_hd__nor2_1 _20383_ (.A(_13986_),
    .B(_13993_),
    .Y(_08246_));
 sky130_fd_sc_hd__or2_1 _20384_ (.A(_13987_),
    .B(_13986_),
    .X(_08247_));
 sky130_fd_sc_hd__a21oi_1 _20385_ (.A1(_13994_),
    .A2(_08247_),
    .B1(_13993_),
    .Y(_08248_));
 sky130_fd_sc_hd__a31oi_4 _20386_ (.A1(_08237_),
    .A2(_08239_),
    .A3(_08246_),
    .B1(_08248_),
    .Y(_08249_));
 sky130_fd_sc_hd__xor2_4 _20387_ (.A(_14001_),
    .B(_08249_),
    .X(\hash.CA1.p4[28] ));
 sky130_fd_sc_hd__inv_1 _20388_ (.A(_12660_),
    .Y(_14005_));
 sky130_fd_sc_hd__inv_1 _20389_ (.A(_13994_),
    .Y(_08250_));
 sky130_fd_sc_hd__o21bai_1 _20390_ (.A1(_08250_),
    .A2(_08245_),
    .B1_N(_13993_),
    .Y(_08251_));
 sky130_fd_sc_hd__a21oi_2 _20391_ (.A1(_14001_),
    .A2(_08251_),
    .B1(_14000_),
    .Y(_08252_));
 sky130_fd_sc_hd__xnor2_4 _20392_ (.A(_14007_),
    .B(_08252_),
    .Y(\hash.CA1.p4[29] ));
 sky130_fd_sc_hd__a21o_1 _20393_ (.A1(_14001_),
    .A2(_13993_),
    .B1(_14000_),
    .X(_08253_));
 sky130_fd_sc_hd__a21o_1 _20394_ (.A1(_14007_),
    .A2(_08253_),
    .B1(_14006_),
    .X(_08254_));
 sky130_fd_sc_hd__nor2_1 _20395_ (.A(_13986_),
    .B(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__a41oi_4 _20396_ (.A1(_13994_),
    .A2(_14001_),
    .A3(_14007_),
    .A4(_08247_),
    .B1(_08254_),
    .Y(_08256_));
 sky130_fd_sc_hd__a31oi_4 _20397_ (.A1(_08237_),
    .A2(_08239_),
    .A3(_08255_),
    .B1(_08256_),
    .Y(_08257_));
 sky130_fd_sc_hd__xor2_4 _20398_ (.A(_14012_),
    .B(_08257_),
    .X(\hash.CA1.p4[30] ));
 sky130_fd_sc_hd__mux2i_1 _20399_ (.A0(\hash.CA2.e_dash[0] ),
    .A1(\hash.CA2.S1.X[0] ),
    .S(_13613_),
    .Y(_08258_));
 sky130_fd_sc_hd__nor2_1 _20400_ (.A(\hash.reset ),
    .B(_08258_),
    .Y(_14029_));
 sky130_fd_sc_hd__mux2i_1 _20401_ (.A0(\hash.CA2.S1.X[2] ),
    .A1(\hash.CA2.e_dash[2] ),
    .S(_06687_),
    .Y(_08259_));
 sky130_fd_sc_hd__nand2_1 _20402_ (.A(_06210_),
    .B(_08259_),
    .Y(_14040_));
 sky130_fd_sc_hd__nor2_1 _20403_ (.A(\hash.CA2.e_dash[3] ),
    .B(\hash.CA1.S1.X[3] ),
    .Y(_08260_));
 sky130_fd_sc_hd__a21oi_1 _20404_ (.A1(_14019_),
    .A2(\hash.CA1.S1.X[3] ),
    .B1(_08260_),
    .Y(_14048_));
 sky130_fd_sc_hd__nand2_1 _20405_ (.A(\hash.CA1.f[4] ),
    .B(\hash.CA1.S1.X[4] ),
    .Y(_08261_));
 sky130_fd_sc_hd__o21ai_0 _20406_ (.A1(_06482_),
    .A2(\hash.CA1.S1.X[4] ),
    .B1(_08261_),
    .Y(_14057_));
 sky130_fd_sc_hd__inv_1 _20407_ (.A(_12687_),
    .Y(_14061_));
 sky130_fd_sc_hd__a21oi_1 _20408_ (.A1(_14056_),
    .A2(_07144_),
    .B1(_14055_),
    .Y(_08262_));
 sky130_fd_sc_hd__xnor2_2 _20409_ (.A(_14066_),
    .B(_08262_),
    .Y(_12695_));
 sky130_fd_sc_hd__mux2_1 _20410_ (.A0(\hash.CA1.f[5] ),
    .A1(\hash.CA2.e_dash[5] ),
    .S(_06707_),
    .X(_14067_));
 sky130_fd_sc_hd__inv_1 _20411_ (.A(_12692_),
    .Y(_14071_));
 sky130_fd_sc_hd__nand2_1 _20412_ (.A(\hash.CA2.e_dash[6] ),
    .B(_06713_),
    .Y(_08263_));
 sky130_fd_sc_hd__nand2_1 _20413_ (.A(\hash.CA1.f[6] ),
    .B(\hash.CA1.S1.X[6] ),
    .Y(_08264_));
 sky130_fd_sc_hd__nand2_1 _20414_ (.A(_08263_),
    .B(_08264_),
    .Y(_14076_));
 sky130_fd_sc_hd__nor2_1 _20415_ (.A(\hash.CA2.S1.X[7] ),
    .B(_06722_),
    .Y(_08265_));
 sky130_fd_sc_hd__a21oi_1 _20416_ (.A1(_12570_),
    .A2(_06722_),
    .B1(_08265_),
    .Y(_14084_));
 sky130_fd_sc_hd__nor2_1 _20417_ (.A(\hash.CA2.S1.X[8] ),
    .B(_06731_),
    .Y(_08266_));
 sky130_fd_sc_hd__a21oi_1 _20418_ (.A1(_12575_),
    .A2(_06731_),
    .B1(_08266_),
    .Y(_14092_));
 sky130_fd_sc_hd__nand2_1 _20419_ (.A(\hash.CA2.e_dash[9] ),
    .B(_06738_),
    .Y(_08267_));
 sky130_fd_sc_hd__nand2_1 _20420_ (.A(\hash.CA1.f[9] ),
    .B(\hash.CA1.S1.X[9] ),
    .Y(_08268_));
 sky130_fd_sc_hd__nand2_1 _20421_ (.A(_08267_),
    .B(_08268_),
    .Y(_14101_));
 sky130_fd_sc_hd__a21oi_1 _20422_ (.A1(_07341_),
    .A2(_07342_),
    .B1(_07183_),
    .Y(_12714_));
 sky130_fd_sc_hd__inv_1 _20423_ (.A(_12712_),
    .Y(_14105_));
 sky130_fd_sc_hd__mux2_1 _20424_ (.A0(_12581_),
    .A1(\hash.CA2.S1.X[10] ),
    .S(\hash.CA1.S1.X[10] ),
    .X(_14110_));
 sky130_fd_sc_hd__nor2_1 _20425_ (.A(\hash.CA2.S1.X[11] ),
    .B(_06758_),
    .Y(_08269_));
 sky130_fd_sc_hd__a21oi_1 _20426_ (.A1(_12586_),
    .A2(_06758_),
    .B1(_08269_),
    .Y(_14119_));
 sky130_fd_sc_hd__inv_1 _20427_ (.A(_12722_),
    .Y(_14123_));
 sky130_fd_sc_hd__nor2_2 _20428_ (.A(_07187_),
    .B(_07189_),
    .Y(_08270_));
 sky130_fd_sc_hd__xnor2_4 _20429_ (.A(_14128_),
    .B(_08270_),
    .Y(_12730_));
 sky130_fd_sc_hd__mux2_1 _20430_ (.A0(\hash.CA2.e_dash[12] ),
    .A1(\hash.CA1.f[12] ),
    .S(\hash.CA1.S1.X[12] ),
    .X(_14129_));
 sky130_fd_sc_hd__xnor2_1 _20431_ (.A(_07207_),
    .B(_07198_),
    .Y(_12729_));
 sky130_fd_sc_hd__inv_1 _20432_ (.A(_12727_),
    .Y(_14133_));
 sky130_fd_sc_hd__nand2_1 _20433_ (.A(_07201_),
    .B(_07202_),
    .Y(_08271_));
 sky130_fd_sc_hd__xor2_4 _20434_ (.A(_14137_),
    .B(_08271_),
    .X(_12735_));
 sky130_fd_sc_hd__nand2_1 _20435_ (.A(_12594_),
    .B(_06775_),
    .Y(_08272_));
 sky130_fd_sc_hd__o21ai_1 _20436_ (.A1(_06631_),
    .A2(_06775_),
    .B1(_08272_),
    .Y(_14138_));
 sky130_fd_sc_hd__xnor2_1 _20437_ (.A(_14141_),
    .B(_07211_),
    .Y(_12734_));
 sky130_fd_sc_hd__mux2_1 _20438_ (.A0(\hash.CA2.e_dash[14] ),
    .A1(\hash.CA1.f[14] ),
    .S(\hash.CA1.S1.X[14] ),
    .X(_14146_));
 sky130_fd_sc_hd__nor2_1 _20439_ (.A(\hash.CA2.S1.X[15] ),
    .B(_06792_),
    .Y(_08273_));
 sky130_fd_sc_hd__a21oi_1 _20440_ (.A1(_12604_),
    .A2(_06792_),
    .B1(_08273_),
    .Y(_14155_));
 sky130_fd_sc_hd__inv_1 _20441_ (.A(_12742_),
    .Y(_14159_));
 sky130_fd_sc_hd__nand3b_2 _20442_ (.A_N(_14153_),
    .B(_07217_),
    .C(_07221_),
    .Y(_08274_));
 sky130_fd_sc_hd__xor2_4 _20443_ (.A(_14164_),
    .B(_08274_),
    .X(_12750_));
 sky130_fd_sc_hd__nor3_1 _20444_ (.A(net523),
    .B(\hash.CA2.e_dash[16] ),
    .C(_06803_),
    .Y(_08275_));
 sky130_fd_sc_hd__a21oi_2 _20445_ (.A1(_06643_),
    .A2(_06804_),
    .B1(_08275_),
    .Y(_14165_));
 sky130_fd_sc_hd__xnor2_1 _20446_ (.A(_14168_),
    .B(_07344_),
    .Y(_12749_));
 sky130_fd_sc_hd__inv_1 _20447_ (.A(_12747_),
    .Y(_14169_));
 sky130_fd_sc_hd__o21ai_2 _20448_ (.A1(_07204_),
    .A2(_07228_),
    .B1(_07231_),
    .Y(_08276_));
 sky130_fd_sc_hd__xnor2_4 _20449_ (.A(_14173_),
    .B(_08276_),
    .Y(_12755_));
 sky130_fd_sc_hd__nand2_1 _20450_ (.A(\hash.CA2.e_dash[17] ),
    .B(_06816_),
    .Y(_08277_));
 sky130_fd_sc_hd__nand2_1 _20451_ (.A(\hash.CA1.f[17] ),
    .B(\hash.CA1.S1.X[17] ),
    .Y(_08278_));
 sky130_fd_sc_hd__nand2_1 _20452_ (.A(_08277_),
    .B(_08278_),
    .Y(_14174_));
 sky130_fd_sc_hd__xnor2_1 _20453_ (.A(_14177_),
    .B(_07346_),
    .Y(_12754_));
 sky130_fd_sc_hd__xor2_4 _20454_ (.A(_14181_),
    .B(_07225_),
    .X(_12760_));
 sky130_fd_sc_hd__nor2_1 _20455_ (.A(\hash.CA2.e_dash[18] ),
    .B(\hash.CA1.S1.X[18] ),
    .Y(_08279_));
 sky130_fd_sc_hd__a21oi_2 _20456_ (.A1(_06649_),
    .A2(\hash.CA1.S1.X[18] ),
    .B1(_08279_),
    .Y(_14182_));
 sky130_fd_sc_hd__xnor2_2 _20457_ (.A(_14185_),
    .B(_07349_),
    .Y(_12759_));
 sky130_fd_sc_hd__nor2_1 _20458_ (.A(_14180_),
    .B(_07234_),
    .Y(_08280_));
 sky130_fd_sc_hd__xnor2_4 _20459_ (.A(_14189_),
    .B(_08280_),
    .Y(_12765_));
 sky130_fd_sc_hd__mux2_1 _20460_ (.A0(\hash.CA1.f[19] ),
    .A1(\hash.CA2.e_dash[19] ),
    .S(_06830_),
    .X(_14190_));
 sky130_fd_sc_hd__xnor2_2 _20461_ (.A(_14193_),
    .B(_07350_),
    .Y(_12764_));
 sky130_fd_sc_hd__mux2_1 _20462_ (.A0(_12623_),
    .A1(\hash.CA2.S1.X[20] ),
    .S(\hash.CA1.S1.X[20] ),
    .X(_14198_));
 sky130_fd_sc_hd__xnor2_1 _20463_ (.A(_14201_),
    .B(_07351_),
    .Y(_12769_));
 sky130_fd_sc_hd__mux2_1 _20464_ (.A0(_12626_),
    .A1(\hash.CA2.S1.X[21] ),
    .S(\hash.CA1.S1.X[21] ),
    .X(_14206_));
 sky130_fd_sc_hd__mux2_1 _20465_ (.A0(_12629_),
    .A1(\hash.CA2.S1.X[22] ),
    .S(_06854_),
    .X(_14215_));
 sky130_fd_sc_hd__inv_1 _20466_ (.A(_12777_),
    .Y(_14219_));
 sky130_fd_sc_hd__mux2_1 _20467_ (.A0(\hash.CA2.S1.X[23] ),
    .A1(_06486_),
    .S(_06864_),
    .X(_14225_));
 sky130_fd_sc_hd__inv_1 _20468_ (.A(_12782_),
    .Y(_14229_));
 sky130_fd_sc_hd__mux2_1 _20469_ (.A0(\hash.CA2.e_dash[24] ),
    .A1(_06668_),
    .S(\hash.CA1.S1.X[24] ),
    .X(_14235_));
 sky130_fd_sc_hd__inv_1 _20470_ (.A(_12787_),
    .Y(_14239_));
 sky130_fd_sc_hd__inv_1 _20471_ (.A(\hash.CA1.S1.X[25] ),
    .Y(_08281_));
 sky130_fd_sc_hd__nor2_1 _20472_ (.A(net1030),
    .B(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__a21oi_1 _20473_ (.A1(_12644_),
    .A2(_08281_),
    .B1(_08282_),
    .Y(_14245_));
 sky130_fd_sc_hd__inv_1 _20474_ (.A(_12792_),
    .Y(_14249_));
 sky130_fd_sc_hd__o21ai_0 _20475_ (.A1(_07227_),
    .A2(_07313_),
    .B1(_07316_),
    .Y(_08283_));
 sky130_fd_sc_hd__a211oi_2 _20476_ (.A1(_14244_),
    .A2(_08283_),
    .B1(_14243_),
    .C1(_14254_),
    .Y(_08284_));
 sky130_fd_sc_hd__nor3_4 _20477_ (.A(_07314_),
    .B(_07317_),
    .C(_08284_),
    .Y(_12800_));
 sky130_fd_sc_hd__nor2_1 _20478_ (.A(\hash.CA2.S1.X[26] ),
    .B(_06886_),
    .Y(_08285_));
 sky130_fd_sc_hd__a21oi_1 _20479_ (.A1(_12649_),
    .A2(_06886_),
    .B1(_08285_),
    .Y(_14255_));
 sky130_fd_sc_hd__xnor2_1 _20480_ (.A(_14258_),
    .B(_07352_),
    .Y(_12799_));
 sky130_fd_sc_hd__inv_1 _20481_ (.A(_12797_),
    .Y(_14259_));
 sky130_fd_sc_hd__nor2_1 _20482_ (.A(net1149),
    .B(_06896_),
    .Y(_08286_));
 sky130_fd_sc_hd__a21oi_1 _20483_ (.A1(_12654_),
    .A2(_06896_),
    .B1(_08286_),
    .Y(_14264_));
 sky130_fd_sc_hd__xor2_4 _20484_ (.A(_14272_),
    .B(_07319_),
    .X(_13027_));
 sky130_fd_sc_hd__mux2_1 _20485_ (.A0(\hash.CA1.f[28] ),
    .A1(\hash.CA2.e_dash[28] ),
    .S(_06903_),
    .X(_14273_));
 sky130_fd_sc_hd__inv_1 _20486_ (.A(_12807_),
    .Y(_14277_));
 sky130_fd_sc_hd__o21bai_1 _20487_ (.A1(_07312_),
    .A2(_07307_),
    .B1_N(_14262_),
    .Y(_08287_));
 sky130_fd_sc_hd__a21oi_2 _20488_ (.A1(_14272_),
    .A2(_08287_),
    .B1(_14271_),
    .Y(_08288_));
 sky130_fd_sc_hd__xnor2_4 _20489_ (.A(_14282_),
    .B(_08288_),
    .Y(_12815_));
 sky130_fd_sc_hd__nand2_1 _20490_ (.A(\hash.CA2.S1.X[29] ),
    .B(\hash.CA1.S1.X[29] ),
    .Y(_08289_));
 sky130_fd_sc_hd__nand2_1 _20491_ (.A(_12662_),
    .B(_06910_),
    .Y(_08290_));
 sky130_fd_sc_hd__nand2_1 _20492_ (.A(_08289_),
    .B(_08290_),
    .Y(_14283_));
 sky130_fd_sc_hd__xnor2_1 _20493_ (.A(_14286_),
    .B(_07354_),
    .Y(_12814_));
 sky130_fd_sc_hd__inv_1 _20494_ (.A(_12812_),
    .Y(_14287_));
 sky130_fd_sc_hd__xor2_4 _20495_ (.A(_14291_),
    .B(_07330_),
    .X(_13041_));
 sky130_fd_sc_hd__mux2_1 _20496_ (.A0(\hash.CA1.f[30] ),
    .A1(\hash.CA2.e_dash[30] ),
    .S(_06917_),
    .X(_14292_));
 sky130_fd_sc_hd__inv_1 _20497_ (.A(_12834_),
    .Y(_14299_));
 sky130_fd_sc_hd__inv_1 _20498_ (.A(_12843_),
    .Y(_14303_));
 sky130_fd_sc_hd__inv_1 _20499_ (.A(_12848_),
    .Y(_14307_));
 sky130_fd_sc_hd__inv_1 _20500_ (.A(_12853_),
    .Y(_14311_));
 sky130_fd_sc_hd__inv_1 _20501_ (.A(_12860_),
    .Y(_14315_));
 sky130_fd_sc_hd__inv_1 _20502_ (.A(_12869_),
    .Y(_14319_));
 sky130_fd_sc_hd__inv_1 _20503_ (.A(_12877_),
    .Y(_14323_));
 sky130_fd_sc_hd__inv_1 _20504_ (.A(_12880_),
    .Y(_12889_));
 sky130_fd_sc_hd__inv_1 _20505_ (.A(_12882_),
    .Y(_14327_));
 sky130_fd_sc_hd__inv_1 _20506_ (.A(_12887_),
    .Y(_12897_));
 sky130_fd_sc_hd__inv_1 _20507_ (.A(_12895_),
    .Y(_12907_));
 sky130_fd_sc_hd__inv_1 _20508_ (.A(_12924_),
    .Y(_12933_));
 sky130_fd_sc_hd__inv_1 _20509_ (.A(_12931_),
    .Y(_12941_));
 sky130_fd_sc_hd__inv_2 _20510_ (.A(_06957_),
    .Y(_12945_));
 sky130_fd_sc_hd__inv_1 _20511_ (.A(_12966_),
    .Y(_12977_));
 sky130_fd_sc_hd__inv_1 _20512_ (.A(_12982_),
    .Y(_12993_));
 sky130_fd_sc_hd__inv_1 _20513_ (.A(_12998_),
    .Y(_13009_));
 sky130_fd_sc_hd__a21oi_1 _20514_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_13403_),
    .B1(_13090_),
    .Y(_08291_));
 sky130_fd_sc_hd__nor2_1 _20515_ (.A(\hash.CA2.a_dash[0] ),
    .B(_13403_),
    .Y(_08292_));
 sky130_fd_sc_hd__o21ai_0 _20516_ (.A1(_08291_),
    .A2(_08292_),
    .B1(net519),
    .Y(_14373_));
 sky130_fd_sc_hd__inv_1 _20517_ (.A(\count_hash2[2] ),
    .Y(_13068_));
 sky130_fd_sc_hd__inv_1 _20518_ (.A(\count_hash1[2] ),
    .Y(_13078_));
 sky130_fd_sc_hd__inv_1 _20519_ (.A(_11754_),
    .Y(_13152_));
 sky130_fd_sc_hd__inv_1 _20520_ (.A(_11762_),
    .Y(_13155_));
 sky130_fd_sc_hd__inv_1 _20521_ (.A(_11770_),
    .Y(_13159_));
 sky130_fd_sc_hd__inv_1 _20522_ (.A(_11781_),
    .Y(_13163_));
 sky130_fd_sc_hd__inv_1 _20523_ (.A(_11789_),
    .Y(_13167_));
 sky130_fd_sc_hd__inv_1 _20524_ (.A(_11797_),
    .Y(_13171_));
 sky130_fd_sc_hd__inv_1 _20525_ (.A(_11805_),
    .Y(_13175_));
 sky130_fd_sc_hd__inv_1 _20526_ (.A(_11813_),
    .Y(_13179_));
 sky130_fd_sc_hd__inv_1 _20527_ (.A(_11821_),
    .Y(_13183_));
 sky130_fd_sc_hd__inv_1 _20528_ (.A(_11829_),
    .Y(_13187_));
 sky130_fd_sc_hd__inv_1 _20529_ (.A(_11837_),
    .Y(_13191_));
 sky130_fd_sc_hd__inv_1 _20530_ (.A(_11845_),
    .Y(_13195_));
 sky130_fd_sc_hd__inv_1 _20531_ (.A(_11853_),
    .Y(_13199_));
 sky130_fd_sc_hd__inv_1 _20532_ (.A(_11861_),
    .Y(_13203_));
 sky130_fd_sc_hd__inv_1 _20533_ (.A(_11869_),
    .Y(_13207_));
 sky130_fd_sc_hd__inv_1 _20534_ (.A(_11877_),
    .Y(_13211_));
 sky130_fd_sc_hd__inv_1 _20535_ (.A(_11885_),
    .Y(_13215_));
 sky130_fd_sc_hd__inv_1 _20536_ (.A(_11893_),
    .Y(_13219_));
 sky130_fd_sc_hd__inv_1 _20537_ (.A(_11901_),
    .Y(_13223_));
 sky130_fd_sc_hd__inv_1 _20538_ (.A(_11909_),
    .Y(_13227_));
 sky130_fd_sc_hd__inv_1 _20539_ (.A(_11917_),
    .Y(_13231_));
 sky130_fd_sc_hd__inv_1 _20540_ (.A(_11925_),
    .Y(_13235_));
 sky130_fd_sc_hd__inv_1 _20541_ (.A(_11933_),
    .Y(_13239_));
 sky130_fd_sc_hd__inv_1 _20542_ (.A(_11941_),
    .Y(_13243_));
 sky130_fd_sc_hd__inv_1 _20543_ (.A(_11949_),
    .Y(_13247_));
 sky130_fd_sc_hd__inv_1 _20544_ (.A(_11957_),
    .Y(_13251_));
 sky130_fd_sc_hd__inv_1 _20545_ (.A(_11965_),
    .Y(_13255_));
 sky130_fd_sc_hd__inv_1 _20546_ (.A(_11973_),
    .Y(_13259_));
 sky130_fd_sc_hd__inv_1 _20547_ (.A(_11981_),
    .Y(_13263_));
 sky130_fd_sc_hd__inv_1 _20548_ (.A(_11989_),
    .Y(_13267_));
 sky130_fd_sc_hd__inv_1 _20549_ (.A(_11997_),
    .Y(_13271_));
 sky130_fd_sc_hd__inv_1 _20550_ (.A(_12002_),
    .Y(_13275_));
 sky130_fd_sc_hd__inv_1 _20551_ (.A(_12010_),
    .Y(_13278_));
 sky130_fd_sc_hd__inv_1 _20552_ (.A(_12018_),
    .Y(_13282_));
 sky130_fd_sc_hd__inv_1 _20553_ (.A(_12029_),
    .Y(_13286_));
 sky130_fd_sc_hd__inv_1 _20554_ (.A(_12037_),
    .Y(_13290_));
 sky130_fd_sc_hd__inv_1 _20555_ (.A(_12045_),
    .Y(_13294_));
 sky130_fd_sc_hd__inv_1 _20556_ (.A(_12053_),
    .Y(_13298_));
 sky130_fd_sc_hd__inv_1 _20557_ (.A(_12061_),
    .Y(_13302_));
 sky130_fd_sc_hd__inv_1 _20558_ (.A(_12069_),
    .Y(_13306_));
 sky130_fd_sc_hd__inv_1 _20559_ (.A(_12077_),
    .Y(_13310_));
 sky130_fd_sc_hd__inv_1 _20560_ (.A(_12085_),
    .Y(_13314_));
 sky130_fd_sc_hd__inv_1 _20561_ (.A(_12093_),
    .Y(_13318_));
 sky130_fd_sc_hd__inv_1 _20562_ (.A(_12101_),
    .Y(_13322_));
 sky130_fd_sc_hd__inv_1 _20563_ (.A(_12109_),
    .Y(_13326_));
 sky130_fd_sc_hd__inv_1 _20564_ (.A(_12117_),
    .Y(_13330_));
 sky130_fd_sc_hd__inv_1 _20565_ (.A(_12125_),
    .Y(_13334_));
 sky130_fd_sc_hd__inv_1 _20566_ (.A(_12133_),
    .Y(_13338_));
 sky130_fd_sc_hd__inv_1 _20567_ (.A(_12141_),
    .Y(_13342_));
 sky130_fd_sc_hd__inv_1 _20568_ (.A(_12149_),
    .Y(_13346_));
 sky130_fd_sc_hd__inv_1 _20569_ (.A(_12157_),
    .Y(_13350_));
 sky130_fd_sc_hd__inv_1 _20570_ (.A(_12165_),
    .Y(_13354_));
 sky130_fd_sc_hd__inv_1 _20571_ (.A(_12173_),
    .Y(_13358_));
 sky130_fd_sc_hd__inv_1 _20572_ (.A(_12181_),
    .Y(_13362_));
 sky130_fd_sc_hd__inv_1 _20573_ (.A(_12189_),
    .Y(_13366_));
 sky130_fd_sc_hd__inv_1 _20574_ (.A(_12197_),
    .Y(_13370_));
 sky130_fd_sc_hd__inv_1 _20575_ (.A(_12205_),
    .Y(_13374_));
 sky130_fd_sc_hd__inv_1 _20576_ (.A(_12213_),
    .Y(_13378_));
 sky130_fd_sc_hd__inv_1 _20577_ (.A(_12221_),
    .Y(_13382_));
 sky130_fd_sc_hd__inv_1 _20578_ (.A(_12229_),
    .Y(_13386_));
 sky130_fd_sc_hd__inv_1 _20579_ (.A(_12237_),
    .Y(_13390_));
 sky130_fd_sc_hd__inv_1 _20580_ (.A(_12245_),
    .Y(_13394_));
 sky130_fd_sc_hd__inv_1 _20581_ (.A(_12250_),
    .Y(_13401_));
 sky130_fd_sc_hd__inv_1 _20582_ (.A(_12263_),
    .Y(_12265_));
 sky130_fd_sc_hd__xnor2_2 _20583_ (.A(\hash.CA2.S1.X[27] ),
    .B(\hash.CA2.S1.X[8] ),
    .Y(_08293_));
 sky130_fd_sc_hd__xnor2_2 _20584_ (.A(\hash.CA2.S1.X[13] ),
    .B(_08293_),
    .Y(_13411_));
 sky130_fd_sc_hd__inv_1 _20585_ (.A(_12272_),
    .Y(_12274_));
 sky130_fd_sc_hd__xnor2_1 _20586_ (.A(\hash.CA2.S1.X[28] ),
    .B(\hash.CA2.S1.X[9] ),
    .Y(_08294_));
 sky130_fd_sc_hd__xnor2_2 _20587_ (.A(\hash.CA2.S1.X[14] ),
    .B(_08294_),
    .Y(_13418_));
 sky130_fd_sc_hd__inv_1 _20588_ (.A(_12286_),
    .Y(_12288_));
 sky130_fd_sc_hd__xnor2_1 _20589_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA2.S1.X[29] ),
    .Y(_08295_));
 sky130_fd_sc_hd__xnor2_2 _20590_ (.A(\hash.CA2.S1.X[15] ),
    .B(_08295_),
    .Y(_13425_));
 sky130_fd_sc_hd__inv_1 _20591_ (.A(_12295_),
    .Y(_12297_));
 sky130_fd_sc_hd__xnor2_2 _20592_ (.A(\hash.CA2.S1.X[16] ),
    .B(\hash.CA2.S1.X[30] ),
    .Y(_08296_));
 sky130_fd_sc_hd__xnor2_2 _20593_ (.A(\hash.CA2.S1.X[11] ),
    .B(_08296_),
    .Y(_13432_));
 sky130_fd_sc_hd__inv_1 _20594_ (.A(_12304_),
    .Y(_12306_));
 sky130_fd_sc_hd__xnor2_1 _20595_ (.A(\hash.CA2.S1.X[12] ),
    .B(\hash.CA2.S1.X[17] ),
    .Y(_08297_));
 sky130_fd_sc_hd__xnor2_2 _20596_ (.A(\hash.CA2.S1.X[31] ),
    .B(_08297_),
    .Y(_13439_));
 sky130_fd_sc_hd__inv_1 _20597_ (.A(_12313_),
    .Y(_12315_));
 sky130_fd_sc_hd__xnor2_1 _20598_ (.A(\hash.CA2.S1.X[18] ),
    .B(\hash.CA2.S1.X[0] ),
    .Y(_08298_));
 sky130_fd_sc_hd__xnor2_1 _20599_ (.A(\hash.CA2.S1.X[13] ),
    .B(_08298_),
    .Y(_13446_));
 sky130_fd_sc_hd__inv_1 _20600_ (.A(_12322_),
    .Y(_12324_));
 sky130_fd_sc_hd__xnor2_1 _20601_ (.A(\hash.CA2.S1.X[1] ),
    .B(\hash.CA2.S1.X[19] ),
    .Y(_08299_));
 sky130_fd_sc_hd__xnor2_1 _20602_ (.A(\hash.CA2.S1.X[14] ),
    .B(_08299_),
    .Y(_13453_));
 sky130_fd_sc_hd__inv_1 _20603_ (.A(_12331_),
    .Y(_12333_));
 sky130_fd_sc_hd__xnor2_2 _20604_ (.A(\hash.CA2.S1.X[15] ),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08300_));
 sky130_fd_sc_hd__xnor2_1 _20605_ (.A(\hash.CA2.S1.X[2] ),
    .B(_08300_),
    .Y(_13460_));
 sky130_fd_sc_hd__inv_1 _20606_ (.A(_12340_),
    .Y(_12342_));
 sky130_fd_sc_hd__xnor2_2 _20607_ (.A(\hash.CA2.S1.X[16] ),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08301_));
 sky130_fd_sc_hd__xnor2_1 _20608_ (.A(\hash.CA2.S1.X[3] ),
    .B(_08301_),
    .Y(_13467_));
 sky130_fd_sc_hd__inv_1 _20609_ (.A(_12349_),
    .Y(_12351_));
 sky130_fd_sc_hd__xnor2_1 _20610_ (.A(\hash.CA2.S1.X[17] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08302_));
 sky130_fd_sc_hd__xnor2_2 _20611_ (.A(\hash.CA2.S1.X[4] ),
    .B(_08302_),
    .Y(_13474_));
 sky130_fd_sc_hd__inv_1 _20612_ (.A(_12358_),
    .Y(_12360_));
 sky130_fd_sc_hd__xnor2_1 _20613_ (.A(\hash.CA2.S1.X[5] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08303_));
 sky130_fd_sc_hd__xnor2_1 _20614_ (.A(\hash.CA2.S1.X[18] ),
    .B(_08303_),
    .Y(_13481_));
 sky130_fd_sc_hd__inv_1 _20615_ (.A(_12367_),
    .Y(_12369_));
 sky130_fd_sc_hd__xnor2_1 _20616_ (.A(net1094),
    .B(\hash.CA2.S1.X[19] ),
    .Y(_08304_));
 sky130_fd_sc_hd__xnor2_1 _20617_ (.A(\hash.CA2.S1.X[24] ),
    .B(_08304_),
    .Y(_13488_));
 sky130_fd_sc_hd__inv_2 _20618_ (.A(_12376_),
    .Y(_12378_));
 sky130_fd_sc_hd__xnor2_1 _20619_ (.A(net1034),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08305_));
 sky130_fd_sc_hd__xnor2_1 _20620_ (.A(\hash.CA2.S1.X[7] ),
    .B(_08305_),
    .Y(_13495_));
 sky130_fd_sc_hd__inv_1 _20621_ (.A(_12385_),
    .Y(_12387_));
 sky130_fd_sc_hd__xnor2_1 _20622_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08306_));
 sky130_fd_sc_hd__xnor2_1 _20623_ (.A(\hash.CA2.S1.X[26] ),
    .B(_08306_),
    .Y(_13502_));
 sky130_fd_sc_hd__inv_1 _20624_ (.A(_12394_),
    .Y(_12396_));
 sky130_fd_sc_hd__xnor2_1 _20625_ (.A(\hash.CA2.S1.X[9] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08307_));
 sky130_fd_sc_hd__xnor2_1 _20626_ (.A(\hash.CA2.S1.X[27] ),
    .B(_08307_),
    .Y(_13509_));
 sky130_fd_sc_hd__inv_1 _20627_ (.A(_12403_),
    .Y(_12405_));
 sky130_fd_sc_hd__xnor2_1 _20628_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08308_));
 sky130_fd_sc_hd__xnor2_1 _20629_ (.A(\hash.CA2.S1.X[28] ),
    .B(_08308_),
    .Y(_13516_));
 sky130_fd_sc_hd__inv_1 _20630_ (.A(_12412_),
    .Y(_12414_));
 sky130_fd_sc_hd__xnor2_1 _20631_ (.A(\hash.CA2.S1.X[24] ),
    .B(\hash.CA2.S1.X[29] ),
    .Y(_08309_));
 sky130_fd_sc_hd__xnor2_2 _20632_ (.A(\hash.CA2.S1.X[11] ),
    .B(_08309_),
    .Y(_13523_));
 sky130_fd_sc_hd__inv_1 _20633_ (.A(_12421_),
    .Y(_12423_));
 sky130_fd_sc_hd__xnor2_1 _20634_ (.A(\hash.CA2.S1.X[12] ),
    .B(\hash.CA2.S1.X[30] ),
    .Y(_08310_));
 sky130_fd_sc_hd__xnor2_1 _20635_ (.A(net1090),
    .B(_08310_),
    .Y(_13530_));
 sky130_fd_sc_hd__inv_1 _20636_ (.A(_12430_),
    .Y(_12432_));
 sky130_fd_sc_hd__xnor2_1 _20637_ (.A(\hash.CA2.S1.X[31] ),
    .B(\hash.CA2.S1.X[26] ),
    .Y(_08311_));
 sky130_fd_sc_hd__xnor2_1 _20638_ (.A(\hash.CA2.S1.X[13] ),
    .B(_08311_),
    .Y(_13537_));
 sky130_fd_sc_hd__inv_1 _20639_ (.A(_12439_),
    .Y(_12441_));
 sky130_fd_sc_hd__xnor2_1 _20640_ (.A(\hash.CA2.S1.X[27] ),
    .B(\hash.CA2.S1.X[0] ),
    .Y(_08312_));
 sky130_fd_sc_hd__xnor2_2 _20641_ (.A(\hash.CA2.S1.X[14] ),
    .B(_08312_),
    .Y(_13544_));
 sky130_fd_sc_hd__inv_1 _20642_ (.A(_12448_),
    .Y(_12450_));
 sky130_fd_sc_hd__xnor2_2 _20643_ (.A(\hash.CA2.S1.X[1] ),
    .B(\hash.CA2.S1.X[15] ),
    .Y(_08313_));
 sky130_fd_sc_hd__xnor2_1 _20644_ (.A(\hash.CA2.S1.X[28] ),
    .B(_08313_),
    .Y(_13551_));
 sky130_fd_sc_hd__inv_1 _20645_ (.A(_12457_),
    .Y(_12459_));
 sky130_fd_sc_hd__xnor2_1 _20646_ (.A(\hash.CA2.S1.X[16] ),
    .B(\hash.CA2.S1.X[29] ),
    .Y(_08314_));
 sky130_fd_sc_hd__xnor2_2 _20647_ (.A(\hash.CA2.S1.X[2] ),
    .B(_08314_),
    .Y(_13558_));
 sky130_fd_sc_hd__inv_1 _20648_ (.A(_12466_),
    .Y(_12468_));
 sky130_fd_sc_hd__xnor2_1 _20649_ (.A(\hash.CA2.S1.X[30] ),
    .B(\hash.CA2.S1.X[17] ),
    .Y(_08315_));
 sky130_fd_sc_hd__xnor2_1 _20650_ (.A(\hash.CA2.S1.X[3] ),
    .B(_08315_),
    .Y(_13565_));
 sky130_fd_sc_hd__inv_1 _20651_ (.A(_12475_),
    .Y(_12477_));
 sky130_fd_sc_hd__xnor2_1 _20652_ (.A(\hash.CA2.S1.X[31] ),
    .B(\hash.CA2.S1.X[4] ),
    .Y(_08316_));
 sky130_fd_sc_hd__xnor2_1 _20653_ (.A(\hash.CA2.S1.X[18] ),
    .B(_08316_),
    .Y(_13572_));
 sky130_fd_sc_hd__inv_1 _20654_ (.A(_12484_),
    .Y(_12486_));
 sky130_fd_sc_hd__xnor2_2 _20655_ (.A(\hash.CA2.S1.X[5] ),
    .B(\hash.CA2.S1.X[19] ),
    .Y(_08317_));
 sky130_fd_sc_hd__xnor2_4 _20656_ (.A(\hash.CA2.S1.X[0] ),
    .B(_08317_),
    .Y(_13579_));
 sky130_fd_sc_hd__inv_1 _20657_ (.A(_12493_),
    .Y(_12495_));
 sky130_fd_sc_hd__xnor2_2 _20658_ (.A(\hash.CA2.S1.X[1] ),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08318_));
 sky130_fd_sc_hd__xnor2_4 _20659_ (.A(net1095),
    .B(_08318_),
    .Y(_13586_));
 sky130_fd_sc_hd__inv_1 _20660_ (.A(_12502_),
    .Y(_12504_));
 sky130_fd_sc_hd__xnor2_2 _20661_ (.A(\hash.CA2.S1.X[7] ),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08319_));
 sky130_fd_sc_hd__xnor2_4 _20662_ (.A(\hash.CA2.S1.X[2] ),
    .B(_08319_),
    .Y(_13593_));
 sky130_fd_sc_hd__inv_1 _20663_ (.A(_12511_),
    .Y(_12513_));
 sky130_fd_sc_hd__xnor2_1 _20664_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08320_));
 sky130_fd_sc_hd__xnor2_2 _20665_ (.A(\hash.CA2.S1.X[3] ),
    .B(_08320_),
    .Y(_13600_));
 sky130_fd_sc_hd__inv_1 _20666_ (.A(_12520_),
    .Y(_12522_));
 sky130_fd_sc_hd__xnor2_1 _20667_ (.A(\hash.CA2.S1.X[4] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08321_));
 sky130_fd_sc_hd__xnor2_2 _20668_ (.A(\hash.CA2.S1.X[9] ),
    .B(_08321_),
    .Y(_13607_));
 sky130_fd_sc_hd__inv_1 _20669_ (.A(_12529_),
    .Y(_12531_));
 sky130_fd_sc_hd__xnor2_2 _20670_ (.A(_04916_),
    .B(_13553_),
    .Y(_13554_));
 sky130_fd_sc_hd__xor2_1 _20671_ (.A(_13609_),
    .B(_04980_),
    .X(_13610_));
 sky130_fd_sc_hd__inv_1 _20672_ (.A(\count_1[2] ),
    .Y(_13695_));
 sky130_fd_sc_hd__inv_1 _20673_ (.A(\count_2[2] ),
    .Y(_13703_));
 sky130_fd_sc_hd__xnor2_2 _20674_ (.A(\hash.CA1.S0.X[4] ),
    .B(_06283_),
    .Y(_08322_));
 sky130_fd_sc_hd__xor2_4 _20675_ (.A(_08322_),
    .B(\hash.CA1.S0.X[24] ),
    .X(_13720_));
 sky130_fd_sc_hd__xnor2_2 _20676_ (.A(_06190_),
    .B(_06291_),
    .Y(_08323_));
 sky130_fd_sc_hd__xnor2_4 _20677_ (.A(\hash.CA1.S0.X[25] ),
    .B(_08323_),
    .Y(_13724_));
 sky130_fd_sc_hd__xnor2_2 _20678_ (.A(\hash.CA1.S0.X[6] ),
    .B(\hash.CA1.S0.X[17] ),
    .Y(_08324_));
 sky130_fd_sc_hd__xnor2_4 _20679_ (.A(\hash.CA1.S0.X[26] ),
    .B(_08324_),
    .Y(_13728_));
 sky130_fd_sc_hd__xor2_2 _20680_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06312_),
    .X(_08325_));
 sky130_fd_sc_hd__xnor2_4 _20681_ (.A(_06402_),
    .B(_08325_),
    .Y(_13732_));
 sky130_fd_sc_hd__xnor2_2 _20682_ (.A(\hash.CA1.S0.X[8] ),
    .B(_06321_),
    .Y(_08326_));
 sky130_fd_sc_hd__xnor2_4 _20683_ (.A(_06412_),
    .B(_08326_),
    .Y(_13736_));
 sky130_fd_sc_hd__xnor2_2 _20684_ (.A(_06227_),
    .B(\hash.CA1.S0.X[20] ),
    .Y(_08327_));
 sky130_fd_sc_hd__xnor2_4 _20685_ (.A(_06417_),
    .B(_08327_),
    .Y(_13740_));
 sky130_fd_sc_hd__xnor2_2 _20686_ (.A(\hash.CA1.S0.X[10] ),
    .B(_06338_),
    .Y(_08328_));
 sky130_fd_sc_hd__xnor2_4 _20687_ (.A(\hash.CA1.S0.X[30] ),
    .B(_08328_),
    .Y(_13744_));
 sky130_fd_sc_hd__xnor2_1 _20688_ (.A(\hash.CA1.S0.X[11] ),
    .B(_06349_),
    .Y(_08329_));
 sky130_fd_sc_hd__xnor2_1 _20689_ (.A(_06462_),
    .B(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__nor2_1 _20690_ (.A(net524),
    .B(_08330_),
    .Y(_13748_));
 sky130_fd_sc_hd__xnor2_1 _20691_ (.A(_13403_),
    .B(_06251_),
    .Y(_08331_));
 sky130_fd_sc_hd__nor2_1 _20692_ (.A(net524),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__xnor2_1 _20693_ (.A(net1128),
    .B(_08332_),
    .Y(_13752_));
 sky130_fd_sc_hd__xnor2_1 _20694_ (.A(_13409_),
    .B(_06258_),
    .Y(_08333_));
 sky130_fd_sc_hd__xnor2_1 _20695_ (.A(_06367_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__nor2_1 _20696_ (.A(net524),
    .B(_08334_),
    .Y(_13756_));
 sky130_fd_sc_hd__xor2_1 _20697_ (.A(_12281_),
    .B(_06273_),
    .X(_08335_));
 sky130_fd_sc_hd__xnor2_1 _20698_ (.A(net1157),
    .B(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__nand2_1 _20699_ (.A(net519),
    .B(_08336_),
    .Y(_13760_));
 sky130_fd_sc_hd__xnor2_1 _20700_ (.A(_06179_),
    .B(_06283_),
    .Y(_08337_));
 sky130_fd_sc_hd__xnor2_1 _20701_ (.A(\hash.CA1.S0.X[26] ),
    .B(_08337_),
    .Y(_13764_));
 sky130_fd_sc_hd__xnor2_1 _20702_ (.A(\hash.CA1.S0.X[4] ),
    .B(_06291_),
    .Y(_08338_));
 sky130_fd_sc_hd__xnor2_2 _20703_ (.A(_06402_),
    .B(_08338_),
    .Y(_13768_));
 sky130_fd_sc_hd__xnor2_1 _20704_ (.A(_06190_),
    .B(\hash.CA1.S0.X[17] ),
    .Y(_08339_));
 sky130_fd_sc_hd__xnor2_1 _20705_ (.A(_06412_),
    .B(_08339_),
    .Y(_13772_));
 sky130_fd_sc_hd__xnor2_1 _20706_ (.A(_06198_),
    .B(_06312_),
    .Y(_08340_));
 sky130_fd_sc_hd__xnor2_1 _20707_ (.A(_06417_),
    .B(_08340_),
    .Y(_13776_));
 sky130_fd_sc_hd__xnor2_1 _20708_ (.A(\hash.CA1.S0.X[7] ),
    .B(\hash.CA1.S0.X[19] ),
    .Y(_08341_));
 sky130_fd_sc_hd__xnor2_1 _20709_ (.A(\hash.CA1.S0.X[30] ),
    .B(_08341_),
    .Y(_13780_));
 sky130_fd_sc_hd__xnor2_1 _20710_ (.A(\hash.CA1.S0.X[8] ),
    .B(\hash.CA1.S0.X[20] ),
    .Y(_08342_));
 sky130_fd_sc_hd__xnor2_1 _20711_ (.A(_06462_),
    .B(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__nor2_1 _20712_ (.A(net524),
    .B(_08343_),
    .Y(_13784_));
 sky130_fd_sc_hd__xor2_1 _20713_ (.A(_13403_),
    .B(_06337_),
    .X(_08344_));
 sky130_fd_sc_hd__nor2_1 _20714_ (.A(net524),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__xnor2_1 _20715_ (.A(\hash.CA1.S0.X[9] ),
    .B(_08345_),
    .Y(_13788_));
 sky130_fd_sc_hd__xor2_1 _20716_ (.A(_13409_),
    .B(_06349_),
    .X(_08346_));
 sky130_fd_sc_hd__nor2_1 _20717_ (.A(net524),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__xnor2_1 _20718_ (.A(\hash.CA1.S0.X[10] ),
    .B(_08347_),
    .Y(_13792_));
 sky130_fd_sc_hd__nor2_1 _20719_ (.A(\hash.CA1.S0.X[2] ),
    .B(net1127),
    .Y(_08348_));
 sky130_fd_sc_hd__a21oi_1 _20720_ (.A1(_12281_),
    .A2(net1127),
    .B1(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__xor2_2 _20721_ (.A(\hash.CA1.S0.X[11] ),
    .B(_08349_),
    .X(_13796_));
 sky130_fd_sc_hd__xnor2_4 _20722_ (.A(\hash.CA1.S0.X[3] ),
    .B(\hash.CA1.S0.X[12] ),
    .Y(_08350_));
 sky130_fd_sc_hd__xnor2_1 _20723_ (.A(\hash.CA1.S0.X[24] ),
    .B(_08350_),
    .Y(_13800_));
 sky130_fd_sc_hd__xnor2_2 _20724_ (.A(\hash.CA1.S0.X[4] ),
    .B(_06259_),
    .Y(_08351_));
 sky130_fd_sc_hd__xnor2_1 _20725_ (.A(_06377_),
    .B(_08351_),
    .Y(_13804_));
 sky130_fd_sc_hd__xnor2_2 _20726_ (.A(_06190_),
    .B(_06274_),
    .Y(_08352_));
 sky130_fd_sc_hd__xnor2_1 _20727_ (.A(\hash.CA1.S0.X[26] ),
    .B(_08352_),
    .Y(_13808_));
 sky130_fd_sc_hd__xnor2_4 _20728_ (.A(\hash.CA1.S0.X[6] ),
    .B(_06283_),
    .Y(_08353_));
 sky130_fd_sc_hd__xnor2_1 _20729_ (.A(_06402_),
    .B(_08353_),
    .Y(_13812_));
 sky130_fd_sc_hd__xnor2_2 _20730_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06291_),
    .Y(_08354_));
 sky130_fd_sc_hd__xnor2_1 _20731_ (.A(_06412_),
    .B(_08354_),
    .Y(_13816_));
 sky130_fd_sc_hd__xnor2_4 _20732_ (.A(_06219_),
    .B(\hash.CA1.S0.X[17] ),
    .Y(_08355_));
 sky130_fd_sc_hd__xnor2_1 _20733_ (.A(_06417_),
    .B(_08355_),
    .Y(_13820_));
 sky130_fd_sc_hd__xnor2_2 _20734_ (.A(\hash.CA1.S0.X[9] ),
    .B(_06312_),
    .Y(_08356_));
 sky130_fd_sc_hd__xnor2_1 _20735_ (.A(\hash.CA1.S0.X[30] ),
    .B(_08356_),
    .Y(_13824_));
 sky130_fd_sc_hd__xnor2_2 _20736_ (.A(_06236_),
    .B(_06321_),
    .Y(_08357_));
 sky130_fd_sc_hd__xnor2_1 _20737_ (.A(_06462_),
    .B(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__nor2_1 _20738_ (.A(net521),
    .B(_08358_),
    .Y(_13828_));
 sky130_fd_sc_hd__nor2_1 _20739_ (.A(\hash.CA1.S0.X[0] ),
    .B(\hash.CA1.S0.X[11] ),
    .Y(_08359_));
 sky130_fd_sc_hd__a21oi_4 _20740_ (.A1(_13403_),
    .A2(\hash.CA1.S0.X[11] ),
    .B1(_08359_),
    .Y(_08360_));
 sky130_fd_sc_hd__xnor2_2 _20741_ (.A(_06332_),
    .B(_08360_),
    .Y(_13832_));
 sky130_fd_sc_hd__inv_1 _20742_ (.A(_12541_),
    .Y(_13836_));
 sky130_fd_sc_hd__inv_1 _20743_ (.A(_12556_),
    .Y(_13844_));
 sky130_fd_sc_hd__inv_1 _20744_ (.A(_12564_),
    .Y(_13856_));
 sky130_fd_sc_hd__inv_1 _20745_ (.A(_12572_),
    .Y(_13868_));
 sky130_fd_sc_hd__inv_1 _20746_ (.A(_06996_),
    .Y(_13871_));
 sky130_fd_sc_hd__inv_1 _20747_ (.A(_12577_),
    .Y(_13875_));
 sky130_fd_sc_hd__inv_1 _20748_ (.A(_12588_),
    .Y(_13892_));
 sky130_fd_sc_hd__inv_1 _20749_ (.A(_12593_),
    .Y(_13899_));
 sky130_fd_sc_hd__inv_1 _20750_ (.A(_12601_),
    .Y(_13911_));
 sky130_fd_sc_hd__inv_1 _20751_ (.A(_12606_),
    .Y(_13918_));
 sky130_fd_sc_hd__inv_1 _20752_ (.A(_12611_),
    .Y(_13925_));
 sky130_fd_sc_hd__inv_1 _20753_ (.A(_07013_),
    .Y(_13928_));
 sky130_fd_sc_hd__inv_1 _20754_ (.A(_12616_),
    .Y(_13932_));
 sky130_fd_sc_hd__inv_1 _20755_ (.A(_12636_),
    .Y(_13964_));
 sky130_fd_sc_hd__inv_1 _20756_ (.A(_12641_),
    .Y(_13971_));
 sky130_fd_sc_hd__nor2b_1 _20757_ (.A(net521),
    .B_N(\hash.CA2.a_dash[24] ),
    .Y(_13974_));
 sky130_fd_sc_hd__inv_1 _20758_ (.A(_12646_),
    .Y(_13978_));
 sky130_fd_sc_hd__inv_1 _20759_ (.A(_12651_),
    .Y(_13985_));
 sky130_fd_sc_hd__inv_1 _20760_ (.A(_12656_),
    .Y(_13992_));
 sky130_fd_sc_hd__inv_1 _20761_ (.A(_12661_),
    .Y(_13999_));
 sky130_fd_sc_hd__inv_1 _20762_ (.A(\hash.CA1.S1.X[1] ),
    .Y(_14022_));
 sky130_fd_sc_hd__xnor2_1 _20763_ (.A(_06731_),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_08361_));
 sky130_fd_sc_hd__xnor2_4 _20764_ (.A(_06896_),
    .B(_08361_),
    .Y(_14041_));
 sky130_fd_sc_hd__xnor2_1 _20765_ (.A(\hash.CA1.S1.X[9] ),
    .B(_06784_),
    .Y(_08362_));
 sky130_fd_sc_hd__xnor2_2 _20766_ (.A(_06903_),
    .B(_08362_),
    .Y(_14049_));
 sky130_fd_sc_hd__inv_1 _20767_ (.A(_12688_),
    .Y(_14052_));
 sky130_fd_sc_hd__xnor2_2 _20768_ (.A(\hash.CA1.S1.X[10] ),
    .B(_06792_),
    .Y(_08363_));
 sky130_fd_sc_hd__xnor2_4 _20769_ (.A(_06910_),
    .B(_08363_),
    .Y(_14058_));
 sky130_fd_sc_hd__inv_1 _20770_ (.A(_12693_),
    .Y(_14062_));
 sky130_fd_sc_hd__xnor2_1 _20771_ (.A(_06758_),
    .B(_06804_),
    .Y(_08364_));
 sky130_fd_sc_hd__xnor2_4 _20772_ (.A(_06917_),
    .B(_08364_),
    .Y(_14068_));
 sky130_fd_sc_hd__xor2_1 _20773_ (.A(\hash.CA1.S1.X[12] ),
    .B(_06816_),
    .X(_08365_));
 sky130_fd_sc_hd__xnor2_4 _20774_ (.A(_06922_),
    .B(_08365_),
    .Y(_14077_));
 sky130_fd_sc_hd__xnor2_1 _20775_ (.A(_13613_),
    .B(_06774_),
    .Y(_08366_));
 sky130_fd_sc_hd__xnor2_1 _20776_ (.A(_06839_),
    .B(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__nor2_1 _20777_ (.A(net524),
    .B(_08367_),
    .Y(_14085_));
 sky130_fd_sc_hd__mux2i_1 _20778_ (.A0(\hash.CA1.S1.X[1] ),
    .A1(_12536_),
    .S(_06830_),
    .Y(_08368_));
 sky130_fd_sc_hd__xnor2_1 _20779_ (.A(_06784_),
    .B(_08368_),
    .Y(_14093_));
 sky130_fd_sc_hd__inv_1 _20780_ (.A(_12713_),
    .Y(_14096_));
 sky130_fd_sc_hd__xnor2_1 _20781_ (.A(\hash.CA1.S1.X[2] ),
    .B(\hash.CA1.S1.X[15] ),
    .Y(_08369_));
 sky130_fd_sc_hd__xnor2_1 _20782_ (.A(\hash.CA1.S1.X[20] ),
    .B(_08369_),
    .Y(_14102_));
 sky130_fd_sc_hd__xnor2_1 _20783_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06804_),
    .Y(_08370_));
 sky130_fd_sc_hd__xnor2_1 _20784_ (.A(\hash.CA1.S1.X[21] ),
    .B(_08370_),
    .Y(_14111_));
 sky130_fd_sc_hd__inv_1 _20785_ (.A(_12723_),
    .Y(_14114_));
 sky130_fd_sc_hd__xnor2_1 _20786_ (.A(_06699_),
    .B(_06816_),
    .Y(_08371_));
 sky130_fd_sc_hd__xnor2_1 _20787_ (.A(_06854_),
    .B(_08371_),
    .Y(_14120_));
 sky130_fd_sc_hd__inv_1 _20788_ (.A(_12728_),
    .Y(_14124_));
 sky130_fd_sc_hd__xnor2_1 _20789_ (.A(_06707_),
    .B(\hash.CA1.S1.X[23] ),
    .Y(_08372_));
 sky130_fd_sc_hd__xnor2_2 _20790_ (.A(_06821_),
    .B(_08372_),
    .Y(_14130_));
 sky130_fd_sc_hd__xnor2_1 _20791_ (.A(_06713_),
    .B(_06830_),
    .Y(_08373_));
 sky130_fd_sc_hd__xnor2_1 _20792_ (.A(\hash.CA1.S1.X[24] ),
    .B(_08373_),
    .Y(_14139_));
 sky130_fd_sc_hd__xnor2_1 _20793_ (.A(\hash.CA1.S1.X[7] ),
    .B(\hash.CA1.S1.X[20] ),
    .Y(_08374_));
 sky130_fd_sc_hd__xnor2_1 _20794_ (.A(\hash.CA1.S1.X[25] ),
    .B(_08374_),
    .Y(_14147_));
 sky130_fd_sc_hd__inv_2 _20795_ (.A(_12743_),
    .Y(_14150_));
 sky130_fd_sc_hd__xnor2_1 _20796_ (.A(\hash.CA1.S1.X[8] ),
    .B(\hash.CA1.S1.X[21] ),
    .Y(_08375_));
 sky130_fd_sc_hd__xnor2_1 _20797_ (.A(\hash.CA1.S1.X[26] ),
    .B(_08375_),
    .Y(_14156_));
 sky130_fd_sc_hd__inv_1 _20798_ (.A(_12748_),
    .Y(_14160_));
 sky130_fd_sc_hd__xnor2_1 _20799_ (.A(_06738_),
    .B(_06854_),
    .Y(_08376_));
 sky130_fd_sc_hd__xnor2_1 _20800_ (.A(_06896_),
    .B(_08376_),
    .Y(_14166_));
 sky130_fd_sc_hd__xnor2_1 _20801_ (.A(\hash.CA1.S1.X[10] ),
    .B(_06864_),
    .Y(_08377_));
 sky130_fd_sc_hd__xnor2_1 _20802_ (.A(_06903_),
    .B(_08377_),
    .Y(_14175_));
 sky130_fd_sc_hd__xnor2_1 _20803_ (.A(_06758_),
    .B(\hash.CA1.S1.X[24] ),
    .Y(_08378_));
 sky130_fd_sc_hd__xnor2_1 _20804_ (.A(_06910_),
    .B(_08378_),
    .Y(_14183_));
 sky130_fd_sc_hd__xor2_1 _20805_ (.A(\hash.CA1.S1.X[12] ),
    .B(\hash.CA1.S1.X[25] ),
    .X(_08379_));
 sky130_fd_sc_hd__xnor2_1 _20806_ (.A(_06917_),
    .B(_08379_),
    .Y(_14191_));
 sky130_fd_sc_hd__xnor2_2 _20807_ (.A(\hash.CA1.S1.X[13] ),
    .B(\hash.CA1.S1.X[26] ),
    .Y(_08380_));
 sky130_fd_sc_hd__xnor2_1 _20808_ (.A(_06922_),
    .B(_08380_),
    .Y(_14199_));
 sky130_fd_sc_hd__mux2i_4 _20809_ (.A0(_13613_),
    .A1(_00781_),
    .S(_06896_),
    .Y(_08381_));
 sky130_fd_sc_hd__xnor2_4 _20810_ (.A(_06784_),
    .B(_08381_),
    .Y(_14207_));
 sky130_fd_sc_hd__inv_2 _20811_ (.A(_12778_),
    .Y(_14210_));
 sky130_fd_sc_hd__nand3_1 _20812_ (.A(_06210_),
    .B(_12536_),
    .C(_06902_),
    .Y(_08382_));
 sky130_fd_sc_hd__o21ai_2 _20813_ (.A1(_12536_),
    .A2(\hash.CA1.S1.X[28] ),
    .B1(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__xnor2_1 _20814_ (.A(_06792_),
    .B(_08383_),
    .Y(_14216_));
 sky130_fd_sc_hd__inv_1 _20815_ (.A(_12783_),
    .Y(_14220_));
 sky130_fd_sc_hd__xnor2_2 _20816_ (.A(_06688_),
    .B(_06804_),
    .Y(_08384_));
 sky130_fd_sc_hd__xnor2_1 _20817_ (.A(_06910_),
    .B(_08384_),
    .Y(_14226_));
 sky130_fd_sc_hd__inv_2 _20818_ (.A(_12788_),
    .Y(_14230_));
 sky130_fd_sc_hd__xnor2_2 _20819_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06816_),
    .Y(_08385_));
 sky130_fd_sc_hd__xnor2_1 _20820_ (.A(_06917_),
    .B(_08385_),
    .Y(_14236_));
 sky130_fd_sc_hd__inv_1 _20821_ (.A(_12793_),
    .Y(_14240_));
 sky130_fd_sc_hd__xnor2_2 _20822_ (.A(_06699_),
    .B(_06821_),
    .Y(_08386_));
 sky130_fd_sc_hd__xnor2_1 _20823_ (.A(_06922_),
    .B(_08386_),
    .Y(_14246_));
 sky130_fd_sc_hd__inv_1 _20824_ (.A(_12798_),
    .Y(_14250_));
 sky130_fd_sc_hd__nor2_1 _20825_ (.A(\hash.CA1.S1.X[0] ),
    .B(_06707_),
    .Y(_08387_));
 sky130_fd_sc_hd__a21oi_4 _20826_ (.A1(_13613_),
    .A2(_06707_),
    .B1(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__xor2_4 _20827_ (.A(_06830_),
    .B(_08388_),
    .X(_14256_));
 sky130_fd_sc_hd__mux2i_4 _20828_ (.A0(_12536_),
    .A1(\hash.CA1.S1.X[1] ),
    .S(\hash.CA1.S1.X[6] ),
    .Y(_08389_));
 sky130_fd_sc_hd__xor2_2 _20829_ (.A(\hash.CA1.S1.X[20] ),
    .B(_08389_),
    .X(_14265_));
 sky130_fd_sc_hd__inv_1 _20830_ (.A(_12808_),
    .Y(_14268_));
 sky130_fd_sc_hd__xnor2_2 _20831_ (.A(\hash.CA1.S1.X[2] ),
    .B(\hash.CA1.S1.X[7] ),
    .Y(_08390_));
 sky130_fd_sc_hd__xnor2_4 _20832_ (.A(\hash.CA1.S1.X[21] ),
    .B(_08390_),
    .Y(_14274_));
 sky130_fd_sc_hd__inv_1 _20833_ (.A(_12813_),
    .Y(_14278_));
 sky130_fd_sc_hd__xnor2_4 _20834_ (.A(_06692_),
    .B(_06731_),
    .Y(_08391_));
 sky130_fd_sc_hd__xnor2_2 _20835_ (.A(_06854_),
    .B(_08391_),
    .Y(_14284_));
 sky130_fd_sc_hd__xnor2_2 _20836_ (.A(_06699_),
    .B(_06738_),
    .Y(_08392_));
 sky130_fd_sc_hd__xnor2_2 _20837_ (.A(\hash.CA1.S1.X[23] ),
    .B(_08392_),
    .Y(_14293_));
 sky130_fd_sc_hd__inv_1 _20838_ (.A(_12823_),
    .Y(_14296_));
 sky130_fd_sc_hd__inv_1 _20839_ (.A(_12844_),
    .Y(_14300_));
 sky130_fd_sc_hd__inv_1 _20840_ (.A(_12849_),
    .Y(_14304_));
 sky130_fd_sc_hd__inv_1 _20841_ (.A(_12854_),
    .Y(_14308_));
 sky130_fd_sc_hd__inv_1 _20842_ (.A(_12861_),
    .Y(_14312_));
 sky130_fd_sc_hd__inv_1 _20843_ (.A(_12870_),
    .Y(_14316_));
 sky130_fd_sc_hd__inv_1 _20844_ (.A(_12878_),
    .Y(_14320_));
 sky130_fd_sc_hd__inv_1 _20845_ (.A(_12883_),
    .Y(_14324_));
 sky130_fd_sc_hd__inv_1 _20846_ (.A(_12888_),
    .Y(_12890_));
 sky130_fd_sc_hd__inv_1 _20847_ (.A(_12896_),
    .Y(_12898_));
 sky130_fd_sc_hd__inv_1 _20848_ (.A(_12925_),
    .Y(_12926_));
 sky130_fd_sc_hd__inv_1 _20849_ (.A(_12932_),
    .Y(_12934_));
 sky130_fd_sc_hd__inv_1 _20850_ (.A(_12967_),
    .Y(_12968_));
 sky130_fd_sc_hd__inv_1 _20851_ (.A(_12983_),
    .Y(_12984_));
 sky130_fd_sc_hd__inv_1 _20852_ (.A(_12999_),
    .Y(_13000_));
 sky130_fd_sc_hd__inv_1 _20853_ (.A(_13049_),
    .Y(_14370_));
 sky130_fd_sc_hd__xor2_2 _20854_ (.A(_12281_),
    .B(_06258_),
    .X(_08393_));
 sky130_fd_sc_hd__xnor2_4 _20855_ (.A(_06349_),
    .B(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__nor2_1 _20856_ (.A(net520),
    .B(_08394_),
    .Y(_14374_));
 sky130_fd_sc_hd__inv_1 _20857_ (.A(_12835_),
    .Y(_14377_));
 sky130_fd_sc_hd__inv_1 _20858_ (.A(_12545_),
    .Y(\hash.CA1.p4[0] ));
 sky130_fd_sc_hd__inv_1 _20859_ (.A(_13400_),
    .Y(_12247_));
 sky130_fd_sc_hd__inv_1 _20860_ (.A(_14024_),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_1 _20861_ (.A(_13713_),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_1 _20862_ (.A(\hash.CA1.p4[1] ),
    .Y(_13064_));
 sky130_fd_sc_hd__inv_1 _20863_ (.A(_14018_),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_1 _20864_ (.A(_14021_),
    .Y(_00824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_976 ();
 sky130_fd_sc_hd__nor2_1 _20866_ (.A(net762),
    .B(\count15_1[1] ),
    .Y(_00907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_975 ();
 sky130_fd_sc_hd__nor2b_1 _20868_ (.A(net762),
    .B_N(_00645_),
    .Y(_00908_));
 sky130_fd_sc_hd__xnor2_1 _20869_ (.A(\count15_1[3] ),
    .B(_13689_),
    .Y(_08397_));
 sky130_fd_sc_hd__nor2_1 _20870_ (.A(net762),
    .B(_08397_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand3_1 _20871_ (.A(net701),
    .B(net696),
    .C(\count15_1[3] ),
    .Y(_08398_));
 sky130_fd_sc_hd__xor2_1 _20872_ (.A(\count15_1[4] ),
    .B(_08398_),
    .X(_08399_));
 sky130_fd_sc_hd__nor2_1 _20873_ (.A(net762),
    .B(_08399_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand3_1 _20874_ (.A(\count15_1[3] ),
    .B(\count15_1[4] ),
    .C(_13689_),
    .Y(_08400_));
 sky130_fd_sc_hd__xor2_1 _20875_ (.A(\count15_1[5] ),
    .B(_08400_),
    .X(_08401_));
 sky130_fd_sc_hd__nor2_1 _20876_ (.A(net762),
    .B(_08401_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _20877_ (.A(_09893_),
    .B(\count15_2[1] ),
    .Y(_00912_));
 sky130_fd_sc_hd__nor2b_1 _20878_ (.A(net762),
    .B_N(_00649_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_1 _20879_ (.A(\count15_2[3] ),
    .B(_13693_),
    .Y(_08402_));
 sky130_fd_sc_hd__nor2_1 _20880_ (.A(net762),
    .B(_08402_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand3_1 _20881_ (.A(net682),
    .B(net677),
    .C(\count15_2[3] ),
    .Y(_08403_));
 sky130_fd_sc_hd__xor2_1 _20882_ (.A(\count15_2[4] ),
    .B(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__nor2_1 _20883_ (.A(net762),
    .B(_08404_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand3_1 _20884_ (.A(\count15_2[3] ),
    .B(\count15_2[4] ),
    .C(_13693_),
    .Y(_08405_));
 sky130_fd_sc_hd__xor2_1 _20885_ (.A(\count15_2[5] ),
    .B(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__nor2_1 _20886_ (.A(net762),
    .B(_08406_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_1 _20887_ (.A(net762),
    .B(\count16_1[1] ),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2b_1 _20888_ (.A(net762),
    .B_N(_00646_),
    .Y(_00918_));
 sky130_fd_sc_hd__xnor2_1 _20889_ (.A(\count16_1[3] ),
    .B(_13690_),
    .Y(_08407_));
 sky130_fd_sc_hd__nor2_1 _20890_ (.A(net762),
    .B(_08407_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand3_1 _20891_ (.A(net663),
    .B(\count16_1[2] ),
    .C(net653),
    .Y(_08408_));
 sky130_fd_sc_hd__xor2_1 _20892_ (.A(\count16_1[4] ),
    .B(_08408_),
    .X(_08409_));
 sky130_fd_sc_hd__nor2_1 _20893_ (.A(net762),
    .B(_08409_),
    .Y(_00920_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_974 ();
 sky130_fd_sc_hd__nand3_1 _20895_ (.A(\count16_1[3] ),
    .B(\count16_1[4] ),
    .C(_13690_),
    .Y(_08411_));
 sky130_fd_sc_hd__xor2_1 _20896_ (.A(\count16_1[5] ),
    .B(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__nor2_1 _20897_ (.A(net762),
    .B(_08412_),
    .Y(_00921_));
 sky130_fd_sc_hd__nor2_1 _20898_ (.A(net762),
    .B(\count16_2[1] ),
    .Y(_00922_));
 sky130_fd_sc_hd__nor2b_1 _20899_ (.A(net762),
    .B_N(_00650_),
    .Y(_00923_));
 sky130_fd_sc_hd__xnor2_1 _20900_ (.A(\count16_2[3] ),
    .B(_13694_),
    .Y(_08413_));
 sky130_fd_sc_hd__nor2_1 _20901_ (.A(net762),
    .B(_08413_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand3_1 _20902_ (.A(net642),
    .B(\count16_2[2] ),
    .C(\count16_2[3] ),
    .Y(_08414_));
 sky130_fd_sc_hd__xor2_1 _20903_ (.A(\count16_2[4] ),
    .B(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__nor2_1 _20904_ (.A(net762),
    .B(_08415_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand3_1 _20905_ (.A(\count16_2[3] ),
    .B(\count16_2[4] ),
    .C(_13694_),
    .Y(_08416_));
 sky130_fd_sc_hd__xor2_1 _20906_ (.A(\count16_2[5] ),
    .B(_08416_),
    .X(_08417_));
 sky130_fd_sc_hd__nor2_1 _20907_ (.A(net762),
    .B(_08417_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_1 _20908_ (.A(_09893_),
    .B(\count2_1[1] ),
    .Y(_00927_));
 sky130_fd_sc_hd__or2_0 _20909_ (.A(net762),
    .B(_00643_),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_1 _20910_ (.A(\count2_1[3] ),
    .B(_13714_),
    .Y(_08418_));
 sky130_fd_sc_hd__nand2_1 _20911_ (.A(_09893_),
    .B(_08418_),
    .Y(_00929_));
 sky130_fd_sc_hd__nand3_1 _20912_ (.A(\count2_1[1] ),
    .B(\count2_1[2] ),
    .C(\count2_1[3] ),
    .Y(_08419_));
 sky130_fd_sc_hd__xor2_1 _20913_ (.A(\count2_1[4] ),
    .B(_08419_),
    .X(_08420_));
 sky130_fd_sc_hd__nor2_1 _20914_ (.A(net762),
    .B(_08420_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand3_1 _20915_ (.A(\count2_1[3] ),
    .B(net614),
    .C(_13714_),
    .Y(_08421_));
 sky130_fd_sc_hd__xor2_1 _20916_ (.A(\count2_1[5] ),
    .B(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__nor2_1 _20917_ (.A(net762),
    .B(_08422_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _20918_ (.A(_09893_),
    .B(\count2_2[1] ),
    .Y(_00932_));
 sky130_fd_sc_hd__or2_0 _20919_ (.A(net762),
    .B(_00647_),
    .X(_00933_));
 sky130_fd_sc_hd__xnor2_1 _20920_ (.A(net598),
    .B(_13691_),
    .Y(_08423_));
 sky130_fd_sc_hd__nand2_1 _20921_ (.A(_09893_),
    .B(_08423_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand3_1 _20922_ (.A(\count2_2[1] ),
    .B(\count2_2[2] ),
    .C(\count2_2[3] ),
    .Y(_08424_));
 sky130_fd_sc_hd__xor2_1 _20923_ (.A(\count2_2[4] ),
    .B(_08424_),
    .X(_08425_));
 sky130_fd_sc_hd__nor2_1 _20924_ (.A(net762),
    .B(_08425_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand3_1 _20925_ (.A(net598),
    .B(\count2_2[4] ),
    .C(_13691_),
    .Y(_08426_));
 sky130_fd_sc_hd__xor2_1 _20926_ (.A(\count2_2[5] ),
    .B(_08426_),
    .X(_08427_));
 sky130_fd_sc_hd__nor2_1 _20927_ (.A(net762),
    .B(_08427_),
    .Y(_00936_));
 sky130_fd_sc_hd__nor2_1 _20928_ (.A(net762),
    .B(\count7_1[1] ),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2b_1 _20929_ (.A(net762),
    .B_N(_00644_),
    .Y(_00938_));
 sky130_fd_sc_hd__xnor2_1 _20930_ (.A(net579),
    .B(_13688_),
    .Y(_08428_));
 sky130_fd_sc_hd__nand2_1 _20931_ (.A(_09893_),
    .B(_08428_),
    .Y(_00939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_973 ();
 sky130_fd_sc_hd__nand3_1 _20933_ (.A(net590),
    .B(\count7_1[2] ),
    .C(\count7_1[3] ),
    .Y(_08430_));
 sky130_fd_sc_hd__xor2_1 _20934_ (.A(\count7_1[4] ),
    .B(_08430_),
    .X(_08431_));
 sky130_fd_sc_hd__nor2_1 _20935_ (.A(net762),
    .B(_08431_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand3_1 _20936_ (.A(net579),
    .B(\count7_1[4] ),
    .C(_13688_),
    .Y(_08432_));
 sky130_fd_sc_hd__xor2_1 _20937_ (.A(\count7_1[5] ),
    .B(_08432_),
    .X(_08433_));
 sky130_fd_sc_hd__nor2_1 _20938_ (.A(net762),
    .B(_08433_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_1 _20939_ (.A(_09893_),
    .B(\count7_2[1] ),
    .Y(_00942_));
 sky130_fd_sc_hd__nor2b_1 _20940_ (.A(net762),
    .B_N(_00648_),
    .Y(_00943_));
 sky130_fd_sc_hd__xnor2_1 _20941_ (.A(\count7_2[3] ),
    .B(_13692_),
    .Y(_08434_));
 sky130_fd_sc_hd__nand2_1 _20942_ (.A(_09893_),
    .B(_08434_),
    .Y(_00944_));
 sky130_fd_sc_hd__nand3_1 _20943_ (.A(net572),
    .B(\count7_2[2] ),
    .C(\count7_2[3] ),
    .Y(_08435_));
 sky130_fd_sc_hd__xor2_1 _20944_ (.A(\count7_2[4] ),
    .B(_08435_),
    .X(_08436_));
 sky130_fd_sc_hd__nor2_1 _20945_ (.A(net762),
    .B(_08436_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand3_1 _20946_ (.A(\count7_2[3] ),
    .B(net556),
    .C(_13692_),
    .Y(_08437_));
 sky130_fd_sc_hd__xor2_1 _20947_ (.A(\count7_2[5] ),
    .B(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__nor2_1 _20948_ (.A(net762),
    .B(_08438_),
    .Y(_00946_));
 sky130_fd_sc_hd__xnor2_1 _20949_ (.A(_00651_),
    .B(_00128_),
    .Y(_08439_));
 sky130_fd_sc_hd__nor2_1 _20950_ (.A(net762),
    .B(_08439_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _20951_ (.A(\count_1[2] ),
    .B(_00128_),
    .Y(_08440_));
 sky130_fd_sc_hd__nand2_1 _20952_ (.A(_00652_),
    .B(_09890_),
    .Y(_08441_));
 sky130_fd_sc_hd__a21oi_1 _20953_ (.A1(_08440_),
    .A2(_08441_),
    .B1(net762),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _20954_ (.A(_13701_),
    .B(_09890_),
    .Y(_08442_));
 sky130_fd_sc_hd__xor2_1 _20955_ (.A(\count_1[3] ),
    .B(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__nor2_1 _20956_ (.A(net762),
    .B(_08443_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand4_1 _20957_ (.A(\count_1[3] ),
    .B(\count_1[2] ),
    .C(\count_1[1] ),
    .D(_09890_),
    .Y(_08444_));
 sky130_fd_sc_hd__xor2_1 _20958_ (.A(\count_1[4] ),
    .B(_08444_),
    .X(_08445_));
 sky130_fd_sc_hd__nand2_1 _20959_ (.A(_09893_),
    .B(_08445_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand4_1 _20960_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C(_13701_),
    .D(_09890_),
    .Y(_08446_));
 sky130_fd_sc_hd__xor2_1 _20961_ (.A(\count_1[5] ),
    .B(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__nor2_1 _20962_ (.A(net762),
    .B(_08447_),
    .Y(_00951_));
 sky130_fd_sc_hd__xnor2_1 _20963_ (.A(_00653_),
    .B(_00128_),
    .Y(_08448_));
 sky130_fd_sc_hd__nor2_1 _20964_ (.A(net762),
    .B(_08448_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand2_1 _20965_ (.A(\count_2[2] ),
    .B(_00128_),
    .Y(_08449_));
 sky130_fd_sc_hd__nand2_1 _20966_ (.A(_00654_),
    .B(_09890_),
    .Y(_08450_));
 sky130_fd_sc_hd__a21oi_1 _20967_ (.A1(_08449_),
    .A2(_08450_),
    .B1(net762),
    .Y(_00953_));
 sky130_fd_sc_hd__xnor2_1 _20968_ (.A(\count_2[3] ),
    .B(_13709_),
    .Y(_08451_));
 sky130_fd_sc_hd__a21oi_1 _20969_ (.A1(_09890_),
    .A2(_08451_),
    .B1(net762),
    .Y(_00954_));
 sky130_fd_sc_hd__nand3_1 _20970_ (.A(\count_2[3] ),
    .B(\count_2[2] ),
    .C(\count_2[1] ),
    .Y(_08452_));
 sky130_fd_sc_hd__xor2_1 _20971_ (.A(\count_2[4] ),
    .B(_08452_),
    .X(_08453_));
 sky130_fd_sc_hd__nand3_1 _20972_ (.A(_09893_),
    .B(_09890_),
    .C(_08453_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand3_1 _20973_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_13709_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand2_1 _20974_ (.A(\count_2[6] ),
    .B(\count_2[5] ),
    .Y(_08455_));
 sky130_fd_sc_hd__nor2_1 _20975_ (.A(_08454_),
    .B(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__a211oi_1 _20976_ (.A1(_09963_),
    .A2(_08454_),
    .B1(_08456_),
    .C1(net762),
    .Y(_00956_));
 sky130_fd_sc_hd__nor2b_1 _20977_ (.A(\count_2[6] ),
    .B_N(_09889_),
    .Y(_08457_));
 sky130_fd_sc_hd__nand2_1 _20978_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .Y(_08458_));
 sky130_fd_sc_hd__nor2_1 _20979_ (.A(_08452_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__mux2i_1 _20980_ (.A0(\count_2[6] ),
    .A1(_08457_),
    .S(_08459_),
    .Y(_08460_));
 sky130_fd_sc_hd__nor2_1 _20981_ (.A(net762),
    .B(_08460_),
    .Y(_00957_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_972 ();
 sky130_fd_sc_hd__nor2_4 _20983_ (.A(\count_hash1[6] ),
    .B(_10033_),
    .Y(_08462_));
 sky130_fd_sc_hd__xnor2_1 _20984_ (.A(_00642_),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nor2_1 _20985_ (.A(net525),
    .B(_08463_),
    .Y(_00958_));
 sky130_fd_sc_hd__nand2_1 _20986_ (.A(\count_hash1[2] ),
    .B(_08462_),
    .Y(_08464_));
 sky130_fd_sc_hd__or2_4 _20987_ (.A(\count_hash1[6] ),
    .B(_10033_),
    .X(_08465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_971 ();
 sky130_fd_sc_hd__nand2_1 _20989_ (.A(_00655_),
    .B(_08465_),
    .Y(_08467_));
 sky130_fd_sc_hd__a21oi_1 _20990_ (.A1(_08464_),
    .A2(_08467_),
    .B1(net525),
    .Y(_00959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_970 ();
 sky130_fd_sc_hd__a21oi_1 _20992_ (.A1(net492),
    .A2(_08465_),
    .B1(net525),
    .Y(_00960_));
 sky130_fd_sc_hd__a21oi_1 _20993_ (.A1(net499),
    .A2(_08465_),
    .B1(net525),
    .Y(_00961_));
 sky130_fd_sc_hd__a21oi_1 _20994_ (.A1(_10508_),
    .A2(_08465_),
    .B1(net525),
    .Y(_00962_));
 sky130_fd_sc_hd__and3_1 _20995_ (.A(\count_hash1[5] ),
    .B(\count_hash1[2] ),
    .C(\count_hash1[1] ),
    .X(_08469_));
 sky130_fd_sc_hd__nand3_1 _20996_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__xor2_1 _20997_ (.A(\count_hash1[6] ),
    .B(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__nor3_1 _20998_ (.A(net525),
    .B(_08462_),
    .C(_08471_),
    .Y(_00963_));
 sky130_fd_sc_hd__xnor2_1 _20999_ (.A(_00656_),
    .B(_08462_),
    .Y(_08472_));
 sky130_fd_sc_hd__nor2_1 _21000_ (.A(net525),
    .B(_08472_),
    .Y(_00964_));
 sky130_fd_sc_hd__nand2_1 _21001_ (.A(\count_hash2[2] ),
    .B(_08462_),
    .Y(_08473_));
 sky130_fd_sc_hd__nand2_1 _21002_ (.A(_00657_),
    .B(_08465_),
    .Y(_08474_));
 sky130_fd_sc_hd__a21oi_1 _21003_ (.A1(_08473_),
    .A2(_08474_),
    .B1(net525),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _21004_ (.A(_13076_),
    .B(_08465_),
    .Y(_08475_));
 sky130_fd_sc_hd__xor2_1 _21005_ (.A(\count_hash2[3] ),
    .B(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__nor2_1 _21006_ (.A(net525),
    .B(_08476_),
    .Y(_00966_));
 sky130_fd_sc_hd__o21ai_0 _21007_ (.A1(_10015_),
    .A2(_08462_),
    .B1(\count_hash2[4] ),
    .Y(_08477_));
 sky130_fd_sc_hd__or3_1 _21008_ (.A(\count_hash2[4] ),
    .B(_10015_),
    .C(_08462_),
    .X(_08478_));
 sky130_fd_sc_hd__a21oi_1 _21009_ (.A1(_08477_),
    .A2(_08478_),
    .B1(net525),
    .Y(_00967_));
 sky130_fd_sc_hd__o21ai_0 _21010_ (.A1(_10026_),
    .A2(_08462_),
    .B1(\count_hash2[5] ),
    .Y(_08479_));
 sky130_fd_sc_hd__or3_1 _21011_ (.A(\count_hash2[5] ),
    .B(_10026_),
    .C(_08462_),
    .X(_08480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_969 ();
 sky130_fd_sc_hd__a21oi_1 _21013_ (.A1(_08479_),
    .A2(_08480_),
    .B1(net525),
    .Y(_00968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_967 ();
 sky130_fd_sc_hd__nor2_2 _21016_ (.A(_13079_),
    .B(_13084_),
    .Y(_08484_));
 sky130_fd_sc_hd__nor3_2 _21017_ (.A(_10564_),
    .B(_10575_),
    .C(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__nor2_4 _21018_ (.A(_13084_),
    .B(_13086_),
    .Y(_08486_));
 sky130_fd_sc_hd__nand2_4 _21019_ (.A(_10503_),
    .B(net507),
    .Y(_08487_));
 sky130_fd_sc_hd__nor3_1 _21020_ (.A(net463),
    .B(_08486_),
    .C(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__nor2_2 _21021_ (.A(_08485_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_964 ();
 sky130_fd_sc_hd__nand2_1 _21025_ (.A(net507),
    .B(net459),
    .Y(_08493_));
 sky130_fd_sc_hd__inv_2 _21026_ (.A(_13086_),
    .Y(_08494_));
 sky130_fd_sc_hd__nor2_2 _21027_ (.A(_08494_),
    .B(net507),
    .Y(_08495_));
 sky130_fd_sc_hd__a22o_1 _21028_ (.A1(_13084_),
    .A2(_08493_),
    .B1(_08495_),
    .B2(net463),
    .X(_08496_));
 sky130_fd_sc_hd__nor2_4 _21029_ (.A(_10512_),
    .B(net463),
    .Y(_08497_));
 sky130_fd_sc_hd__nand2_4 _21030_ (.A(_10512_),
    .B(net459),
    .Y(_08498_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_963 ();
 sky130_fd_sc_hd__clkinvlp_4 _21032_ (.A(_13080_),
    .Y(_08500_));
 sky130_fd_sc_hd__a21oi_1 _21033_ (.A1(_10532_),
    .A2(_08498_),
    .B1(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__a221oi_1 _21034_ (.A1(_10512_),
    .A2(_08496_),
    .B1(_08497_),
    .B2(_08495_),
    .C1(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__nor2_8 _21035_ (.A(_10503_),
    .B(net507),
    .Y(_08503_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_962 ();
 sky130_fd_sc_hd__nor2_2 _21037_ (.A(net461),
    .B(_10575_),
    .Y(_08505_));
 sky130_fd_sc_hd__o21ai_1 _21038_ (.A1(_13079_),
    .A2(_13080_),
    .B1(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__nor2_1 _21039_ (.A(_13080_),
    .B(_13086_),
    .Y(_08507_));
 sky130_fd_sc_hd__nor2_2 _21040_ (.A(net461),
    .B(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__nand2_1 _21041_ (.A(_08503_),
    .B(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__nand2_1 _21042_ (.A(_08506_),
    .B(_08509_),
    .Y(_08510_));
 sky130_fd_sc_hd__nand2_1 _21043_ (.A(_13079_),
    .B(_08503_),
    .Y(_08511_));
 sky130_fd_sc_hd__o21ai_0 _21044_ (.A1(_13084_),
    .A2(_13086_),
    .B1(_10513_),
    .Y(_08512_));
 sky130_fd_sc_hd__a21oi_2 _21045_ (.A1(_08511_),
    .A2(_08512_),
    .B1(net463),
    .Y(_08513_));
 sky130_fd_sc_hd__a311oi_4 _21046_ (.A1(_13084_),
    .A2(net459),
    .A3(_08503_),
    .B1(_08510_),
    .C1(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__nor2_4 _21047_ (.A(_10503_),
    .B(net459),
    .Y(_08515_));
 sky130_fd_sc_hd__nor2_1 _21048_ (.A(_13079_),
    .B(_13080_),
    .Y(_08516_));
 sky130_fd_sc_hd__o22ai_2 _21049_ (.A1(net463),
    .A2(_08486_),
    .B1(_08515_),
    .B2(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__nor2_4 _21050_ (.A(_10503_),
    .B(net490),
    .Y(_08518_));
 sky130_fd_sc_hd__or2_2 _21051_ (.A(_13080_),
    .B(_13084_),
    .X(_08519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_961 ();
 sky130_fd_sc_hd__a22oi_1 _21053_ (.A1(_13086_),
    .A2(_08503_),
    .B1(_08518_),
    .B2(_08519_),
    .Y(_08521_));
 sky130_fd_sc_hd__nor3_1 _21054_ (.A(_13079_),
    .B(_13080_),
    .C(_13084_),
    .Y(_08522_));
 sky130_fd_sc_hd__nand2_1 _21055_ (.A(_10512_),
    .B(net461),
    .Y(_08523_));
 sky130_fd_sc_hd__or3_2 _21056_ (.A(net507),
    .B(_08522_),
    .C(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__o21ai_2 _21057_ (.A1(net459),
    .A2(_08521_),
    .B1(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__a21oi_1 _21058_ (.A1(net507),
    .A2(_08517_),
    .B1(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__nand2_1 _21059_ (.A(_13079_),
    .B(_10512_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand2_1 _21060_ (.A(_13084_),
    .B(_10503_),
    .Y(_08528_));
 sky130_fd_sc_hd__a31oi_1 _21061_ (.A1(_08494_),
    .A2(_08527_),
    .A3(_08528_),
    .B1(_10532_),
    .Y(_08529_));
 sky130_fd_sc_hd__nor2_1 _21062_ (.A(_10575_),
    .B(_08522_),
    .Y(_08530_));
 sky130_fd_sc_hd__o21ai_1 _21063_ (.A1(_08529_),
    .A2(_08530_),
    .B1(net461),
    .Y(_08531_));
 sky130_fd_sc_hd__and3_4 _21064_ (.A(_08514_),
    .B(_08526_),
    .C(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_960 ();
 sky130_fd_sc_hd__nand2b_4 _21066_ (.A_N(_08532_),
    .B(_10573_),
    .Y(_08534_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_958 ();
 sky130_fd_sc_hd__a21oi_2 _21069_ (.A1(_08489_),
    .A2(_08502_),
    .B1(_08534_),
    .Y(_00969_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_957 ();
 sky130_fd_sc_hd__nor2_1 _21071_ (.A(_08500_),
    .B(_10512_),
    .Y(_08538_));
 sky130_fd_sc_hd__a21oi_1 _21072_ (.A1(_13084_),
    .A2(_10512_),
    .B1(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__nor3_1 _21073_ (.A(_10512_),
    .B(net503),
    .C(net459),
    .Y(_08540_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_956 ();
 sky130_fd_sc_hd__nand2_2 _21075_ (.A(net503),
    .B(net461),
    .Y(_08542_));
 sky130_fd_sc_hd__a21oi_1 _21076_ (.A1(_13084_),
    .A2(_08542_),
    .B1(_10503_),
    .Y(_08543_));
 sky130_fd_sc_hd__nand2_1 _21077_ (.A(net507),
    .B(_08497_),
    .Y(_08544_));
 sky130_fd_sc_hd__a21oi_1 _21078_ (.A1(_13084_),
    .A2(_08544_),
    .B1(_13080_),
    .Y(_08545_));
 sky130_fd_sc_hd__nor3_1 _21079_ (.A(_10513_),
    .B(_08543_),
    .C(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__nor2_1 _21080_ (.A(_13079_),
    .B(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__a311oi_1 _21081_ (.A1(net503),
    .A2(net459),
    .A3(_08539_),
    .B1(_08540_),
    .C1(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__nor2_8 _21082_ (.A(\count_hash1[6] ),
    .B(_10034_),
    .Y(_08549_));
 sky130_fd_sc_hd__o21ai_0 _21083_ (.A1(_08532_),
    .A2(_08548_),
    .B1(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__nand2b_1 _21084_ (.A_N(net525),
    .B(_08550_),
    .Y(_00970_));
 sky130_fd_sc_hd__nor2_1 _21085_ (.A(_10512_),
    .B(_10532_),
    .Y(_08551_));
 sky130_fd_sc_hd__nand2_1 _21086_ (.A(net463),
    .B(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_955 ();
 sky130_fd_sc_hd__a31oi_1 _21088_ (.A1(_13080_),
    .A2(_10564_),
    .A3(_08503_),
    .B1(_08532_),
    .Y(_08554_));
 sky130_fd_sc_hd__o21ai_1 _21089_ (.A1(_08486_),
    .A2(_08552_),
    .B1(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__nand2_2 _21090_ (.A(net463),
    .B(_08503_),
    .Y(_08556_));
 sky130_fd_sc_hd__o21ai_0 _21091_ (.A1(_08494_),
    .A2(_08556_),
    .B1(_08524_),
    .Y(_08557_));
 sky130_fd_sc_hd__nand2_1 _21092_ (.A(_10512_),
    .B(net507),
    .Y(_08558_));
 sky130_fd_sc_hd__nand2_2 _21093_ (.A(_10575_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__a222oi_1 _21094_ (.A1(_13084_),
    .A2(_10512_),
    .B1(_10513_),
    .B2(_08495_),
    .C1(_08559_),
    .C2(_13079_),
    .Y(_08560_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_954 ();
 sky130_fd_sc_hd__a22oi_1 _21096_ (.A1(_13084_),
    .A2(_08515_),
    .B1(_08497_),
    .B2(_13079_),
    .Y(_08562_));
 sky130_fd_sc_hd__nand2_1 _21097_ (.A(_13080_),
    .B(_10564_),
    .Y(_08563_));
 sky130_fd_sc_hd__nand2_1 _21098_ (.A(_13079_),
    .B(net463),
    .Y(_08564_));
 sky130_fd_sc_hd__a21oi_1 _21099_ (.A1(_08563_),
    .A2(_08564_),
    .B1(_10575_),
    .Y(_08565_));
 sky130_fd_sc_hd__nor2_1 _21100_ (.A(_08488_),
    .B(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__o221ai_1 _21101_ (.A1(net463),
    .A2(_08560_),
    .B1(_08562_),
    .B2(_10532_),
    .C1(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__nor3_1 _21102_ (.A(_08555_),
    .B(_08557_),
    .C(_08567_),
    .Y(_08568_));
 sky130_fd_sc_hd__o21bai_1 _21103_ (.A1(_10571_),
    .A2(_08568_),
    .B1_N(net525),
    .Y(_00971_));
 sky130_fd_sc_hd__nand2_1 _21104_ (.A(_13079_),
    .B(_10513_),
    .Y(_08569_));
 sky130_fd_sc_hd__nor2_1 _21105_ (.A(net459),
    .B(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__nand2_1 _21106_ (.A(_13080_),
    .B(_08551_),
    .Y(_08571_));
 sky130_fd_sc_hd__nor2_1 _21107_ (.A(net463),
    .B(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__nor2_1 _21108_ (.A(_08570_),
    .B(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_953 ();
 sky130_fd_sc_hd__nand3_1 _21110_ (.A(_13084_),
    .B(net459),
    .C(_10513_),
    .Y(_08575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_951 ();
 sky130_fd_sc_hd__nor2_1 _21113_ (.A(_13079_),
    .B(net461),
    .Y(_08578_));
 sky130_fd_sc_hd__nor2_1 _21114_ (.A(_10503_),
    .B(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_950 ();
 sky130_fd_sc_hd__nor2_1 _21116_ (.A(_10532_),
    .B(_08497_),
    .Y(_08581_));
 sky130_fd_sc_hd__o221ai_4 _21117_ (.A1(_13086_),
    .A2(_08523_),
    .B1(_08579_),
    .B2(_13084_),
    .C1(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__a41oi_1 _21118_ (.A1(_08511_),
    .A2(_08573_),
    .A3(_08575_),
    .A4(_08582_),
    .B1(_08534_),
    .Y(_00972_));
 sky130_fd_sc_hd__a22o_1 _21119_ (.A1(_13079_),
    .A2(_08518_),
    .B1(_08519_),
    .B2(_08503_),
    .X(_08583_));
 sky130_fd_sc_hd__a21oi_1 _21120_ (.A1(net461),
    .A2(_08583_),
    .B1(_08532_),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_2 _21121_ (.A(_13084_),
    .B(_10513_),
    .Y(_08585_));
 sky130_fd_sc_hd__nand2_1 _21122_ (.A(_08511_),
    .B(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__nand2_1 _21123_ (.A(_13086_),
    .B(_08503_),
    .Y(_08587_));
 sky130_fd_sc_hd__nand2_1 _21124_ (.A(_13080_),
    .B(_08518_),
    .Y(_08588_));
 sky130_fd_sc_hd__nand3_1 _21125_ (.A(net463),
    .B(_08587_),
    .C(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__o21ai_1 _21126_ (.A1(net463),
    .A2(_08586_),
    .B1(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_949 ();
 sky130_fd_sc_hd__nor3_1 _21128_ (.A(_13079_),
    .B(_13084_),
    .C(_10503_),
    .Y(_08592_));
 sky130_fd_sc_hd__a21oi_1 _21129_ (.A1(_10503_),
    .A2(_08486_),
    .B1(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__o21bai_1 _21130_ (.A1(_13080_),
    .A2(_08593_),
    .B1_N(_08493_),
    .Y(_08594_));
 sky130_fd_sc_hd__nor2_2 _21131_ (.A(net459),
    .B(_08487_),
    .Y(_08595_));
 sky130_fd_sc_hd__a21boi_0 _21132_ (.A1(_13086_),
    .A2(_08595_),
    .B1_N(_08569_),
    .Y(_08596_));
 sky130_fd_sc_hd__nand4_1 _21133_ (.A(_08584_),
    .B(_08590_),
    .C(_08594_),
    .D(_08596_),
    .Y(_08597_));
 sky130_fd_sc_hd__a21o_1 _21134_ (.A1(_08549_),
    .A2(_08597_),
    .B1(net525),
    .X(_00973_));
 sky130_fd_sc_hd__nand2_1 _21135_ (.A(_08489_),
    .B(_08582_),
    .Y(_08598_));
 sky130_fd_sc_hd__nor2_1 _21136_ (.A(_08510_),
    .B(_08598_),
    .Y(_08599_));
 sky130_fd_sc_hd__a21oi_1 _21137_ (.A1(_08590_),
    .A2(_08599_),
    .B1(_08534_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand2_1 _21138_ (.A(_08556_),
    .B(_08487_),
    .Y(_08600_));
 sky130_fd_sc_hd__a22oi_1 _21139_ (.A1(_13086_),
    .A2(_08595_),
    .B1(_08600_),
    .B2(_13079_),
    .Y(_08601_));
 sky130_fd_sc_hd__nand2_1 _21140_ (.A(net507),
    .B(_08498_),
    .Y(_08602_));
 sky130_fd_sc_hd__a21oi_1 _21141_ (.A1(_13084_),
    .A2(net507),
    .B1(_13086_),
    .Y(_08603_));
 sky130_fd_sc_hd__nor2_1 _21142_ (.A(_08498_),
    .B(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__a21oi_1 _21143_ (.A1(_13080_),
    .A2(_08602_),
    .B1(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__a31oi_1 _21144_ (.A1(_08489_),
    .A2(_08601_),
    .A3(_08605_),
    .B1(_08534_),
    .Y(_00975_));
 sky130_fd_sc_hd__o21ai_0 _21145_ (.A1(_13080_),
    .A2(net463),
    .B1(net507),
    .Y(_08606_));
 sky130_fd_sc_hd__nor2_1 _21146_ (.A(_13079_),
    .B(_08542_),
    .Y(_08607_));
 sky130_fd_sc_hd__nor2_2 _21147_ (.A(net507),
    .B(net463),
    .Y(_08608_));
 sky130_fd_sc_hd__a2111oi_2 _21148_ (.A1(_08494_),
    .A2(_08606_),
    .B1(_08607_),
    .C1(_08608_),
    .D1(_10503_),
    .Y(_08609_));
 sky130_fd_sc_hd__a31oi_1 _21149_ (.A1(_13084_),
    .A2(net463),
    .A3(_08503_),
    .B1(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__a32oi_4 _21150_ (.A1(_13080_),
    .A2(net463),
    .A3(_10513_),
    .B1(_08497_),
    .B2(_13086_),
    .Y(_08611_));
 sky130_fd_sc_hd__a31oi_1 _21151_ (.A1(_08601_),
    .A2(_08610_),
    .A3(_08611_),
    .B1(_08534_),
    .Y(_00976_));
 sky130_fd_sc_hd__a21oi_1 _21152_ (.A1(_10503_),
    .A2(_08542_),
    .B1(_13084_),
    .Y(_08612_));
 sky130_fd_sc_hd__nor2_1 _21153_ (.A(_08515_),
    .B(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__nor2_1 _21154_ (.A(_13086_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__a21oi_1 _21155_ (.A1(_13086_),
    .A2(_10575_),
    .B1(_08519_),
    .Y(_08615_));
 sky130_fd_sc_hd__nor2_1 _21156_ (.A(net459),
    .B(_08558_),
    .Y(_08616_));
 sky130_fd_sc_hd__o21ai_0 _21157_ (.A1(_08505_),
    .A2(_08616_),
    .B1(_13080_),
    .Y(_08617_));
 sky130_fd_sc_hd__o21ai_0 _21158_ (.A1(_08515_),
    .A2(_08497_),
    .B1(_13079_),
    .Y(_08618_));
 sky130_fd_sc_hd__o21ai_0 _21159_ (.A1(_13084_),
    .A2(_08495_),
    .B1(_08505_),
    .Y(_08619_));
 sky130_fd_sc_hd__o21ai_0 _21160_ (.A1(_10532_),
    .A2(_08618_),
    .B1(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__nor2_1 _21161_ (.A(_08532_),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__o311ai_2 _21162_ (.A1(_08608_),
    .A2(_08614_),
    .A3(_08615_),
    .B1(_08617_),
    .C1(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_948 ();
 sky130_fd_sc_hd__a21o_1 _21164_ (.A1(_08549_),
    .A2(_08622_),
    .B1(net525),
    .X(_00977_));
 sky130_fd_sc_hd__o21ai_0 _21165_ (.A1(_13086_),
    .A2(_08519_),
    .B1(_08503_),
    .Y(_08624_));
 sky130_fd_sc_hd__a21oi_1 _21166_ (.A1(_08569_),
    .A2(_08624_),
    .B1(net463),
    .Y(_08625_));
 sky130_fd_sc_hd__nor2_2 _21167_ (.A(_10503_),
    .B(net463),
    .Y(_08626_));
 sky130_fd_sc_hd__a21oi_1 _21168_ (.A1(_13084_),
    .A2(_08626_),
    .B1(_13086_),
    .Y(_08627_));
 sky130_fd_sc_hd__nor2_1 _21169_ (.A(_10532_),
    .B(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__nand2_1 _21170_ (.A(_13086_),
    .B(_10564_),
    .Y(_08629_));
 sky130_fd_sc_hd__nand2_1 _21171_ (.A(_13084_),
    .B(net463),
    .Y(_08630_));
 sky130_fd_sc_hd__o21ai_0 _21172_ (.A1(net507),
    .A2(net463),
    .B1(_13080_),
    .Y(_08631_));
 sky130_fd_sc_hd__a31oi_1 _21173_ (.A1(_08629_),
    .A2(_08630_),
    .A3(_08631_),
    .B1(_10512_),
    .Y(_08632_));
 sky130_fd_sc_hd__nor3_1 _21174_ (.A(_08625_),
    .B(_08628_),
    .C(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__nor2_1 _21175_ (.A(_08534_),
    .B(_08633_),
    .Y(_00978_));
 sky130_fd_sc_hd__a21oi_1 _21176_ (.A1(_08516_),
    .A2(_08486_),
    .B1(net463),
    .Y(_08634_));
 sky130_fd_sc_hd__a21oi_1 _21177_ (.A1(_08518_),
    .A2(_08634_),
    .B1(_08532_),
    .Y(_08635_));
 sky130_fd_sc_hd__nand2_1 _21178_ (.A(_10564_),
    .B(_08559_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_2 _21179_ (.A(_13079_),
    .B(_10503_),
    .Y(_08637_));
 sky130_fd_sc_hd__a21oi_2 _21180_ (.A1(_08585_),
    .A2(_08637_),
    .B1(net463),
    .Y(_08638_));
 sky130_fd_sc_hd__a31oi_1 _21181_ (.A1(_13080_),
    .A2(_08556_),
    .A3(_08636_),
    .B1(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__o21ai_1 _21182_ (.A1(net507),
    .A2(_08498_),
    .B1(_08552_),
    .Y(_08640_));
 sky130_fd_sc_hd__nor2_1 _21183_ (.A(_08494_),
    .B(_10532_),
    .Y(_08641_));
 sky130_fd_sc_hd__a21oi_1 _21184_ (.A1(_13084_),
    .A2(_10532_),
    .B1(_08641_),
    .Y(_08642_));
 sky130_fd_sc_hd__nand2_1 _21185_ (.A(_13079_),
    .B(_08608_),
    .Y(_08643_));
 sky130_fd_sc_hd__o21ai_0 _21186_ (.A1(_10564_),
    .A2(_08642_),
    .B1(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__a21oi_1 _21187_ (.A1(_08556_),
    .A2(_08544_),
    .B1(_08494_),
    .Y(_08645_));
 sky130_fd_sc_hd__a221oi_2 _21188_ (.A1(_13084_),
    .A2(_08640_),
    .B1(_08644_),
    .B2(_10512_),
    .C1(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__nand3_1 _21189_ (.A(_08635_),
    .B(_08639_),
    .C(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__a21o_1 _21190_ (.A1(_08549_),
    .A2(_08647_),
    .B1(net525),
    .X(_00979_));
 sky130_fd_sc_hd__a211o_1 _21191_ (.A1(_13080_),
    .A2(_10532_),
    .B1(_08641_),
    .C1(_13084_),
    .X(_08648_));
 sky130_fd_sc_hd__nand3_1 _21192_ (.A(net461),
    .B(_08518_),
    .C(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__o31ai_1 _21193_ (.A1(_08500_),
    .A2(net461),
    .A3(_10575_),
    .B1(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__o21ai_0 _21194_ (.A1(_13079_),
    .A2(_13084_),
    .B1(_10532_),
    .Y(_08651_));
 sky130_fd_sc_hd__a21oi_2 _21195_ (.A1(_08571_),
    .A2(_08651_),
    .B1(net459),
    .Y(_08652_));
 sky130_fd_sc_hd__nor2_1 _21196_ (.A(net490),
    .B(_08507_),
    .Y(_08653_));
 sky130_fd_sc_hd__o21ai_0 _21197_ (.A1(_13084_),
    .A2(_08653_),
    .B1(_08626_),
    .Y(_08654_));
 sky130_fd_sc_hd__o21ai_0 _21198_ (.A1(_08542_),
    .A2(_08637_),
    .B1(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__a2111oi_1 _21199_ (.A1(_08503_),
    .A2(_08508_),
    .B1(_08650_),
    .C1(_08652_),
    .D1(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__nor2_1 _21200_ (.A(_08534_),
    .B(_08656_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _21201_ (.A(_13086_),
    .B(_10503_),
    .Y(_08657_));
 sky130_fd_sc_hd__a221oi_1 _21202_ (.A1(_13080_),
    .A2(_10512_),
    .B1(_10575_),
    .B2(_13084_),
    .C1(net463),
    .Y(_08658_));
 sky130_fd_sc_hd__o21ai_1 _21203_ (.A1(_08494_),
    .A2(_08558_),
    .B1(_08585_),
    .Y(_08659_));
 sky130_fd_sc_hd__o21ai_0 _21204_ (.A1(_08484_),
    .A2(_08487_),
    .B1(_08587_),
    .Y(_08660_));
 sky130_fd_sc_hd__a2111oi_0 _21205_ (.A1(_13080_),
    .A2(_08558_),
    .B1(_08659_),
    .C1(_08660_),
    .D1(_10564_),
    .Y(_08661_));
 sky130_fd_sc_hd__a211oi_1 _21206_ (.A1(_08657_),
    .A2(_08658_),
    .B1(_08661_),
    .C1(_08534_),
    .Y(_00981_));
 sky130_fd_sc_hd__a21oi_1 _21207_ (.A1(net507),
    .A2(_08519_),
    .B1(_08495_),
    .Y(_08662_));
 sky130_fd_sc_hd__o22a_1 _21208_ (.A1(_08484_),
    .A2(_08552_),
    .B1(_08662_),
    .B2(_08498_),
    .X(_08663_));
 sky130_fd_sc_hd__a22oi_1 _21209_ (.A1(_13079_),
    .A2(_08505_),
    .B1(_08515_),
    .B2(_08648_),
    .Y(_08664_));
 sky130_fd_sc_hd__a31oi_2 _21210_ (.A1(_08611_),
    .A2(_08663_),
    .A3(_08664_),
    .B1(_08534_),
    .Y(_00982_));
 sky130_fd_sc_hd__a32oi_1 _21211_ (.A1(_13079_),
    .A2(net459),
    .A3(_10575_),
    .B1(_08616_),
    .B2(_13084_),
    .Y(_08665_));
 sky130_fd_sc_hd__o21ai_0 _21212_ (.A1(net463),
    .A2(_10575_),
    .B1(_08558_),
    .Y(_08666_));
 sky130_fd_sc_hd__a21oi_1 _21213_ (.A1(_13080_),
    .A2(_08666_),
    .B1(_08652_),
    .Y(_08667_));
 sky130_fd_sc_hd__a21oi_1 _21214_ (.A1(_08665_),
    .A2(_08667_),
    .B1(_08534_),
    .Y(_00983_));
 sky130_fd_sc_hd__a21oi_2 _21215_ (.A1(_13084_),
    .A2(_08595_),
    .B1(_08525_),
    .Y(_08668_));
 sky130_fd_sc_hd__a22oi_1 _21216_ (.A1(_13086_),
    .A2(_08608_),
    .B1(_08640_),
    .B2(_13080_),
    .Y(_08669_));
 sky130_fd_sc_hd__nand4_1 _21217_ (.A(_08566_),
    .B(_08635_),
    .C(_08668_),
    .D(_08669_),
    .Y(_08670_));
 sky130_fd_sc_hd__a21o_1 _21218_ (.A1(_08549_),
    .A2(_08670_),
    .B1(net525),
    .X(_00984_));
 sky130_fd_sc_hd__a31oi_1 _21219_ (.A1(_13084_),
    .A2(net459),
    .A3(_08551_),
    .B1(_08652_),
    .Y(_08671_));
 sky130_fd_sc_hd__a21oi_1 _21220_ (.A1(_08514_),
    .A2(_08671_),
    .B1(_08534_),
    .Y(_00985_));
 sky130_fd_sc_hd__nor2_1 _21221_ (.A(_10532_),
    .B(_08562_),
    .Y(_08672_));
 sky130_fd_sc_hd__a21oi_1 _21222_ (.A1(_13084_),
    .A2(net507),
    .B1(_13080_),
    .Y(_08673_));
 sky130_fd_sc_hd__nor3_1 _21223_ (.A(_10512_),
    .B(_10564_),
    .C(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand2_1 _21224_ (.A(_13079_),
    .B(_10532_),
    .Y(_08675_));
 sky130_fd_sc_hd__nand2_1 _21225_ (.A(_13080_),
    .B(net507),
    .Y(_08676_));
 sky130_fd_sc_hd__and3_1 _21226_ (.A(_10512_),
    .B(_08675_),
    .C(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__a21oi_1 _21227_ (.A1(_10503_),
    .A2(_08629_),
    .B1(_08677_),
    .Y(_08678_));
 sky130_fd_sc_hd__nor3_1 _21228_ (.A(_08672_),
    .B(_08674_),
    .C(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__a21oi_1 _21229_ (.A1(_08554_),
    .A2(_08679_),
    .B1(_10571_),
    .Y(_08680_));
 sky130_fd_sc_hd__or2_0 _21230_ (.A(net525),
    .B(_08680_),
    .X(_00986_));
 sky130_fd_sc_hd__nor2_1 _21231_ (.A(_08515_),
    .B(_08497_),
    .Y(_08681_));
 sky130_fd_sc_hd__nand2_1 _21232_ (.A(_13079_),
    .B(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__o21ai_0 _21233_ (.A1(_08507_),
    .A2(_08498_),
    .B1(_08682_),
    .Y(_08683_));
 sky130_fd_sc_hd__a2111oi_1 _21234_ (.A1(net507),
    .A2(_08683_),
    .B1(_08572_),
    .C1(_08570_),
    .D1(_08513_),
    .Y(_08684_));
 sky130_fd_sc_hd__a21oi_1 _21235_ (.A1(_13079_),
    .A2(_08505_),
    .B1(_08525_),
    .Y(_08685_));
 sky130_fd_sc_hd__a21oi_1 _21236_ (.A1(_08684_),
    .A2(_08685_),
    .B1(_08534_),
    .Y(_00987_));
 sky130_fd_sc_hd__a21oi_1 _21237_ (.A1(net463),
    .A2(_08659_),
    .B1(_08625_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand2_1 _21238_ (.A(_13080_),
    .B(_08681_),
    .Y(_08687_));
 sky130_fd_sc_hd__o21ai_0 _21239_ (.A1(net459),
    .A2(_08657_),
    .B1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__nand2_1 _21240_ (.A(net507),
    .B(_08688_),
    .Y(_08689_));
 sky130_fd_sc_hd__a31oi_2 _21241_ (.A1(_08524_),
    .A2(_08686_),
    .A3(_08689_),
    .B1(_08534_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _21242_ (.A(net461),
    .B(_08518_),
    .Y(_08690_));
 sky130_fd_sc_hd__a21oi_1 _21243_ (.A1(_13086_),
    .A2(_10512_),
    .B1(_13084_),
    .Y(_08691_));
 sky130_fd_sc_hd__o21ai_0 _21244_ (.A1(net461),
    .A2(_08691_),
    .B1(_08500_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand3_1 _21245_ (.A(_10575_),
    .B(_08690_),
    .C(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__a21oi_2 _21246_ (.A1(_08531_),
    .A2(_08693_),
    .B1(_08534_),
    .Y(_00989_));
 sky130_fd_sc_hd__a21oi_1 _21247_ (.A1(_08585_),
    .A2(_08637_),
    .B1(net459),
    .Y(_08694_));
 sky130_fd_sc_hd__nor2_1 _21248_ (.A(_08513_),
    .B(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__o21ai_0 _21249_ (.A1(_08503_),
    .A2(_08595_),
    .B1(_13084_),
    .Y(_08696_));
 sky130_fd_sc_hd__a21oi_1 _21250_ (.A1(_08508_),
    .A2(_08551_),
    .B1(_08609_),
    .Y(_08697_));
 sky130_fd_sc_hd__a31oi_1 _21251_ (.A1(_08695_),
    .A2(_08696_),
    .A3(_08697_),
    .B1(_08534_),
    .Y(_00990_));
 sky130_fd_sc_hd__nor3b_1 _21252_ (.A(_08674_),
    .B(_08510_),
    .C_N(_08524_),
    .Y(_08698_));
 sky130_fd_sc_hd__a21oi_1 _21253_ (.A1(_08684_),
    .A2(_08698_),
    .B1(_08534_),
    .Y(_00991_));
 sky130_fd_sc_hd__o22ai_1 _21254_ (.A1(_13084_),
    .A2(_10512_),
    .B1(net507),
    .B2(_13086_),
    .Y(_08699_));
 sky130_fd_sc_hd__o211ai_1 _21255_ (.A1(_13086_),
    .A2(_10503_),
    .B1(net507),
    .C1(_10564_),
    .Y(_08700_));
 sky130_fd_sc_hd__o211ai_1 _21256_ (.A1(_13084_),
    .A2(_10532_),
    .B1(net463),
    .C1(_10512_),
    .Y(_08701_));
 sky130_fd_sc_hd__a22oi_1 _21257_ (.A1(_08500_),
    .A2(_08699_),
    .B1(_08700_),
    .B2(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__nor3_1 _21258_ (.A(_08555_),
    .B(_08638_),
    .C(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__o21bai_1 _21259_ (.A1(_10571_),
    .A2(_08703_),
    .B1_N(net525),
    .Y(_00992_));
 sky130_fd_sc_hd__nand2_1 _21260_ (.A(_13079_),
    .B(_08559_),
    .Y(_08704_));
 sky130_fd_sc_hd__o21ai_0 _21261_ (.A1(_13080_),
    .A2(_08641_),
    .B1(_10503_),
    .Y(_08705_));
 sky130_fd_sc_hd__a21oi_1 _21262_ (.A1(_08704_),
    .A2(_08705_),
    .B1(net459),
    .Y(_08706_));
 sky130_fd_sc_hd__o221ai_1 _21263_ (.A1(_08494_),
    .A2(_08556_),
    .B1(_08493_),
    .B2(_08637_),
    .C1(_08594_),
    .Y(_08707_));
 sky130_fd_sc_hd__nor3_1 _21264_ (.A(_08650_),
    .B(_08706_),
    .C(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__nor2_1 _21265_ (.A(_08534_),
    .B(_08708_),
    .Y(_00993_));
 sky130_fd_sc_hd__nor2_1 _21266_ (.A(_13079_),
    .B(_13086_),
    .Y(_08709_));
 sky130_fd_sc_hd__nor2_1 _21267_ (.A(net458),
    .B(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__a21oi_1 _21268_ (.A1(_13084_),
    .A2(net458),
    .B1(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_1 _21269_ (.A(_10532_),
    .B(_08516_),
    .Y(_08712_));
 sky130_fd_sc_hd__nand2_1 _21270_ (.A(net507),
    .B(_08486_),
    .Y(_08713_));
 sky130_fd_sc_hd__a31oi_4 _21271_ (.A1(_08626_),
    .A2(_08712_),
    .A3(_08713_),
    .B1(_08485_),
    .Y(_08714_));
 sky130_fd_sc_hd__o2111ai_1 _21272_ (.A1(_08487_),
    .A2(_08711_),
    .B1(_08714_),
    .C1(_08584_),
    .D1(_08506_),
    .Y(_08715_));
 sky130_fd_sc_hd__a21o_1 _21273_ (.A1(_08549_),
    .A2(_08715_),
    .B1(net525),
    .X(_00994_));
 sky130_fd_sc_hd__nand2_1 _21274_ (.A(_13080_),
    .B(_10512_),
    .Y(_08716_));
 sky130_fd_sc_hd__o21ai_0 _21275_ (.A1(_10512_),
    .A2(_08709_),
    .B1(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__a22oi_1 _21276_ (.A1(_13084_),
    .A2(_08498_),
    .B1(_08717_),
    .B2(net463),
    .Y(_08718_));
 sky130_fd_sc_hd__a21oi_1 _21277_ (.A1(net507),
    .A2(_08484_),
    .B1(net463),
    .Y(_08719_));
 sky130_fd_sc_hd__nand2_1 _21278_ (.A(_08486_),
    .B(_08608_),
    .Y(_08720_));
 sky130_fd_sc_hd__o2111ai_1 _21279_ (.A1(_13080_),
    .A2(_08719_),
    .B1(_08720_),
    .C1(_10512_),
    .D1(_08542_),
    .Y(_08721_));
 sky130_fd_sc_hd__o21ai_0 _21280_ (.A1(_10532_),
    .A2(_08718_),
    .B1(_08721_),
    .Y(_08722_));
 sky130_fd_sc_hd__a2111oi_1 _21281_ (.A1(net463),
    .A2(_08659_),
    .B1(_08722_),
    .C1(_08532_),
    .D1(_08638_),
    .Y(_08723_));
 sky130_fd_sc_hd__o21bai_1 _21282_ (.A1(_10571_),
    .A2(_08723_),
    .B1_N(net525),
    .Y(_00995_));
 sky130_fd_sc_hd__o21ai_0 _21283_ (.A1(_08626_),
    .A2(_08595_),
    .B1(_13084_),
    .Y(_08724_));
 sky130_fd_sc_hd__o21ai_0 _21284_ (.A1(_08507_),
    .A2(_08498_),
    .B1(_08637_),
    .Y(_08725_));
 sky130_fd_sc_hd__nor2_1 _21285_ (.A(net459),
    .B(_08539_),
    .Y(_08726_));
 sky130_fd_sc_hd__a221oi_1 _21286_ (.A1(_08497_),
    .A2(_08641_),
    .B1(_08725_),
    .B2(net503),
    .C1(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__a31oi_1 _21287_ (.A1(_08506_),
    .A2(_08724_),
    .A3(_08727_),
    .B1(_08534_),
    .Y(_00996_));
 sky130_fd_sc_hd__nand3_1 _21288_ (.A(_08585_),
    .B(_08588_),
    .C(_08637_),
    .Y(_08728_));
 sky130_fd_sc_hd__o21ai_0 _21289_ (.A1(_08690_),
    .A2(_08709_),
    .B1(_08714_),
    .Y(_08729_));
 sky130_fd_sc_hd__a21oi_1 _21290_ (.A1(net459),
    .A2(_08728_),
    .B1(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__a21oi_1 _21291_ (.A1(_08668_),
    .A2(_08730_),
    .B1(_08534_),
    .Y(_00997_));
 sky130_fd_sc_hd__nor3_1 _21292_ (.A(_13079_),
    .B(_13080_),
    .C(_13086_),
    .Y(_08731_));
 sky130_fd_sc_hd__o21bai_1 _21293_ (.A1(_08556_),
    .A2(_08731_),
    .B1_N(_08532_),
    .Y(_08732_));
 sky130_fd_sc_hd__a22oi_1 _21294_ (.A1(net495),
    .A2(_08508_),
    .B1(_08515_),
    .B2(_13084_),
    .Y(_08733_));
 sky130_fd_sc_hd__o21ai_0 _21295_ (.A1(_13079_),
    .A2(_08495_),
    .B1(_08505_),
    .Y(_08734_));
 sky130_fd_sc_hd__o21ai_0 _21296_ (.A1(net490),
    .A2(_08733_),
    .B1(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__nor4_1 _21297_ (.A(_08655_),
    .B(_08706_),
    .C(_08732_),
    .D(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__o21bai_1 _21298_ (.A1(_10571_),
    .A2(_08736_),
    .B1_N(net525),
    .Y(_00998_));
 sky130_fd_sc_hd__o21ai_0 _21299_ (.A1(_13086_),
    .A2(_08519_),
    .B1(_08515_),
    .Y(_08737_));
 sky130_fd_sc_hd__a21oi_1 _21300_ (.A1(_08618_),
    .A2(_08737_),
    .B1(_10532_),
    .Y(_08738_));
 sky130_fd_sc_hd__a21oi_1 _21301_ (.A1(_08563_),
    .A2(_08569_),
    .B1(_10512_),
    .Y(_08739_));
 sky130_fd_sc_hd__nand2_1 _21302_ (.A(_10564_),
    .B(_08586_),
    .Y(_08740_));
 sky130_fd_sc_hd__nand2_1 _21303_ (.A(_08663_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__nor4_1 _21304_ (.A(_08732_),
    .B(_08738_),
    .C(_08739_),
    .D(_08741_),
    .Y(_08742_));
 sky130_fd_sc_hd__o21bai_1 _21305_ (.A1(_10571_),
    .A2(_08742_),
    .B1_N(net525),
    .Y(_00999_));
 sky130_fd_sc_hd__a22oi_1 _21306_ (.A1(_13084_),
    .A2(_08518_),
    .B1(_08559_),
    .B2(_13080_),
    .Y(_08743_));
 sky130_fd_sc_hd__o2111ai_1 _21307_ (.A1(net458),
    .A2(_08743_),
    .B1(_08714_),
    .C1(_08689_),
    .D1(_08621_),
    .Y(_08744_));
 sky130_fd_sc_hd__a21o_1 _21308_ (.A1(_08549_),
    .A2(_08744_),
    .B1(net525),
    .X(_01000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_946 ();
 sky130_fd_sc_hd__xnor2_4 _21311_ (.A(\count_hash2[4] ),
    .B(_10015_),
    .Y(_08747_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_945 ();
 sky130_fd_sc_hd__nand2_4 _21313_ (.A(_08747_),
    .B(net518),
    .Y(_08749_));
 sky130_fd_sc_hd__xnor2_4 _21314_ (.A(\count_hash2[3] ),
    .B(_13076_),
    .Y(_08750_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_944 ();
 sky130_fd_sc_hd__xor2_4 _21316_ (.A(\count_hash2[5] ),
    .B(_10026_),
    .X(_08752_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_943 ();
 sky130_fd_sc_hd__nor2_2 _21318_ (.A(_08747_),
    .B(_08752_),
    .Y(_08754_));
 sky130_fd_sc_hd__nand2_1 _21319_ (.A(_08750_),
    .B(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__nand2_1 _21320_ (.A(_08749_),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__nand2_1 _21321_ (.A(_13072_),
    .B(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_941 ();
 sky130_fd_sc_hd__or3_4 _21324_ (.A(_13069_),
    .B(_13072_),
    .C(_13074_),
    .X(_08760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_940 ();
 sky130_fd_sc_hd__nor2_4 _21326_ (.A(_13070_),
    .B(_08760_),
    .Y(_08762_));
 sky130_fd_sc_hd__nand2_1 _21327_ (.A(_10016_),
    .B(_08750_),
    .Y(_08763_));
 sky130_fd_sc_hd__or2_4 _21328_ (.A(_13069_),
    .B(_13070_),
    .X(_08764_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_939 ();
 sky130_fd_sc_hd__nor2_1 _21330_ (.A(_13074_),
    .B(_08764_),
    .Y(_08766_));
 sky130_fd_sc_hd__o22ai_1 _21331_ (.A1(_08762_),
    .A2(_08763_),
    .B1(_08766_),
    .B2(_08749_),
    .Y(_08767_));
 sky130_fd_sc_hd__nor2_2 _21332_ (.A(net518),
    .B(_08752_),
    .Y(_08768_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_938 ();
 sky130_fd_sc_hd__nand2_2 _21334_ (.A(_13069_),
    .B(_10016_),
    .Y(_08770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_937 ();
 sky130_fd_sc_hd__nand2_2 _21336_ (.A(_08747_),
    .B(_08752_),
    .Y(_08772_));
 sky130_fd_sc_hd__nand2_1 _21337_ (.A(_13074_),
    .B(_08772_),
    .Y(_08773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_936 ();
 sky130_fd_sc_hd__a21oi_1 _21339_ (.A1(_08770_),
    .A2(_08773_),
    .B1(_08750_),
    .Y(_08775_));
 sky130_fd_sc_hd__a221oi_1 _21340_ (.A1(_08752_),
    .A2(_08767_),
    .B1(_08768_),
    .B2(_08764_),
    .C1(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_935 ();
 sky130_fd_sc_hd__o21ai_4 _21342_ (.A1(_13070_),
    .A2(_08760_),
    .B1(_10573_),
    .Y(_08778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_934 ();
 sky130_fd_sc_hd__a21oi_1 _21344_ (.A1(_08757_),
    .A2(_08776_),
    .B1(_08778_),
    .Y(_08780_));
 sky130_fd_sc_hd__or2_0 _21345_ (.A(net525),
    .B(_08780_),
    .X(_01001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_933 ();
 sky130_fd_sc_hd__nor2_1 _21347_ (.A(_08750_),
    .B(_10027_),
    .Y(_08782_));
 sky130_fd_sc_hd__nor2_1 _21348_ (.A(_08768_),
    .B(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_932 ();
 sky130_fd_sc_hd__a221oi_1 _21350_ (.A1(_13069_),
    .A2(_08768_),
    .B1(_08783_),
    .B2(_13072_),
    .C1(_10016_),
    .Y(_08785_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_931 ();
 sky130_fd_sc_hd__nor2_1 _21352_ (.A(_13072_),
    .B(_13074_),
    .Y(_08787_));
 sky130_fd_sc_hd__nand2_1 _21353_ (.A(_13069_),
    .B(_08750_),
    .Y(_08788_));
 sky130_fd_sc_hd__o21ai_1 _21354_ (.A1(_08750_),
    .A2(_08787_),
    .B1(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_930 ();
 sky130_fd_sc_hd__a221oi_1 _21356_ (.A1(_13070_),
    .A2(_08750_),
    .B1(_10027_),
    .B2(_08789_),
    .C1(_08747_),
    .Y(_08791_));
 sky130_fd_sc_hd__clkinv_2 _21357_ (.A(_13069_),
    .Y(_08792_));
 sky130_fd_sc_hd__nand2_2 _21358_ (.A(net518),
    .B(_08752_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand2_1 _21359_ (.A(_13070_),
    .B(_08768_),
    .Y(_08794_));
 sky130_fd_sc_hd__o21ai_0 _21360_ (.A1(_08792_),
    .A2(_08793_),
    .B1(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__o21ai_0 _21361_ (.A1(net518),
    .A2(_08754_),
    .B1(_08772_),
    .Y(_08796_));
 sky130_fd_sc_hd__a22o_1 _21362_ (.A1(_08747_),
    .A2(_08795_),
    .B1(_08796_),
    .B2(_13074_),
    .X(_08797_));
 sky130_fd_sc_hd__o22ai_4 _21363_ (.A1(_13070_),
    .A2(_08760_),
    .B1(_08770_),
    .B2(_08793_),
    .Y(_08798_));
 sky130_fd_sc_hd__nor2_1 _21364_ (.A(_08797_),
    .B(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__o21ai_0 _21365_ (.A1(_08785_),
    .A2(_08791_),
    .B1(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__a21o_1 _21366_ (.A1(_08549_),
    .A2(_08800_),
    .B1(net525),
    .X(_01002_));
 sky130_fd_sc_hd__a21oi_1 _21367_ (.A1(_13074_),
    .A2(_10016_),
    .B1(_13069_),
    .Y(_08801_));
 sky130_fd_sc_hd__nand2_1 _21368_ (.A(_13070_),
    .B(_08747_),
    .Y(_08802_));
 sky130_fd_sc_hd__o21ai_0 _21369_ (.A1(_08750_),
    .A2(_08801_),
    .B1(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__nor2_2 _21370_ (.A(_13072_),
    .B(_08764_),
    .Y(_08804_));
 sky130_fd_sc_hd__nor3_1 _21371_ (.A(_08752_),
    .B(_08763_),
    .C(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__a21oi_1 _21372_ (.A1(_08752_),
    .A2(_08803_),
    .B1(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_929 ();
 sky130_fd_sc_hd__nor2_1 _21374_ (.A(_08747_),
    .B(net518),
    .Y(_08808_));
 sky130_fd_sc_hd__a31oi_1 _21375_ (.A1(_08752_),
    .A2(_08808_),
    .A3(_08764_),
    .B1(_08762_),
    .Y(_08809_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_928 ();
 sky130_fd_sc_hd__or2_2 _21377_ (.A(_13070_),
    .B(_13072_),
    .X(_08811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_927 ();
 sky130_fd_sc_hd__nor2_2 _21379_ (.A(net512),
    .B(_08752_),
    .Y(_08813_));
 sky130_fd_sc_hd__o21ai_0 _21380_ (.A1(_08750_),
    .A2(_08811_),
    .B1(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__a31oi_1 _21381_ (.A1(_08806_),
    .A2(_08809_),
    .A3(_08814_),
    .B1(net454),
    .Y(_01003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_925 ();
 sky130_fd_sc_hd__nand2_1 _21384_ (.A(_08750_),
    .B(net466),
    .Y(_08817_));
 sky130_fd_sc_hd__nand2_1 _21385_ (.A(_08817_),
    .B(_08793_),
    .Y(_08818_));
 sky130_fd_sc_hd__nor2_1 _21386_ (.A(_10016_),
    .B(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__nor2_1 _21387_ (.A(_08747_),
    .B(_08783_),
    .Y(_08820_));
 sky130_fd_sc_hd__nor2_1 _21388_ (.A(_08819_),
    .B(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__nor2_4 _21389_ (.A(_08747_),
    .B(_08750_),
    .Y(_08822_));
 sky130_fd_sc_hd__nor2_1 _21390_ (.A(net512),
    .B(net518),
    .Y(_08823_));
 sky130_fd_sc_hd__nor2_2 _21391_ (.A(_08822_),
    .B(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__a22oi_1 _21392_ (.A1(_08760_),
    .A2(_08822_),
    .B1(_08824_),
    .B2(_13072_),
    .Y(_08825_));
 sky130_fd_sc_hd__nor2_2 _21393_ (.A(_08747_),
    .B(net466),
    .Y(_08826_));
 sky130_fd_sc_hd__nand2_4 _21394_ (.A(_08747_),
    .B(_10027_),
    .Y(_08827_));
 sky130_fd_sc_hd__nor2_2 _21395_ (.A(_08750_),
    .B(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_924 ();
 sky130_fd_sc_hd__o21ai_0 _21397_ (.A1(_08826_),
    .A2(_08828_),
    .B1(_13070_),
    .Y(_08830_));
 sky130_fd_sc_hd__o21ai_0 _21398_ (.A1(_10027_),
    .A2(_08825_),
    .B1(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__a21oi_1 _21399_ (.A1(_13069_),
    .A2(_08821_),
    .B1(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__nor2_1 _21400_ (.A(_08778_),
    .B(_08832_),
    .Y(_01004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_923 ();
 sky130_fd_sc_hd__inv_2 _21402_ (.A(_13072_),
    .Y(_08834_));
 sky130_fd_sc_hd__nand2_2 _21403_ (.A(_08792_),
    .B(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__nand2_1 _21404_ (.A(_08747_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__nor2_1 _21405_ (.A(_13070_),
    .B(_13074_),
    .Y(_08837_));
 sky130_fd_sc_hd__nor2_1 _21406_ (.A(net512),
    .B(_08750_),
    .Y(_08838_));
 sky130_fd_sc_hd__a211o_1 _21407_ (.A1(_08836_),
    .A2(_08837_),
    .B1(_08752_),
    .C1(_08838_),
    .X(_08839_));
 sky130_fd_sc_hd__nor2_1 _21408_ (.A(_13070_),
    .B(_13072_),
    .Y(_08840_));
 sky130_fd_sc_hd__nand2_1 _21409_ (.A(_10016_),
    .B(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__nor2_1 _21410_ (.A(_13069_),
    .B(_13070_),
    .Y(_08842_));
 sky130_fd_sc_hd__nand2_1 _21411_ (.A(_08747_),
    .B(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__a31oi_2 _21412_ (.A1(_08782_),
    .A2(_08841_),
    .A3(_08843_),
    .B1(_08798_),
    .Y(_08844_));
 sky130_fd_sc_hd__nand2_4 _21413_ (.A(_08750_),
    .B(_08752_),
    .Y(_08845_));
 sky130_fd_sc_hd__nor2_2 _21414_ (.A(_08750_),
    .B(_08752_),
    .Y(_08846_));
 sky130_fd_sc_hd__o21ai_1 _21415_ (.A1(_13074_),
    .A2(_08811_),
    .B1(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__o21ai_0 _21416_ (.A1(_08792_),
    .A2(_08845_),
    .B1(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nand2_1 _21417_ (.A(_08747_),
    .B(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__a31oi_1 _21418_ (.A1(_08839_),
    .A2(_08844_),
    .A3(_08849_),
    .B1(net454),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _21419_ (.A(_13070_),
    .B(_08752_),
    .Y(_08850_));
 sky130_fd_sc_hd__nand2_2 _21420_ (.A(_13074_),
    .B(net518),
    .Y(_08851_));
 sky130_fd_sc_hd__nand3_1 _21421_ (.A(_10016_),
    .B(_08850_),
    .C(_08851_),
    .Y(_08852_));
 sky130_fd_sc_hd__a21oi_1 _21422_ (.A1(_13069_),
    .A2(_08817_),
    .B1(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__a21oi_1 _21423_ (.A1(_08747_),
    .A2(_08847_),
    .B1(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__nor2_4 _21424_ (.A(net454),
    .B(_08762_),
    .Y(_08855_));
 sky130_fd_sc_hd__o21ai_2 _21425_ (.A1(_08797_),
    .A2(_08854_),
    .B1(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__nand2b_1 _21426_ (.A_N(net525),
    .B(_08856_),
    .Y(_01006_));
 sky130_fd_sc_hd__nor2_2 _21427_ (.A(net512),
    .B(net466),
    .Y(_08857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_922 ();
 sky130_fd_sc_hd__o21ai_0 _21429_ (.A1(net518),
    .A2(_08804_),
    .B1(_08851_),
    .Y(_08859_));
 sky130_fd_sc_hd__nand2_1 _21430_ (.A(_13072_),
    .B(_08752_),
    .Y(_08860_));
 sky130_fd_sc_hd__nand2_1 _21431_ (.A(_13070_),
    .B(net511),
    .Y(_08861_));
 sky130_fd_sc_hd__nor2_4 _21432_ (.A(_08857_),
    .B(_08754_),
    .Y(_08862_));
 sky130_fd_sc_hd__a221oi_1 _21433_ (.A1(_13072_),
    .A2(_08813_),
    .B1(_08862_),
    .B2(_13069_),
    .C1(net518),
    .Y(_08863_));
 sky130_fd_sc_hd__a31oi_1 _21434_ (.A1(net518),
    .A2(_08860_),
    .A3(_08861_),
    .B1(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__a21oi_1 _21435_ (.A1(_08857_),
    .A2(_08859_),
    .B1(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__nor2_1 _21436_ (.A(_08778_),
    .B(_08865_),
    .Y(_01007_));
 sky130_fd_sc_hd__a22oi_1 _21437_ (.A1(_13069_),
    .A2(_08813_),
    .B1(_08862_),
    .B2(_13070_),
    .Y(_08866_));
 sky130_fd_sc_hd__nand2_2 _21438_ (.A(_10016_),
    .B(net518),
    .Y(_08867_));
 sky130_fd_sc_hd__o21bai_1 _21439_ (.A1(_10027_),
    .A2(_08804_),
    .B1_N(_13074_),
    .Y(_08868_));
 sky130_fd_sc_hd__nor2_1 _21440_ (.A(_13074_),
    .B(_08835_),
    .Y(_08869_));
 sky130_fd_sc_hd__o21ai_0 _21441_ (.A1(_08869_),
    .A2(_08857_),
    .B1(_08750_),
    .Y(_08870_));
 sky130_fd_sc_hd__nand2_1 _21442_ (.A(_13072_),
    .B(net466),
    .Y(_08871_));
 sky130_fd_sc_hd__a21boi_1 _21443_ (.A1(_13074_),
    .A2(_08752_),
    .B1_N(_08871_),
    .Y(_08872_));
 sky130_fd_sc_hd__o22ai_4 _21444_ (.A1(_08845_),
    .A2(_08802_),
    .B1(_08867_),
    .B2(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__a31oi_1 _21445_ (.A1(_08867_),
    .A2(_08868_),
    .A3(_08870_),
    .B1(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__o21ai_1 _21446_ (.A1(_08750_),
    .A2(_08866_),
    .B1(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__a21o_1 _21447_ (.A1(_08855_),
    .A2(_08875_),
    .B1(net525),
    .X(_01008_));
 sky130_fd_sc_hd__nand2_1 _21448_ (.A(_08755_),
    .B(_08793_),
    .Y(_08876_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_921 ();
 sky130_fd_sc_hd__o21ai_0 _21450_ (.A1(_13074_),
    .A2(_08845_),
    .B1(_08749_),
    .Y(_08878_));
 sky130_fd_sc_hd__a22o_1 _21451_ (.A1(_13074_),
    .A2(_08838_),
    .B1(_08837_),
    .B2(_08835_),
    .X(_08879_));
 sky130_fd_sc_hd__a21oi_1 _21452_ (.A1(_13070_),
    .A2(_08878_),
    .B1(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__a221oi_1 _21453_ (.A1(_13069_),
    .A2(_08828_),
    .B1(_08876_),
    .B2(_13072_),
    .C1(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__o21bai_2 _21454_ (.A1(_10571_),
    .A2(_08881_),
    .B1_N(net525),
    .Y(_01009_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_920 ();
 sky130_fd_sc_hd__o21ai_0 _21456_ (.A1(_08747_),
    .A2(_08845_),
    .B1(_08827_),
    .Y(_08883_));
 sky130_fd_sc_hd__a21oi_1 _21457_ (.A1(_13074_),
    .A2(_08747_),
    .B1(_13069_),
    .Y(_08884_));
 sky130_fd_sc_hd__a21oi_1 _21458_ (.A1(_08861_),
    .A2(_08884_),
    .B1(_08845_),
    .Y(_08885_));
 sky130_fd_sc_hd__o21ai_0 _21459_ (.A1(_13070_),
    .A2(_08752_),
    .B1(_08747_),
    .Y(_08886_));
 sky130_fd_sc_hd__a32o_1 _21460_ (.A1(_08792_),
    .A2(net518),
    .A3(_08860_),
    .B1(_08857_),
    .B2(_08834_),
    .X(_08887_));
 sky130_fd_sc_hd__a21oi_1 _21461_ (.A1(_08750_),
    .A2(_08886_),
    .B1(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__a211oi_1 _21462_ (.A1(_13074_),
    .A2(_08883_),
    .B1(_08885_),
    .C1(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__o21bai_1 _21463_ (.A1(_08778_),
    .A2(_08889_),
    .B1_N(net525),
    .Y(_01010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_919 ();
 sky130_fd_sc_hd__nand2_1 _21465_ (.A(_08834_),
    .B(net511),
    .Y(_08891_));
 sky130_fd_sc_hd__a21oi_1 _21466_ (.A1(_08843_),
    .A2(_08891_),
    .B1(_13074_),
    .Y(_08892_));
 sky130_fd_sc_hd__nor3_1 _21467_ (.A(net517),
    .B(_08862_),
    .C(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__a31oi_1 _21468_ (.A1(net466),
    .A2(_08835_),
    .A3(_08822_),
    .B1(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__a21oi_1 _21469_ (.A1(_08750_),
    .A2(_08811_),
    .B1(_10016_),
    .Y(_08895_));
 sky130_fd_sc_hd__a311oi_1 _21470_ (.A1(_10016_),
    .A2(_08788_),
    .A3(_08851_),
    .B1(_08895_),
    .C1(_08752_),
    .Y(_08896_));
 sky130_fd_sc_hd__a31oi_2 _21471_ (.A1(_13070_),
    .A2(_10016_),
    .A3(_08783_),
    .B1(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__a31oi_1 _21472_ (.A1(_08844_),
    .A2(_08894_),
    .A3(_08897_),
    .B1(net454),
    .Y(_01011_));
 sky130_fd_sc_hd__nor2_1 _21473_ (.A(_10016_),
    .B(_08845_),
    .Y(_08898_));
 sky130_fd_sc_hd__o21ai_0 _21474_ (.A1(_08846_),
    .A2(_08898_),
    .B1(_13074_),
    .Y(_08899_));
 sky130_fd_sc_hd__nand3_1 _21475_ (.A(_13069_),
    .B(_08845_),
    .C(_08827_),
    .Y(_08900_));
 sky130_fd_sc_hd__a22oi_1 _21476_ (.A1(_13072_),
    .A2(_08818_),
    .B1(_08811_),
    .B2(_08747_),
    .Y(_08901_));
 sky130_fd_sc_hd__a31oi_2 _21477_ (.A1(_08899_),
    .A2(_08900_),
    .A3(_08901_),
    .B1(_08778_),
    .Y(_01012_));
 sky130_fd_sc_hd__a21oi_1 _21478_ (.A1(_08749_),
    .A2(_08811_),
    .B1(_13069_),
    .Y(_08902_));
 sky130_fd_sc_hd__a21oi_1 _21479_ (.A1(_08840_),
    .A2(_08823_),
    .B1(_08902_),
    .Y(_08903_));
 sky130_fd_sc_hd__o22ai_1 _21480_ (.A1(_08811_),
    .A2(_08867_),
    .B1(_08903_),
    .B2(_13074_),
    .Y(_08904_));
 sky130_fd_sc_hd__nand2_1 _21481_ (.A(_13072_),
    .B(_08747_),
    .Y(_08905_));
 sky130_fd_sc_hd__nor2_1 _21482_ (.A(_13069_),
    .B(net518),
    .Y(_08906_));
 sky130_fd_sc_hd__a32oi_1 _21483_ (.A1(_08861_),
    .A2(_08905_),
    .A3(_08906_),
    .B1(_08822_),
    .B2(_08834_),
    .Y(_08907_));
 sky130_fd_sc_hd__o221ai_1 _21484_ (.A1(_08749_),
    .A2(_08811_),
    .B1(_08907_),
    .B2(_13074_),
    .C1(net466),
    .Y(_08908_));
 sky130_fd_sc_hd__o21ai_1 _21485_ (.A1(net466),
    .A2(_08904_),
    .B1(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__a21o_1 _21486_ (.A1(_08855_),
    .A2(_08909_),
    .B1(net525),
    .X(_01013_));
 sky130_fd_sc_hd__nand2_1 _21487_ (.A(_08770_),
    .B(_08802_),
    .Y(_08910_));
 sky130_fd_sc_hd__o21ai_0 _21488_ (.A1(_13074_),
    .A2(_08910_),
    .B1(_08750_),
    .Y(_08911_));
 sky130_fd_sc_hd__a21oi_1 _21489_ (.A1(_08834_),
    .A2(_08911_),
    .B1(_08822_),
    .Y(_08912_));
 sky130_fd_sc_hd__o2bb2ai_1 _21490_ (.A1_N(_08754_),
    .A2_N(_08804_),
    .B1(_08912_),
    .B2(net466),
    .Y(_08913_));
 sky130_fd_sc_hd__nand2_1 _21491_ (.A(_08750_),
    .B(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__nor2_1 _21492_ (.A(_13074_),
    .B(net512),
    .Y(_08915_));
 sky130_fd_sc_hd__o21ai_0 _21493_ (.A1(_08822_),
    .A2(_08915_),
    .B1(_08792_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand2_1 _21494_ (.A(net518),
    .B(_08915_),
    .Y(_08917_));
 sky130_fd_sc_hd__a21oi_1 _21495_ (.A1(_08916_),
    .A2(_08917_),
    .B1(_13070_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand2_1 _21496_ (.A(_08752_),
    .B(_08912_),
    .Y(_08919_));
 sky130_fd_sc_hd__o21ai_0 _21497_ (.A1(_08826_),
    .A2(_08918_),
    .B1(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__a31o_1 _21498_ (.A1(_08855_),
    .A2(_08914_),
    .A3(_08920_),
    .B1(net525),
    .X(_01014_));
 sky130_fd_sc_hd__a21oi_1 _21499_ (.A1(_13069_),
    .A2(net518),
    .B1(_13072_),
    .Y(_08921_));
 sky130_fd_sc_hd__o21ai_1 _21500_ (.A1(net518),
    .A2(_08827_),
    .B1(_13070_),
    .Y(_08922_));
 sky130_fd_sc_hd__nor2_1 _21501_ (.A(_13072_),
    .B(_10027_),
    .Y(_08923_));
 sky130_fd_sc_hd__nor3_1 _21502_ (.A(_08750_),
    .B(_08752_),
    .C(_08764_),
    .Y(_08924_));
 sky130_fd_sc_hd__o21ai_1 _21503_ (.A1(_08923_),
    .A2(_08924_),
    .B1(_10016_),
    .Y(_08925_));
 sky130_fd_sc_hd__o311ai_4 _21504_ (.A1(_13069_),
    .A2(_08750_),
    .A3(_08772_),
    .B1(_08925_),
    .C1(_08855_),
    .Y(_08926_));
 sky130_fd_sc_hd__a21oi_4 _21505_ (.A1(_08921_),
    .A2(_08922_),
    .B1(_08926_),
    .Y(_01015_));
 sky130_fd_sc_hd__a21oi_1 _21506_ (.A1(_13070_),
    .A2(net512),
    .B1(_13072_),
    .Y(_08927_));
 sky130_fd_sc_hd__nand2_1 _21507_ (.A(_13074_),
    .B(_08823_),
    .Y(_08928_));
 sky130_fd_sc_hd__o21ai_2 _21508_ (.A1(_08750_),
    .A2(_08927_),
    .B1(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__nand3_1 _21509_ (.A(_08750_),
    .B(_08835_),
    .C(_08862_),
    .Y(_08930_));
 sky130_fd_sc_hd__or2_0 _21510_ (.A(_13069_),
    .B(_13074_),
    .X(_08931_));
 sky130_fd_sc_hd__a21oi_2 _21511_ (.A1(_08828_),
    .A2(_08931_),
    .B1(_08762_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand2_1 _21512_ (.A(_08930_),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__a211oi_4 _21513_ (.A1(_08752_),
    .A2(_08929_),
    .B1(_08933_),
    .C1(_08873_),
    .Y(_08934_));
 sky130_fd_sc_hd__nor2_1 _21514_ (.A(net454),
    .B(_08934_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _21515_ (.A(_13072_),
    .B(net518),
    .Y(_08935_));
 sky130_fd_sc_hd__nand2_1 _21516_ (.A(_13074_),
    .B(_08750_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand3_1 _21517_ (.A(_08747_),
    .B(_08935_),
    .C(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__nand2_1 _21518_ (.A(_08752_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__a21oi_1 _21519_ (.A1(_08760_),
    .A2(_08867_),
    .B1(_13070_),
    .Y(_08939_));
 sky130_fd_sc_hd__o21ai_1 _21520_ (.A1(_08938_),
    .A2(_08939_),
    .B1(_08900_),
    .Y(_08940_));
 sky130_fd_sc_hd__a21o_1 _21521_ (.A1(_08855_),
    .A2(_08940_),
    .B1(net525),
    .X(_01017_));
 sky130_fd_sc_hd__nand2_1 _21522_ (.A(_13070_),
    .B(_08813_),
    .Y(_08941_));
 sky130_fd_sc_hd__o21ai_0 _21523_ (.A1(_08792_),
    .A2(_08862_),
    .B1(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__a21oi_2 _21524_ (.A1(net518),
    .A2(_08942_),
    .B1(_08762_),
    .Y(_08943_));
 sky130_fd_sc_hd__nor2_1 _21525_ (.A(_08766_),
    .B(_08846_),
    .Y(_08944_));
 sky130_fd_sc_hd__a21oi_1 _21526_ (.A1(_08752_),
    .A2(_08851_),
    .B1(_08747_),
    .Y(_08945_));
 sky130_fd_sc_hd__o21ai_1 _21527_ (.A1(_13072_),
    .A2(_08944_),
    .B1(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__o21ai_0 _21528_ (.A1(_10016_),
    .A2(_08787_),
    .B1(_08850_),
    .Y(_08947_));
 sky130_fd_sc_hd__nand2_1 _21529_ (.A(_08750_),
    .B(_08947_),
    .Y(_08948_));
 sky130_fd_sc_hd__a31oi_4 _21530_ (.A1(_08943_),
    .A2(_08946_),
    .A3(_08948_),
    .B1(_10035_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand3_1 _21531_ (.A(_08750_),
    .B(_10027_),
    .C(_08760_),
    .Y(_08949_));
 sky130_fd_sc_hd__o21ai_0 _21532_ (.A1(_08750_),
    .A2(_08804_),
    .B1(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__nor2_1 _21533_ (.A(_08770_),
    .B(_08793_),
    .Y(_08951_));
 sky130_fd_sc_hd__a21oi_2 _21534_ (.A1(_08747_),
    .A2(_08950_),
    .B1(_08951_),
    .Y(_08952_));
 sky130_fd_sc_hd__a21oi_1 _21535_ (.A1(_08894_),
    .A2(_08952_),
    .B1(_08778_),
    .Y(_01019_));
 sky130_fd_sc_hd__a21oi_1 _21536_ (.A1(_13069_),
    .A2(net518),
    .B1(_13074_),
    .Y(_08953_));
 sky130_fd_sc_hd__o22ai_1 _21537_ (.A1(_08817_),
    .A2(_08840_),
    .B1(_08953_),
    .B2(net466),
    .Y(_08954_));
 sky130_fd_sc_hd__a21oi_1 _21538_ (.A1(_10016_),
    .A2(_08764_),
    .B1(_13072_),
    .Y(_08955_));
 sky130_fd_sc_hd__a31oi_1 _21539_ (.A1(_13069_),
    .A2(_08747_),
    .A3(net518),
    .B1(_13074_),
    .Y(_08956_));
 sky130_fd_sc_hd__o22ai_1 _21540_ (.A1(_08845_),
    .A2(_08955_),
    .B1(_08956_),
    .B2(_08752_),
    .Y(_08957_));
 sky130_fd_sc_hd__a21oi_1 _21541_ (.A1(_08747_),
    .A2(_08954_),
    .B1(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__nor2_2 _21542_ (.A(_08778_),
    .B(_08958_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_1 _21543_ (.A(_13070_),
    .B(_08846_),
    .Y(_08959_));
 sky130_fd_sc_hd__o21ai_0 _21544_ (.A1(_08845_),
    .A2(_08787_),
    .B1(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__a21oi_1 _21545_ (.A1(_13069_),
    .A2(_08750_),
    .B1(_13074_),
    .Y(_08961_));
 sky130_fd_sc_hd__o22ai_1 _21546_ (.A1(_08862_),
    .A2(_08935_),
    .B1(_08961_),
    .B2(_08827_),
    .Y(_08962_));
 sky130_fd_sc_hd__a21oi_1 _21547_ (.A1(_10016_),
    .A2(_08960_),
    .B1(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__a21oi_1 _21548_ (.A1(_08806_),
    .A2(_08963_),
    .B1(_08778_),
    .Y(_08964_));
 sky130_fd_sc_hd__or2_0 _21549_ (.A(net525),
    .B(_08964_),
    .X(_01021_));
 sky130_fd_sc_hd__a22oi_2 _21550_ (.A1(_08747_),
    .A2(_08764_),
    .B1(_08827_),
    .B2(_13074_),
    .Y(_08965_));
 sky130_fd_sc_hd__a22oi_1 _21551_ (.A1(_13074_),
    .A2(_08838_),
    .B1(_08824_),
    .B2(_13072_),
    .Y(_08966_));
 sky130_fd_sc_hd__nand2_1 _21552_ (.A(net512),
    .B(net466),
    .Y(_08967_));
 sky130_fd_sc_hd__a222oi_1 _21553_ (.A1(_13070_),
    .A2(_08808_),
    .B1(_08838_),
    .B2(_13074_),
    .C1(_08824_),
    .C2(_13069_),
    .Y(_08968_));
 sky130_fd_sc_hd__o22a_1 _21554_ (.A1(_08967_),
    .A2(_08851_),
    .B1(_08968_),
    .B2(net466),
    .X(_08969_));
 sky130_fd_sc_hd__o221ai_2 _21555_ (.A1(net518),
    .A2(_08965_),
    .B1(_08966_),
    .B2(_08752_),
    .C1(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__a21o_2 _21556_ (.A1(_08855_),
    .A2(_08970_),
    .B1(net525),
    .X(_01022_));
 sky130_fd_sc_hd__nand2_1 _21557_ (.A(_13070_),
    .B(_08818_),
    .Y(_08971_));
 sky130_fd_sc_hd__a221oi_1 _21558_ (.A1(_13069_),
    .A2(_08768_),
    .B1(_08868_),
    .B2(net518),
    .C1(_10016_),
    .Y(_08972_));
 sky130_fd_sc_hd__a31oi_1 _21559_ (.A1(_10016_),
    .A2(_08935_),
    .A3(_08971_),
    .B1(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__o21a_1 _21560_ (.A1(_08885_),
    .A2(_08973_),
    .B1(_08855_),
    .X(_01023_));
 sky130_fd_sc_hd__nor2_1 _21561_ (.A(_08752_),
    .B(_08915_),
    .Y(_08974_));
 sky130_fd_sc_hd__nor2_1 _21562_ (.A(_08750_),
    .B(_08857_),
    .Y(_08975_));
 sky130_fd_sc_hd__o221ai_1 _21563_ (.A1(_08835_),
    .A2(_08967_),
    .B1(_08974_),
    .B2(_13070_),
    .C1(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__o21ai_0 _21564_ (.A1(_13072_),
    .A2(_08910_),
    .B1(_08768_),
    .Y(_08977_));
 sky130_fd_sc_hd__nand4b_1 _21565_ (.A_N(_08798_),
    .B(_08919_),
    .C(_08976_),
    .D(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__a21o_2 _21566_ (.A1(_08549_),
    .A2(_08978_),
    .B1(net525),
    .X(_01024_));
 sky130_fd_sc_hd__a221o_1 _21567_ (.A1(net518),
    .A2(_08835_),
    .B1(_08824_),
    .B2(_13070_),
    .C1(_08752_),
    .X(_08979_));
 sky130_fd_sc_hd__o21ai_0 _21568_ (.A1(net466),
    .A2(_08929_),
    .B1(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__a21oi_2 _21569_ (.A1(_08969_),
    .A2(_08980_),
    .B1(_08778_),
    .Y(_01025_));
 sky130_fd_sc_hd__o22ai_1 _21570_ (.A1(_13072_),
    .A2(_08827_),
    .B1(_08862_),
    .B2(_13074_),
    .Y(_08981_));
 sky130_fd_sc_hd__a21oi_1 _21571_ (.A1(_08750_),
    .A2(_08842_),
    .B1(_10016_),
    .Y(_08982_));
 sky130_fd_sc_hd__o21ai_0 _21572_ (.A1(_13072_),
    .A2(_08982_),
    .B1(_08763_),
    .Y(_08983_));
 sky130_fd_sc_hd__nor3_1 _21573_ (.A(_13072_),
    .B(_13074_),
    .C(_08752_),
    .Y(_08984_));
 sky130_fd_sc_hd__a221o_1 _21574_ (.A1(net518),
    .A2(_08981_),
    .B1(_08983_),
    .B2(_08752_),
    .C1(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__a21oi_1 _21575_ (.A1(_08932_),
    .A2(_08985_),
    .B1(_10035_),
    .Y(_01026_));
 sky130_fd_sc_hd__a22oi_1 _21576_ (.A1(_13069_),
    .A2(_10027_),
    .B1(_08826_),
    .B2(_13074_),
    .Y(_08986_));
 sky130_fd_sc_hd__nor2_1 _21577_ (.A(net518),
    .B(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__o22ai_1 _21578_ (.A1(_13070_),
    .A2(_10027_),
    .B1(_08755_),
    .B2(_13074_),
    .Y(_08988_));
 sky130_fd_sc_hd__nor2_1 _21579_ (.A(_08747_),
    .B(_08846_),
    .Y(_08989_));
 sky130_fd_sc_hd__o21ai_0 _21580_ (.A1(_13070_),
    .A2(_08989_),
    .B1(_08749_),
    .Y(_08990_));
 sky130_fd_sc_hd__a21oi_1 _21581_ (.A1(_08834_),
    .A2(_08988_),
    .B1(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__a2111oi_1 _21582_ (.A1(_13070_),
    .A2(_08828_),
    .B1(_08987_),
    .C1(_08991_),
    .D1(_08762_),
    .Y(_08992_));
 sky130_fd_sc_hd__o21bai_1 _21583_ (.A1(_10571_),
    .A2(_08992_),
    .B1_N(net525),
    .Y(_01027_));
 sky130_fd_sc_hd__nand2_1 _21584_ (.A(_13074_),
    .B(_08756_),
    .Y(_08993_));
 sky130_fd_sc_hd__nand2_1 _21585_ (.A(_13069_),
    .B(_08862_),
    .Y(_08994_));
 sky130_fd_sc_hd__a21oi_1 _21586_ (.A1(_08860_),
    .A2(_08994_),
    .B1(net518),
    .Y(_08995_));
 sky130_fd_sc_hd__o21ai_0 _21587_ (.A1(_10016_),
    .A2(_08846_),
    .B1(_13072_),
    .Y(_08996_));
 sky130_fd_sc_hd__o21ai_0 _21588_ (.A1(net518),
    .A2(_08813_),
    .B1(_13070_),
    .Y(_08997_));
 sky130_fd_sc_hd__nand2_1 _21589_ (.A(_08996_),
    .B(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__a311oi_1 _21590_ (.A1(_13069_),
    .A2(_10016_),
    .A3(_08846_),
    .B1(_08995_),
    .C1(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__a21oi_1 _21591_ (.A1(_08993_),
    .A2(_08999_),
    .B1(_08778_),
    .Y(_01028_));
 sky130_fd_sc_hd__nor2_1 _21592_ (.A(_08857_),
    .B(_08921_),
    .Y(_09000_));
 sky130_fd_sc_hd__o211ai_1 _21593_ (.A1(_13070_),
    .A2(_09000_),
    .B1(_08967_),
    .C1(_08749_),
    .Y(_09001_));
 sky130_fd_sc_hd__nand3_1 _21594_ (.A(_08747_),
    .B(_08752_),
    .C(_08835_),
    .Y(_09002_));
 sky130_fd_sc_hd__o21ai_0 _21595_ (.A1(_08862_),
    .A2(_08837_),
    .B1(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand2_1 _21596_ (.A(net518),
    .B(_09003_),
    .Y(_09004_));
 sky130_fd_sc_hd__a31oi_2 _21597_ (.A1(_08849_),
    .A2(_09001_),
    .A3(_09004_),
    .B1(_08778_),
    .Y(_01029_));
 sky130_fd_sc_hd__o21ai_0 _21598_ (.A1(_08820_),
    .A2(_08828_),
    .B1(_13072_),
    .Y(_09005_));
 sky130_fd_sc_hd__o22ai_1 _21599_ (.A1(_08747_),
    .A2(_08793_),
    .B1(_08827_),
    .B2(net518),
    .Y(_09006_));
 sky130_fd_sc_hd__a21oi_1 _21600_ (.A1(_08752_),
    .A2(_08760_),
    .B1(_13070_),
    .Y(_09007_));
 sky130_fd_sc_hd__nor2_1 _21601_ (.A(net518),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__a21oi_1 _21602_ (.A1(_13069_),
    .A2(_09006_),
    .B1(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__nand3_1 _21603_ (.A(_08943_),
    .B(_09005_),
    .C(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__a21o_1 _21604_ (.A1(_08549_),
    .A2(_09010_),
    .B1(net525),
    .X(_01030_));
 sky130_fd_sc_hd__o21ai_0 _21605_ (.A1(_13072_),
    .A2(net518),
    .B1(_08826_),
    .Y(_09011_));
 sky130_fd_sc_hd__a21oi_1 _21606_ (.A1(_13069_),
    .A2(_08827_),
    .B1(_08762_),
    .Y(_09012_));
 sky130_fd_sc_hd__a21o_1 _21607_ (.A1(_10027_),
    .A2(_08824_),
    .B1(_08898_),
    .X(_09013_));
 sky130_fd_sc_hd__nand2_1 _21608_ (.A(_13072_),
    .B(_08782_),
    .Y(_09014_));
 sky130_fd_sc_hd__a21oi_1 _21609_ (.A1(_08971_),
    .A2(_09014_),
    .B1(_10016_),
    .Y(_09015_));
 sky130_fd_sc_hd__a21oi_1 _21610_ (.A1(_13074_),
    .A2(_09013_),
    .B1(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__a31oi_1 _21611_ (.A1(_09011_),
    .A2(_09012_),
    .A3(_09016_),
    .B1(_10035_),
    .Y(_01031_));
 sky130_fd_sc_hd__o2111ai_1 _21612_ (.A1(_08842_),
    .A2(_08845_),
    .B1(_08851_),
    .C1(_08871_),
    .D1(_10016_),
    .Y(_09017_));
 sky130_fd_sc_hd__o21ai_1 _21613_ (.A1(_10016_),
    .A2(_08954_),
    .B1(_09017_),
    .Y(_09018_));
 sky130_fd_sc_hd__a21oi_1 _21614_ (.A1(_08932_),
    .A2(_09018_),
    .B1(_10035_),
    .Y(_01032_));
 sky130_fd_sc_hd__nor2_2 _21615_ (.A(net525),
    .B(_08465_),
    .Y(_01033_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_918 ();
 sky130_fd_sc_hd__nand2_8 _21617_ (.A(_09907_),
    .B(_04982_),
    .Y(_09020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_917 ();
 sky130_fd_sc_hd__nor2_1 _21619_ (.A(_04988_),
    .B(_09020_),
    .Y(_01034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_916 ();
 sky130_fd_sc_hd__nor2_1 _21621_ (.A(_05062_),
    .B(_09020_),
    .Y(_01035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_915 ();
 sky130_fd_sc_hd__nor2_1 _21623_ (.A(_05077_),
    .B(_09020_),
    .Y(_01036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_914 ();
 sky130_fd_sc_hd__nor2_1 _21625_ (.A(_05087_),
    .B(_09020_),
    .Y(_01037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_913 ();
 sky130_fd_sc_hd__nor2_1 _21627_ (.A(_05095_),
    .B(_09020_),
    .Y(_01038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_912 ();
 sky130_fd_sc_hd__nor2_1 _21629_ (.A(_05102_),
    .B(_09020_),
    .Y(_01039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_911 ();
 sky130_fd_sc_hd__nor2_1 _21631_ (.A(_05112_),
    .B(_09020_),
    .Y(_01040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_910 ();
 sky130_fd_sc_hd__nor2_1 _21633_ (.A(_05121_),
    .B(_09020_),
    .Y(_01041_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_909 ();
 sky130_fd_sc_hd__nor2_1 _21635_ (.A(_05128_),
    .B(_09020_),
    .Y(_01042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_908 ();
 sky130_fd_sc_hd__nor2_1 _21637_ (.A(_05137_),
    .B(_09020_),
    .Y(_01043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_906 ();
 sky130_fd_sc_hd__nor2_1 _21640_ (.A(_05154_),
    .B(_09020_),
    .Y(_01044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_905 ();
 sky130_fd_sc_hd__nor2_1 _21642_ (.A(_04992_),
    .B(_09020_),
    .Y(_01045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_904 ();
 sky130_fd_sc_hd__nor2_1 _21644_ (.A(_05167_),
    .B(_09020_),
    .Y(_01046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_903 ();
 sky130_fd_sc_hd__nor2_1 _21646_ (.A(_05175_),
    .B(_09020_),
    .Y(_01047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_902 ();
 sky130_fd_sc_hd__nor2_1 _21648_ (.A(_05184_),
    .B(_09020_),
    .Y(_01048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_901 ();
 sky130_fd_sc_hd__nor2_1 _21650_ (.A(_05196_),
    .B(_09020_),
    .Y(_01049_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_900 ();
 sky130_fd_sc_hd__nor2_1 _21652_ (.A(_05206_),
    .B(_09020_),
    .Y(_01050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_899 ();
 sky130_fd_sc_hd__nor2_1 _21654_ (.A(_05214_),
    .B(_09020_),
    .Y(_01051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_898 ();
 sky130_fd_sc_hd__nor2_1 _21656_ (.A(_05224_),
    .B(_09020_),
    .Y(_01052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_897 ();
 sky130_fd_sc_hd__nor2_1 _21658_ (.A(_05236_),
    .B(_09020_),
    .Y(_01053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_895 ();
 sky130_fd_sc_hd__nor2_1 _21661_ (.A(_05243_),
    .B(_09020_),
    .Y(_01054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_894 ();
 sky130_fd_sc_hd__nor2_1 _21663_ (.A(_05251_),
    .B(_09020_),
    .Y(_01055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_893 ();
 sky130_fd_sc_hd__nor2_1 _21665_ (.A(_04995_),
    .B(_09020_),
    .Y(_01056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_892 ();
 sky130_fd_sc_hd__nor2_1 _21667_ (.A(_05260_),
    .B(_09020_),
    .Y(_01057_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_891 ();
 sky130_fd_sc_hd__nor2_1 _21669_ (.A(_05310_),
    .B(_09020_),
    .Y(_01058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_890 ();
 sky130_fd_sc_hd__nor2_1 _21671_ (.A(_05003_),
    .B(_09020_),
    .Y(_01059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_889 ();
 sky130_fd_sc_hd__nor2_1 _21673_ (.A(_05012_),
    .B(_09020_),
    .Y(_01060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_888 ();
 sky130_fd_sc_hd__nor2_1 _21675_ (.A(_05021_),
    .B(_09020_),
    .Y(_01061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_887 ();
 sky130_fd_sc_hd__nor2_1 _21677_ (.A(_05032_),
    .B(_09020_),
    .Y(_01062_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_886 ();
 sky130_fd_sc_hd__nor2_1 _21679_ (.A(_05039_),
    .B(_09020_),
    .Y(_01063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_885 ();
 sky130_fd_sc_hd__nor2_1 _21681_ (.A(_05048_),
    .B(_09020_),
    .Y(_01064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_884 ();
 sky130_fd_sc_hd__nor2_1 _21683_ (.A(_05055_),
    .B(_09020_),
    .Y(_01065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_883 ();
 sky130_fd_sc_hd__nand2_8 _21685_ (.A(_09956_),
    .B(_05313_),
    .Y(_09056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_882 ();
 sky130_fd_sc_hd__nor2_1 _21687_ (.A(_05317_),
    .B(_09056_),
    .Y(_01066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_881 ();
 sky130_fd_sc_hd__nor2_1 _21689_ (.A(_05388_),
    .B(_09056_),
    .Y(_01067_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_880 ();
 sky130_fd_sc_hd__nor2_1 _21691_ (.A(_05402_),
    .B(_09056_),
    .Y(_01068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_879 ();
 sky130_fd_sc_hd__nor2_1 _21693_ (.A(_05412_),
    .B(_09056_),
    .Y(_01069_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_878 ();
 sky130_fd_sc_hd__nor2_1 _21695_ (.A(_05419_),
    .B(_09056_),
    .Y(_01070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_877 ();
 sky130_fd_sc_hd__nor2_1 _21697_ (.A(_05426_),
    .B(_09056_),
    .Y(_01071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_876 ();
 sky130_fd_sc_hd__nor2_1 _21699_ (.A(_05438_),
    .B(_09056_),
    .Y(_01072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_875 ();
 sky130_fd_sc_hd__nor2_1 _21701_ (.A(_05447_),
    .B(_09056_),
    .Y(_01073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_874 ();
 sky130_fd_sc_hd__nor2_1 _21703_ (.A(_05453_),
    .B(_09056_),
    .Y(_01074_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_873 ();
 sky130_fd_sc_hd__nor2_1 _21705_ (.A(_05465_),
    .B(_09056_),
    .Y(_01075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_871 ();
 sky130_fd_sc_hd__nor2_1 _21708_ (.A(_05480_),
    .B(_09056_),
    .Y(_01076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_870 ();
 sky130_fd_sc_hd__nor2_1 _21710_ (.A(_05321_),
    .B(_09056_),
    .Y(_01077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_869 ();
 sky130_fd_sc_hd__nor2_1 _21712_ (.A(_05488_),
    .B(_09056_),
    .Y(_01078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_868 ();
 sky130_fd_sc_hd__nor2_1 _21714_ (.A(_05498_),
    .B(_09056_),
    .Y(_01079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_867 ();
 sky130_fd_sc_hd__nor2_1 _21716_ (.A(_05509_),
    .B(_09056_),
    .Y(_01080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_866 ();
 sky130_fd_sc_hd__nor2_1 _21718_ (.A(_05515_),
    .B(_09056_),
    .Y(_01081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_865 ();
 sky130_fd_sc_hd__nor2_1 _21720_ (.A(_05523_),
    .B(_09056_),
    .Y(_01082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_864 ();
 sky130_fd_sc_hd__nor2_1 _21722_ (.A(_05535_),
    .B(_09056_),
    .Y(_01083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_863 ();
 sky130_fd_sc_hd__nor2_1 _21724_ (.A(_05542_),
    .B(_09056_),
    .Y(_01084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_862 ();
 sky130_fd_sc_hd__nor2_1 _21726_ (.A(_05551_),
    .B(_09056_),
    .Y(_01085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_860 ();
 sky130_fd_sc_hd__nor2_1 _21729_ (.A(_05559_),
    .B(_09056_),
    .Y(_01086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_859 ();
 sky130_fd_sc_hd__nor2_1 _21731_ (.A(_05567_),
    .B(_09056_),
    .Y(_01087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_858 ();
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(_05324_),
    .B(_09056_),
    .Y(_01088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_857 ();
 sky130_fd_sc_hd__nor2_1 _21735_ (.A(_05573_),
    .B(_09056_),
    .Y(_01089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_856 ();
 sky130_fd_sc_hd__nor2_1 _21737_ (.A(_05611_),
    .B(_09056_),
    .Y(_01090_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_855 ();
 sky130_fd_sc_hd__nor2_1 _21739_ (.A(_05330_),
    .B(_09056_),
    .Y(_01091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_854 ();
 sky130_fd_sc_hd__nor2_1 _21741_ (.A(_05338_),
    .B(_09056_),
    .Y(_01092_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_853 ();
 sky130_fd_sc_hd__nor2_1 _21743_ (.A(_05347_),
    .B(_09056_),
    .Y(_01093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_852 ();
 sky130_fd_sc_hd__nor2_1 _21745_ (.A(_05354_),
    .B(_09056_),
    .Y(_01094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_851 ();
 sky130_fd_sc_hd__nor2_1 _21747_ (.A(_05360_),
    .B(_09056_),
    .Y(_01095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_850 ();
 sky130_fd_sc_hd__nor2_1 _21749_ (.A(_05371_),
    .B(_09056_),
    .Y(_01096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_849 ();
 sky130_fd_sc_hd__nor2_1 _21751_ (.A(_05380_),
    .B(_09056_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_8 _21752_ (.A(_09907_),
    .B(_05614_),
    .Y(_09091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_848 ();
 sky130_fd_sc_hd__nor2_1 _21754_ (.A(_04988_),
    .B(_09091_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_1 _21755_ (.A(_05062_),
    .B(_09091_),
    .Y(_01099_));
 sky130_fd_sc_hd__nor2_1 _21756_ (.A(_05077_),
    .B(_09091_),
    .Y(_01100_));
 sky130_fd_sc_hd__nor2_1 _21757_ (.A(_05087_),
    .B(_09091_),
    .Y(_01101_));
 sky130_fd_sc_hd__nor2_1 _21758_ (.A(_05095_),
    .B(_09091_),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_1 _21759_ (.A(_05102_),
    .B(_09091_),
    .Y(_01103_));
 sky130_fd_sc_hd__nor2_1 _21760_ (.A(_05112_),
    .B(_09091_),
    .Y(_01104_));
 sky130_fd_sc_hd__nor2_1 _21761_ (.A(_05121_),
    .B(_09091_),
    .Y(_01105_));
 sky130_fd_sc_hd__nor2_1 _21762_ (.A(_05128_),
    .B(_09091_),
    .Y(_01106_));
 sky130_fd_sc_hd__nor2_1 _21763_ (.A(_05137_),
    .B(_09091_),
    .Y(_01107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_847 ();
 sky130_fd_sc_hd__nor2_1 _21765_ (.A(_05154_),
    .B(_09091_),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _21766_ (.A(_04992_),
    .B(_09091_),
    .Y(_01109_));
 sky130_fd_sc_hd__nor2_1 _21767_ (.A(_05167_),
    .B(_09091_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2_1 _21768_ (.A(_05175_),
    .B(_09091_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_1 _21769_ (.A(_05184_),
    .B(_09091_),
    .Y(_01112_));
 sky130_fd_sc_hd__nor2_1 _21770_ (.A(_05196_),
    .B(_09091_),
    .Y(_01113_));
 sky130_fd_sc_hd__nor2_1 _21771_ (.A(_05206_),
    .B(_09091_),
    .Y(_01114_));
 sky130_fd_sc_hd__nor2_1 _21772_ (.A(_05214_),
    .B(_09091_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _21773_ (.A(_05224_),
    .B(_09091_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor2_1 _21774_ (.A(_05236_),
    .B(_09091_),
    .Y(_01117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_846 ();
 sky130_fd_sc_hd__nor2_1 _21776_ (.A(_05243_),
    .B(_09091_),
    .Y(_01118_));
 sky130_fd_sc_hd__nor2_1 _21777_ (.A(_05251_),
    .B(_09091_),
    .Y(_01119_));
 sky130_fd_sc_hd__nor2_1 _21778_ (.A(_04995_),
    .B(_09091_),
    .Y(_01120_));
 sky130_fd_sc_hd__nor2_1 _21779_ (.A(_05260_),
    .B(_09091_),
    .Y(_01121_));
 sky130_fd_sc_hd__nor2_1 _21780_ (.A(_05310_),
    .B(_09091_),
    .Y(_01122_));
 sky130_fd_sc_hd__nor2_1 _21781_ (.A(_05003_),
    .B(_09091_),
    .Y(_01123_));
 sky130_fd_sc_hd__nor2_1 _21782_ (.A(_05012_),
    .B(_09091_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _21783_ (.A(_05021_),
    .B(_09091_),
    .Y(_01125_));
 sky130_fd_sc_hd__nor2_1 _21784_ (.A(_05032_),
    .B(_09091_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_1 _21785_ (.A(_05039_),
    .B(_09091_),
    .Y(_01127_));
 sky130_fd_sc_hd__nor2_1 _21786_ (.A(_05048_),
    .B(_09091_),
    .Y(_01128_));
 sky130_fd_sc_hd__nor2_1 _21787_ (.A(_05055_),
    .B(_09091_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_8 _21788_ (.A(_09956_),
    .B(_05655_),
    .Y(_09095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_845 ();
 sky130_fd_sc_hd__nor2_1 _21790_ (.A(_05317_),
    .B(_09095_),
    .Y(_01130_));
 sky130_fd_sc_hd__nor2_1 _21791_ (.A(_05388_),
    .B(_09095_),
    .Y(_01131_));
 sky130_fd_sc_hd__nor2_1 _21792_ (.A(_05402_),
    .B(_09095_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_1 _21793_ (.A(_05412_),
    .B(_09095_),
    .Y(_01133_));
 sky130_fd_sc_hd__nor2_1 _21794_ (.A(_05419_),
    .B(_09095_),
    .Y(_01134_));
 sky130_fd_sc_hd__nor2_1 _21795_ (.A(_05426_),
    .B(_09095_),
    .Y(_01135_));
 sky130_fd_sc_hd__nor2_1 _21796_ (.A(_05438_),
    .B(_09095_),
    .Y(_01136_));
 sky130_fd_sc_hd__nor2_1 _21797_ (.A(_05447_),
    .B(_09095_),
    .Y(_01137_));
 sky130_fd_sc_hd__nor2_1 _21798_ (.A(_05453_),
    .B(_09095_),
    .Y(_01138_));
 sky130_fd_sc_hd__nor2_1 _21799_ (.A(_05465_),
    .B(_09095_),
    .Y(_01139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_844 ();
 sky130_fd_sc_hd__nor2_1 _21801_ (.A(_05480_),
    .B(_09095_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _21802_ (.A(_05321_),
    .B(_09095_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _21803_ (.A(_05488_),
    .B(_09095_),
    .Y(_01142_));
 sky130_fd_sc_hd__nor2_1 _21804_ (.A(_05498_),
    .B(_09095_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_1 _21805_ (.A(_05509_),
    .B(_09095_),
    .Y(_01144_));
 sky130_fd_sc_hd__nor2_1 _21806_ (.A(_05515_),
    .B(_09095_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _21807_ (.A(_05523_),
    .B(_09095_),
    .Y(_01146_));
 sky130_fd_sc_hd__nor2_1 _21808_ (.A(_05535_),
    .B(_09095_),
    .Y(_01147_));
 sky130_fd_sc_hd__nor2_1 _21809_ (.A(_05542_),
    .B(_09095_),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_1 _21810_ (.A(_05551_),
    .B(_09095_),
    .Y(_01149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_843 ();
 sky130_fd_sc_hd__nor2_1 _21812_ (.A(_05559_),
    .B(_09095_),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_1 _21813_ (.A(_05567_),
    .B(_09095_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _21814_ (.A(_05324_),
    .B(_09095_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor2_1 _21815_ (.A(_05573_),
    .B(_09095_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor2_1 _21816_ (.A(_05611_),
    .B(_09095_),
    .Y(_01154_));
 sky130_fd_sc_hd__nor2_1 _21817_ (.A(_05330_),
    .B(_09095_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _21818_ (.A(_05338_),
    .B(_09095_),
    .Y(_01156_));
 sky130_fd_sc_hd__nor2_1 _21819_ (.A(_05347_),
    .B(_09095_),
    .Y(_01157_));
 sky130_fd_sc_hd__nor2_1 _21820_ (.A(_05354_),
    .B(_09095_),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _21821_ (.A(_05360_),
    .B(_09095_),
    .Y(_01159_));
 sky130_fd_sc_hd__nor2_1 _21822_ (.A(_05371_),
    .B(_09095_),
    .Y(_01160_));
 sky130_fd_sc_hd__nor2_1 _21823_ (.A(_05380_),
    .B(_09095_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2_8 _21824_ (.A(_09907_),
    .B(_05696_),
    .Y(_09099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_842 ();
 sky130_fd_sc_hd__nor2_1 _21826_ (.A(_04988_),
    .B(_09099_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_1 _21827_ (.A(_05062_),
    .B(_09099_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_1 _21828_ (.A(_05077_),
    .B(_09099_),
    .Y(_01164_));
 sky130_fd_sc_hd__nor2_1 _21829_ (.A(_05087_),
    .B(_09099_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _21830_ (.A(_05095_),
    .B(_09099_),
    .Y(_01166_));
 sky130_fd_sc_hd__nor2_1 _21831_ (.A(_05102_),
    .B(_09099_),
    .Y(_01167_));
 sky130_fd_sc_hd__nor2_1 _21832_ (.A(_05112_),
    .B(_09099_),
    .Y(_01168_));
 sky130_fd_sc_hd__nor2_1 _21833_ (.A(_05121_),
    .B(_09099_),
    .Y(_01169_));
 sky130_fd_sc_hd__nor2_1 _21834_ (.A(_05128_),
    .B(_09099_),
    .Y(_01170_));
 sky130_fd_sc_hd__nor2_1 _21835_ (.A(_05137_),
    .B(_09099_),
    .Y(_01171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_841 ();
 sky130_fd_sc_hd__nor2_1 _21837_ (.A(_05154_),
    .B(_09099_),
    .Y(_01172_));
 sky130_fd_sc_hd__nor2_1 _21838_ (.A(_04992_),
    .B(_09099_),
    .Y(_01173_));
 sky130_fd_sc_hd__nor2_1 _21839_ (.A(_05167_),
    .B(_09099_),
    .Y(_01174_));
 sky130_fd_sc_hd__nor2_1 _21840_ (.A(_05175_),
    .B(_09099_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor2_1 _21841_ (.A(_05184_),
    .B(_09099_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2_1 _21842_ (.A(_05196_),
    .B(_09099_),
    .Y(_01177_));
 sky130_fd_sc_hd__nor2_1 _21843_ (.A(_05206_),
    .B(_09099_),
    .Y(_01178_));
 sky130_fd_sc_hd__nor2_1 _21844_ (.A(_05214_),
    .B(_09099_),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_1 _21845_ (.A(_05224_),
    .B(_09099_),
    .Y(_01180_));
 sky130_fd_sc_hd__nor2_1 _21846_ (.A(_05236_),
    .B(_09099_),
    .Y(_01181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_840 ();
 sky130_fd_sc_hd__nor2_1 _21848_ (.A(_05243_),
    .B(_09099_),
    .Y(_01182_));
 sky130_fd_sc_hd__nor2_1 _21849_ (.A(_05251_),
    .B(_09099_),
    .Y(_01183_));
 sky130_fd_sc_hd__nor2_1 _21850_ (.A(_04995_),
    .B(_09099_),
    .Y(_01184_));
 sky130_fd_sc_hd__nor2_1 _21851_ (.A(_05260_),
    .B(_09099_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_1 _21852_ (.A(_05310_),
    .B(_09099_),
    .Y(_01186_));
 sky130_fd_sc_hd__nor2_1 _21853_ (.A(_05003_),
    .B(_09099_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_1 _21854_ (.A(_05012_),
    .B(_09099_),
    .Y(_01188_));
 sky130_fd_sc_hd__nor2_1 _21855_ (.A(_05021_),
    .B(_09099_),
    .Y(_01189_));
 sky130_fd_sc_hd__nor2_1 _21856_ (.A(_05032_),
    .B(_09099_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _21857_ (.A(_05039_),
    .B(_09099_),
    .Y(_01191_));
 sky130_fd_sc_hd__nor2_1 _21858_ (.A(_05048_),
    .B(_09099_),
    .Y(_01192_));
 sky130_fd_sc_hd__nor2_1 _21859_ (.A(_05055_),
    .B(_09099_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_8 _21860_ (.A(_09956_),
    .B(_05737_),
    .Y(_09103_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_839 ();
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(_05317_),
    .B(_09103_),
    .Y(_01194_));
 sky130_fd_sc_hd__nor2_1 _21863_ (.A(_05388_),
    .B(_09103_),
    .Y(_01195_));
 sky130_fd_sc_hd__nor2_1 _21864_ (.A(_05402_),
    .B(_09103_),
    .Y(_01196_));
 sky130_fd_sc_hd__nor2_1 _21865_ (.A(_05412_),
    .B(_09103_),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_1 _21866_ (.A(_05419_),
    .B(_09103_),
    .Y(_01198_));
 sky130_fd_sc_hd__nor2_1 _21867_ (.A(_05426_),
    .B(_09103_),
    .Y(_01199_));
 sky130_fd_sc_hd__nor2_1 _21868_ (.A(_05438_),
    .B(_09103_),
    .Y(_01200_));
 sky130_fd_sc_hd__nor2_1 _21869_ (.A(_05447_),
    .B(_09103_),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _21870_ (.A(_05453_),
    .B(_09103_),
    .Y(_01202_));
 sky130_fd_sc_hd__nor2_1 _21871_ (.A(_05465_),
    .B(_09103_),
    .Y(_01203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_838 ();
 sky130_fd_sc_hd__nor2_1 _21873_ (.A(_05480_),
    .B(_09103_),
    .Y(_01204_));
 sky130_fd_sc_hd__nor2_1 _21874_ (.A(_05321_),
    .B(_09103_),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_1 _21875_ (.A(_05488_),
    .B(_09103_),
    .Y(_01206_));
 sky130_fd_sc_hd__nor2_1 _21876_ (.A(_05498_),
    .B(_09103_),
    .Y(_01207_));
 sky130_fd_sc_hd__nor2_1 _21877_ (.A(_05509_),
    .B(_09103_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _21878_ (.A(_05515_),
    .B(_09103_),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_1 _21879_ (.A(_05523_),
    .B(_09103_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor2_1 _21880_ (.A(_05535_),
    .B(_09103_),
    .Y(_01211_));
 sky130_fd_sc_hd__nor2_1 _21881_ (.A(_05542_),
    .B(_09103_),
    .Y(_01212_));
 sky130_fd_sc_hd__nor2_1 _21882_ (.A(_05551_),
    .B(_09103_),
    .Y(_01213_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_837 ();
 sky130_fd_sc_hd__nor2_1 _21884_ (.A(_05559_),
    .B(_09103_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_1 _21885_ (.A(_05567_),
    .B(_09103_),
    .Y(_01215_));
 sky130_fd_sc_hd__nor2_1 _21886_ (.A(_05324_),
    .B(_09103_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_1 _21887_ (.A(_05573_),
    .B(_09103_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _21888_ (.A(_05611_),
    .B(_09103_),
    .Y(_01218_));
 sky130_fd_sc_hd__nor2_1 _21889_ (.A(_05330_),
    .B(_09103_),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_1 _21890_ (.A(_05338_),
    .B(_09103_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor2_1 _21891_ (.A(_05347_),
    .B(_09103_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _21892_ (.A(_05354_),
    .B(_09103_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_1 _21893_ (.A(_05360_),
    .B(_09103_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_1 _21894_ (.A(_05371_),
    .B(_09103_),
    .Y(_01224_));
 sky130_fd_sc_hd__nor2_1 _21895_ (.A(_05380_),
    .B(_09103_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_8 _21896_ (.A(_09907_),
    .B(_05778_),
    .Y(_09107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_836 ();
 sky130_fd_sc_hd__nor2_1 _21898_ (.A(_04988_),
    .B(_09107_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _21899_ (.A(_05062_),
    .B(_09107_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor2_1 _21900_ (.A(_05077_),
    .B(_09107_),
    .Y(_01228_));
 sky130_fd_sc_hd__nor2_1 _21901_ (.A(_05087_),
    .B(_09107_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_1 _21902_ (.A(_05095_),
    .B(_09107_),
    .Y(_01230_));
 sky130_fd_sc_hd__nor2_1 _21903_ (.A(_05102_),
    .B(_09107_),
    .Y(_01231_));
 sky130_fd_sc_hd__nor2_1 _21904_ (.A(_05112_),
    .B(_09107_),
    .Y(_01232_));
 sky130_fd_sc_hd__nor2_1 _21905_ (.A(_05121_),
    .B(_09107_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_1 _21906_ (.A(_05128_),
    .B(_09107_),
    .Y(_01234_));
 sky130_fd_sc_hd__nor2_1 _21907_ (.A(_05137_),
    .B(_09107_),
    .Y(_01235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_835 ();
 sky130_fd_sc_hd__nor2_1 _21909_ (.A(_05154_),
    .B(_09107_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_1 _21910_ (.A(_04992_),
    .B(_09107_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _21911_ (.A(_05167_),
    .B(_09107_),
    .Y(_01238_));
 sky130_fd_sc_hd__nor2_1 _21912_ (.A(_05175_),
    .B(_09107_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _21913_ (.A(_05184_),
    .B(_09107_),
    .Y(_01240_));
 sky130_fd_sc_hd__nor2_1 _21914_ (.A(_05196_),
    .B(_09107_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_1 _21915_ (.A(_05206_),
    .B(_09107_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_1 _21916_ (.A(_05214_),
    .B(_09107_),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _21917_ (.A(_05224_),
    .B(_09107_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _21918_ (.A(_05236_),
    .B(_09107_),
    .Y(_01245_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_834 ();
 sky130_fd_sc_hd__nor2_1 _21920_ (.A(_05243_),
    .B(_09107_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _21921_ (.A(_05251_),
    .B(_09107_),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_1 _21922_ (.A(_04995_),
    .B(_09107_),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _21923_ (.A(_05260_),
    .B(_09107_),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_1 _21924_ (.A(_05310_),
    .B(_09107_),
    .Y(_01250_));
 sky130_fd_sc_hd__nor2_1 _21925_ (.A(_05003_),
    .B(_09107_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor2_1 _21926_ (.A(_05012_),
    .B(_09107_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _21927_ (.A(_05021_),
    .B(_09107_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor2_1 _21928_ (.A(_05032_),
    .B(_09107_),
    .Y(_01254_));
 sky130_fd_sc_hd__nor2_1 _21929_ (.A(_05039_),
    .B(_09107_),
    .Y(_01255_));
 sky130_fd_sc_hd__nor2_1 _21930_ (.A(_05048_),
    .B(_09107_),
    .Y(_01256_));
 sky130_fd_sc_hd__nor2_1 _21931_ (.A(_05055_),
    .B(_09107_),
    .Y(_01257_));
 sky130_fd_sc_hd__or3_4 _21932_ (.A(net762),
    .B(_09955_),
    .C(_09964_),
    .X(_09111_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_832 ();
 sky130_fd_sc_hd__nor2_1 _21935_ (.A(_05317_),
    .B(_09111_),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _21936_ (.A(_05388_),
    .B(_09111_),
    .Y(_01259_));
 sky130_fd_sc_hd__nor2_1 _21937_ (.A(_05402_),
    .B(_09111_),
    .Y(_01260_));
 sky130_fd_sc_hd__nor2_1 _21938_ (.A(_05412_),
    .B(_09111_),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_1 _21939_ (.A(_05419_),
    .B(_09111_),
    .Y(_01262_));
 sky130_fd_sc_hd__nor2_1 _21940_ (.A(_05426_),
    .B(_09111_),
    .Y(_01263_));
 sky130_fd_sc_hd__nor2_1 _21941_ (.A(_05438_),
    .B(_09111_),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_1 _21942_ (.A(_05447_),
    .B(_09111_),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _21943_ (.A(_05453_),
    .B(_09111_),
    .Y(_01266_));
 sky130_fd_sc_hd__nor2_1 _21944_ (.A(_05465_),
    .B(_09111_),
    .Y(_01267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_831 ();
 sky130_fd_sc_hd__nor2_1 _21946_ (.A(_05480_),
    .B(_09111_),
    .Y(_01268_));
 sky130_fd_sc_hd__nor2_1 _21947_ (.A(_05321_),
    .B(_09111_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_1 _21948_ (.A(_05488_),
    .B(_09111_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _21949_ (.A(_05498_),
    .B(_09111_),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_1 _21950_ (.A(_05509_),
    .B(_09111_),
    .Y(_01272_));
 sky130_fd_sc_hd__nor2_1 _21951_ (.A(_05515_),
    .B(_09111_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor2_1 _21952_ (.A(_05523_),
    .B(_09111_),
    .Y(_01274_));
 sky130_fd_sc_hd__nor2_1 _21953_ (.A(_05535_),
    .B(_09111_),
    .Y(_01275_));
 sky130_fd_sc_hd__nor2_1 _21954_ (.A(_05542_),
    .B(_09111_),
    .Y(_01276_));
 sky130_fd_sc_hd__nor2_1 _21955_ (.A(_05551_),
    .B(_09111_),
    .Y(_01277_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_830 ();
 sky130_fd_sc_hd__nor2_1 _21957_ (.A(_05559_),
    .B(_09111_),
    .Y(_01278_));
 sky130_fd_sc_hd__nor2_1 _21958_ (.A(_05567_),
    .B(_09111_),
    .Y(_01279_));
 sky130_fd_sc_hd__nor2_1 _21959_ (.A(_05324_),
    .B(_09111_),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_1 _21960_ (.A(_05573_),
    .B(_09111_),
    .Y(_01281_));
 sky130_fd_sc_hd__nor2_1 _21961_ (.A(_05611_),
    .B(_09111_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor2_1 _21962_ (.A(_05330_),
    .B(_09111_),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_1 _21963_ (.A(_05338_),
    .B(_09111_),
    .Y(_01284_));
 sky130_fd_sc_hd__nor2_1 _21964_ (.A(_05347_),
    .B(_09111_),
    .Y(_01285_));
 sky130_fd_sc_hd__nor2_1 _21965_ (.A(_05354_),
    .B(_09111_),
    .Y(_01286_));
 sky130_fd_sc_hd__nor2_1 _21966_ (.A(_05360_),
    .B(_09111_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_1 _21967_ (.A(_05371_),
    .B(_09111_),
    .Y(_01288_));
 sky130_fd_sc_hd__nor2_1 _21968_ (.A(_05380_),
    .B(_09111_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_8 _21969_ (.A(_09913_),
    .B(_04982_),
    .Y(_09116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_829 ();
 sky130_fd_sc_hd__nor2_1 _21971_ (.A(_04988_),
    .B(_09116_),
    .Y(_01290_));
 sky130_fd_sc_hd__nor2_1 _21972_ (.A(_05062_),
    .B(_09116_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_1 _21973_ (.A(_05077_),
    .B(_09116_),
    .Y(_01292_));
 sky130_fd_sc_hd__nor2_1 _21974_ (.A(_05087_),
    .B(_09116_),
    .Y(_01293_));
 sky130_fd_sc_hd__nor2_1 _21975_ (.A(_05095_),
    .B(_09116_),
    .Y(_01294_));
 sky130_fd_sc_hd__nor2_1 _21976_ (.A(_05102_),
    .B(_09116_),
    .Y(_01295_));
 sky130_fd_sc_hd__nor2_1 _21977_ (.A(_05112_),
    .B(_09116_),
    .Y(_01296_));
 sky130_fd_sc_hd__nor2_1 _21978_ (.A(_05121_),
    .B(_09116_),
    .Y(_01297_));
 sky130_fd_sc_hd__nor2_1 _21979_ (.A(_05128_),
    .B(_09116_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_1 _21980_ (.A(_05137_),
    .B(_09116_),
    .Y(_01299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_828 ();
 sky130_fd_sc_hd__nor2_1 _21982_ (.A(_05154_),
    .B(_09116_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _21983_ (.A(_04992_),
    .B(_09116_),
    .Y(_01301_));
 sky130_fd_sc_hd__nor2_1 _21984_ (.A(_05167_),
    .B(_09116_),
    .Y(_01302_));
 sky130_fd_sc_hd__nor2_1 _21985_ (.A(_05175_),
    .B(_09116_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_1 _21986_ (.A(_05184_),
    .B(_09116_),
    .Y(_01304_));
 sky130_fd_sc_hd__nor2_1 _21987_ (.A(_05196_),
    .B(_09116_),
    .Y(_01305_));
 sky130_fd_sc_hd__nor2_1 _21988_ (.A(_05206_),
    .B(_09116_),
    .Y(_01306_));
 sky130_fd_sc_hd__nor2_1 _21989_ (.A(_05214_),
    .B(_09116_),
    .Y(_01307_));
 sky130_fd_sc_hd__nor2_1 _21990_ (.A(_05224_),
    .B(_09116_),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_1 _21991_ (.A(_05236_),
    .B(_09116_),
    .Y(_01309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_827 ();
 sky130_fd_sc_hd__nor2_1 _21993_ (.A(_05243_),
    .B(_09116_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor2_1 _21994_ (.A(_05251_),
    .B(_09116_),
    .Y(_01311_));
 sky130_fd_sc_hd__nor2_1 _21995_ (.A(_04995_),
    .B(_09116_),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _21996_ (.A(_05260_),
    .B(_09116_),
    .Y(_01313_));
 sky130_fd_sc_hd__nor2_1 _21997_ (.A(_05310_),
    .B(_09116_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_1 _21998_ (.A(_05003_),
    .B(_09116_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2_1 _21999_ (.A(_05012_),
    .B(_09116_),
    .Y(_01316_));
 sky130_fd_sc_hd__nor2_1 _22000_ (.A(_05021_),
    .B(_09116_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_1 _22001_ (.A(_05032_),
    .B(_09116_),
    .Y(_01318_));
 sky130_fd_sc_hd__nor2_1 _22002_ (.A(_05039_),
    .B(_09116_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_1 _22003_ (.A(_05048_),
    .B(_09116_),
    .Y(_01320_));
 sky130_fd_sc_hd__nor2_1 _22004_ (.A(_05055_),
    .B(_09116_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_8 _22005_ (.A(_09966_),
    .B(_05313_),
    .Y(_09120_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_826 ();
 sky130_fd_sc_hd__nor2_1 _22007_ (.A(_05317_),
    .B(_09120_),
    .Y(_01322_));
 sky130_fd_sc_hd__nor2_1 _22008_ (.A(_05388_),
    .B(_09120_),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2_1 _22009_ (.A(_05402_),
    .B(_09120_),
    .Y(_01324_));
 sky130_fd_sc_hd__nor2_1 _22010_ (.A(_05412_),
    .B(_09120_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_1 _22011_ (.A(_05419_),
    .B(_09120_),
    .Y(_01326_));
 sky130_fd_sc_hd__nor2_1 _22012_ (.A(_05426_),
    .B(_09120_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_1 _22013_ (.A(_05438_),
    .B(_09120_),
    .Y(_01328_));
 sky130_fd_sc_hd__nor2_1 _22014_ (.A(_05447_),
    .B(_09120_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _22015_ (.A(_05453_),
    .B(_09120_),
    .Y(_01330_));
 sky130_fd_sc_hd__nor2_1 _22016_ (.A(_05465_),
    .B(_09120_),
    .Y(_01331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_825 ();
 sky130_fd_sc_hd__nor2_1 _22018_ (.A(_05480_),
    .B(_09120_),
    .Y(_01332_));
 sky130_fd_sc_hd__nor2_1 _22019_ (.A(_05321_),
    .B(_09120_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2_1 _22020_ (.A(_05488_),
    .B(_09120_),
    .Y(_01334_));
 sky130_fd_sc_hd__nor2_1 _22021_ (.A(_05498_),
    .B(_09120_),
    .Y(_01335_));
 sky130_fd_sc_hd__nor2_1 _22022_ (.A(_05509_),
    .B(_09120_),
    .Y(_01336_));
 sky130_fd_sc_hd__nor2_1 _22023_ (.A(_05515_),
    .B(_09120_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2_1 _22024_ (.A(_05523_),
    .B(_09120_),
    .Y(_01338_));
 sky130_fd_sc_hd__nor2_1 _22025_ (.A(_05535_),
    .B(_09120_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2_1 _22026_ (.A(_05542_),
    .B(_09120_),
    .Y(_01340_));
 sky130_fd_sc_hd__nor2_1 _22027_ (.A(_05551_),
    .B(_09120_),
    .Y(_01341_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_824 ();
 sky130_fd_sc_hd__nor2_1 _22029_ (.A(_05559_),
    .B(_09120_),
    .Y(_01342_));
 sky130_fd_sc_hd__nor2_1 _22030_ (.A(_05567_),
    .B(_09120_),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_1 _22031_ (.A(_05324_),
    .B(_09120_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _22032_ (.A(_05573_),
    .B(_09120_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _22033_ (.A(_05611_),
    .B(_09120_),
    .Y(_01346_));
 sky130_fd_sc_hd__nor2_1 _22034_ (.A(_05330_),
    .B(_09120_),
    .Y(_01347_));
 sky130_fd_sc_hd__nor2_1 _22035_ (.A(_05338_),
    .B(_09120_),
    .Y(_01348_));
 sky130_fd_sc_hd__nor2_1 _22036_ (.A(_05347_),
    .B(_09120_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2_1 _22037_ (.A(_05354_),
    .B(_09120_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor2_1 _22038_ (.A(_05360_),
    .B(_09120_),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2_1 _22039_ (.A(_05371_),
    .B(_09120_),
    .Y(_01352_));
 sky130_fd_sc_hd__nor2_1 _22040_ (.A(_05380_),
    .B(_09120_),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_8 _22041_ (.A(_09913_),
    .B(_05614_),
    .Y(_09124_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_823 ();
 sky130_fd_sc_hd__nor2_1 _22043_ (.A(_04988_),
    .B(_09124_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor2_1 _22044_ (.A(_05062_),
    .B(_09124_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2_1 _22045_ (.A(_05077_),
    .B(_09124_),
    .Y(_01356_));
 sky130_fd_sc_hd__nor2_1 _22046_ (.A(_05087_),
    .B(_09124_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_1 _22047_ (.A(_05095_),
    .B(_09124_),
    .Y(_01358_));
 sky130_fd_sc_hd__nor2_1 _22048_ (.A(_05102_),
    .B(_09124_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _22049_ (.A(_05112_),
    .B(_09124_),
    .Y(_01360_));
 sky130_fd_sc_hd__nor2_1 _22050_ (.A(_05121_),
    .B(_09124_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2_1 _22051_ (.A(_05128_),
    .B(_09124_),
    .Y(_01362_));
 sky130_fd_sc_hd__nor2_1 _22052_ (.A(_05137_),
    .B(_09124_),
    .Y(_01363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_822 ();
 sky130_fd_sc_hd__nor2_1 _22054_ (.A(_05154_),
    .B(_09124_),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_1 _22055_ (.A(_04992_),
    .B(_09124_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_1 _22056_ (.A(_05167_),
    .B(_09124_),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_1 _22057_ (.A(_05175_),
    .B(_09124_),
    .Y(_01367_));
 sky130_fd_sc_hd__nor2_1 _22058_ (.A(_05184_),
    .B(_09124_),
    .Y(_01368_));
 sky130_fd_sc_hd__nor2_1 _22059_ (.A(_05196_),
    .B(_09124_),
    .Y(_01369_));
 sky130_fd_sc_hd__nor2_1 _22060_ (.A(_05206_),
    .B(_09124_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _22061_ (.A(_05214_),
    .B(_09124_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_1 _22062_ (.A(_05224_),
    .B(_09124_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_1 _22063_ (.A(_05236_),
    .B(_09124_),
    .Y(_01373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_821 ();
 sky130_fd_sc_hd__nor2_1 _22065_ (.A(_05243_),
    .B(_09124_),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_1 _22066_ (.A(_05251_),
    .B(_09124_),
    .Y(_01375_));
 sky130_fd_sc_hd__nor2_1 _22067_ (.A(_04995_),
    .B(_09124_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _22068_ (.A(_05260_),
    .B(_09124_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _22069_ (.A(_05310_),
    .B(_09124_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_1 _22070_ (.A(_05003_),
    .B(_09124_),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_1 _22071_ (.A(_05012_),
    .B(_09124_),
    .Y(_01380_));
 sky130_fd_sc_hd__nor2_1 _22072_ (.A(_05021_),
    .B(_09124_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _22073_ (.A(_05032_),
    .B(_09124_),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_1 _22074_ (.A(_05039_),
    .B(_09124_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _22075_ (.A(_05048_),
    .B(_09124_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_1 _22076_ (.A(_05055_),
    .B(_09124_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_8 _22077_ (.A(_09966_),
    .B(_05655_),
    .Y(_09128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_820 ();
 sky130_fd_sc_hd__nor2_1 _22079_ (.A(_05317_),
    .B(_09128_),
    .Y(_01386_));
 sky130_fd_sc_hd__nor2_1 _22080_ (.A(_05388_),
    .B(_09128_),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_1 _22081_ (.A(_05402_),
    .B(_09128_),
    .Y(_01388_));
 sky130_fd_sc_hd__nor2_1 _22082_ (.A(_05412_),
    .B(_09128_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _22083_ (.A(_05419_),
    .B(_09128_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_1 _22084_ (.A(_05426_),
    .B(_09128_),
    .Y(_01391_));
 sky130_fd_sc_hd__nor2_1 _22085_ (.A(_05438_),
    .B(_09128_),
    .Y(_01392_));
 sky130_fd_sc_hd__nor2_1 _22086_ (.A(_05447_),
    .B(_09128_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _22087_ (.A(_05453_),
    .B(_09128_),
    .Y(_01394_));
 sky130_fd_sc_hd__nor2_1 _22088_ (.A(_05465_),
    .B(_09128_),
    .Y(_01395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_819 ();
 sky130_fd_sc_hd__nor2_1 _22090_ (.A(_05480_),
    .B(_09128_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _22091_ (.A(_05321_),
    .B(_09128_),
    .Y(_01397_));
 sky130_fd_sc_hd__nor2_1 _22092_ (.A(_05488_),
    .B(_09128_),
    .Y(_01398_));
 sky130_fd_sc_hd__nor2_1 _22093_ (.A(_05498_),
    .B(_09128_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor2_1 _22094_ (.A(_05509_),
    .B(_09128_),
    .Y(_01400_));
 sky130_fd_sc_hd__nor2_1 _22095_ (.A(_05515_),
    .B(_09128_),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_1 _22096_ (.A(_05523_),
    .B(_09128_),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_1 _22097_ (.A(_05535_),
    .B(_09128_),
    .Y(_01403_));
 sky130_fd_sc_hd__nor2_1 _22098_ (.A(_05542_),
    .B(_09128_),
    .Y(_01404_));
 sky130_fd_sc_hd__nor2_1 _22099_ (.A(_05551_),
    .B(_09128_),
    .Y(_01405_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_818 ();
 sky130_fd_sc_hd__nor2_1 _22101_ (.A(_05559_),
    .B(_09128_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _22102_ (.A(_05567_),
    .B(_09128_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _22103_ (.A(_05324_),
    .B(_09128_),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_1 _22104_ (.A(_05573_),
    .B(_09128_),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_1 _22105_ (.A(_05611_),
    .B(_09128_),
    .Y(_01410_));
 sky130_fd_sc_hd__nor2_1 _22106_ (.A(_05330_),
    .B(_09128_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor2_1 _22107_ (.A(_05338_),
    .B(_09128_),
    .Y(_01412_));
 sky130_fd_sc_hd__nor2_1 _22108_ (.A(_05347_),
    .B(_09128_),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_1 _22109_ (.A(_05354_),
    .B(_09128_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _22110_ (.A(_05360_),
    .B(_09128_),
    .Y(_01415_));
 sky130_fd_sc_hd__nor2_1 _22111_ (.A(_05371_),
    .B(_09128_),
    .Y(_01416_));
 sky130_fd_sc_hd__nor2_1 _22112_ (.A(_05380_),
    .B(_09128_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_8 _22113_ (.A(_09913_),
    .B(_05696_),
    .Y(_09132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_817 ();
 sky130_fd_sc_hd__nor2_1 _22115_ (.A(_04988_),
    .B(_09132_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _22116_ (.A(_05062_),
    .B(_09132_),
    .Y(_01419_));
 sky130_fd_sc_hd__nor2_1 _22117_ (.A(_05077_),
    .B(_09132_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_1 _22118_ (.A(_05087_),
    .B(_09132_),
    .Y(_01421_));
 sky130_fd_sc_hd__nor2_1 _22119_ (.A(_05095_),
    .B(_09132_),
    .Y(_01422_));
 sky130_fd_sc_hd__nor2_1 _22120_ (.A(_05102_),
    .B(_09132_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _22121_ (.A(_05112_),
    .B(_09132_),
    .Y(_01424_));
 sky130_fd_sc_hd__nor2_1 _22122_ (.A(_05121_),
    .B(_09132_),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_1 _22123_ (.A(_05128_),
    .B(_09132_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_1 _22124_ (.A(_05137_),
    .B(_09132_),
    .Y(_01427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_816 ();
 sky130_fd_sc_hd__nor2_1 _22126_ (.A(_05154_),
    .B(_09132_),
    .Y(_01428_));
 sky130_fd_sc_hd__nor2_1 _22127_ (.A(_04992_),
    .B(_09132_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _22128_ (.A(_05167_),
    .B(_09132_),
    .Y(_01430_));
 sky130_fd_sc_hd__nor2_1 _22129_ (.A(_05175_),
    .B(_09132_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_1 _22130_ (.A(_05184_),
    .B(_09132_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_1 _22131_ (.A(_05196_),
    .B(_09132_),
    .Y(_01433_));
 sky130_fd_sc_hd__nor2_1 _22132_ (.A(_05206_),
    .B(_09132_),
    .Y(_01434_));
 sky130_fd_sc_hd__nor2_1 _22133_ (.A(_05214_),
    .B(_09132_),
    .Y(_01435_));
 sky130_fd_sc_hd__nor2_1 _22134_ (.A(_05224_),
    .B(_09132_),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_1 _22135_ (.A(_05236_),
    .B(_09132_),
    .Y(_01437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_815 ();
 sky130_fd_sc_hd__nor2_1 _22137_ (.A(_05243_),
    .B(_09132_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _22138_ (.A(_05251_),
    .B(_09132_),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_1 _22139_ (.A(_04995_),
    .B(_09132_),
    .Y(_01440_));
 sky130_fd_sc_hd__nor2_1 _22140_ (.A(_05260_),
    .B(_09132_),
    .Y(_01441_));
 sky130_fd_sc_hd__nor2_1 _22141_ (.A(_05310_),
    .B(_09132_),
    .Y(_01442_));
 sky130_fd_sc_hd__nor2_1 _22142_ (.A(_05003_),
    .B(_09132_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2_1 _22143_ (.A(_05012_),
    .B(_09132_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _22144_ (.A(_05021_),
    .B(_09132_),
    .Y(_01445_));
 sky130_fd_sc_hd__nor2_1 _22145_ (.A(_05032_),
    .B(_09132_),
    .Y(_01446_));
 sky130_fd_sc_hd__nor2_1 _22146_ (.A(_05039_),
    .B(_09132_),
    .Y(_01447_));
 sky130_fd_sc_hd__nor2_1 _22147_ (.A(_05048_),
    .B(_09132_),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_1 _22148_ (.A(_05055_),
    .B(_09132_),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_8 _22149_ (.A(_09966_),
    .B(_05737_),
    .Y(_09136_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_814 ();
 sky130_fd_sc_hd__nor2_1 _22151_ (.A(_05317_),
    .B(_09136_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _22152_ (.A(_05388_),
    .B(_09136_),
    .Y(_01451_));
 sky130_fd_sc_hd__nor2_1 _22153_ (.A(_05402_),
    .B(_09136_),
    .Y(_01452_));
 sky130_fd_sc_hd__nor2_1 _22154_ (.A(_05412_),
    .B(_09136_),
    .Y(_01453_));
 sky130_fd_sc_hd__nor2_1 _22155_ (.A(_05419_),
    .B(_09136_),
    .Y(_01454_));
 sky130_fd_sc_hd__nor2_1 _22156_ (.A(_05426_),
    .B(_09136_),
    .Y(_01455_));
 sky130_fd_sc_hd__nor2_1 _22157_ (.A(_05438_),
    .B(_09136_),
    .Y(_01456_));
 sky130_fd_sc_hd__nor2_1 _22158_ (.A(_05447_),
    .B(_09136_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor2_1 _22159_ (.A(_05453_),
    .B(_09136_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_1 _22160_ (.A(_05465_),
    .B(_09136_),
    .Y(_01459_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_813 ();
 sky130_fd_sc_hd__nor2_1 _22162_ (.A(_05480_),
    .B(_09136_),
    .Y(_01460_));
 sky130_fd_sc_hd__nor2_1 _22163_ (.A(_05321_),
    .B(_09136_),
    .Y(_01461_));
 sky130_fd_sc_hd__nor2_1 _22164_ (.A(_05488_),
    .B(_09136_),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_1 _22165_ (.A(_05498_),
    .B(_09136_),
    .Y(_01463_));
 sky130_fd_sc_hd__nor2_1 _22166_ (.A(_05509_),
    .B(_09136_),
    .Y(_01464_));
 sky130_fd_sc_hd__nor2_1 _22167_ (.A(_05515_),
    .B(_09136_),
    .Y(_01465_));
 sky130_fd_sc_hd__nor2_1 _22168_ (.A(_05523_),
    .B(_09136_),
    .Y(_01466_));
 sky130_fd_sc_hd__nor2_1 _22169_ (.A(_05535_),
    .B(_09136_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _22170_ (.A(_05542_),
    .B(_09136_),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_1 _22171_ (.A(_05551_),
    .B(_09136_),
    .Y(_01469_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_812 ();
 sky130_fd_sc_hd__nor2_1 _22173_ (.A(_05559_),
    .B(_09136_),
    .Y(_01470_));
 sky130_fd_sc_hd__nor2_1 _22174_ (.A(_05567_),
    .B(_09136_),
    .Y(_01471_));
 sky130_fd_sc_hd__nor2_1 _22175_ (.A(_05324_),
    .B(_09136_),
    .Y(_01472_));
 sky130_fd_sc_hd__nor2_1 _22176_ (.A(_05573_),
    .B(_09136_),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_1 _22177_ (.A(_05611_),
    .B(_09136_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor2_1 _22178_ (.A(_05330_),
    .B(_09136_),
    .Y(_01475_));
 sky130_fd_sc_hd__nor2_1 _22179_ (.A(_05338_),
    .B(_09136_),
    .Y(_01476_));
 sky130_fd_sc_hd__nor2_1 _22180_ (.A(_05347_),
    .B(_09136_),
    .Y(_01477_));
 sky130_fd_sc_hd__nor2_1 _22181_ (.A(_05354_),
    .B(_09136_),
    .Y(_01478_));
 sky130_fd_sc_hd__nor2_1 _22182_ (.A(_05360_),
    .B(_09136_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_1 _22183_ (.A(_05371_),
    .B(_09136_),
    .Y(_01480_));
 sky130_fd_sc_hd__nor2_1 _22184_ (.A(_05380_),
    .B(_09136_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand2_8 _22185_ (.A(_09913_),
    .B(_05778_),
    .Y(_09140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_811 ();
 sky130_fd_sc_hd__nor2_1 _22187_ (.A(_04988_),
    .B(_09140_),
    .Y(_01482_));
 sky130_fd_sc_hd__nor2_1 _22188_ (.A(_05062_),
    .B(_09140_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _22189_ (.A(_05077_),
    .B(_09140_),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_1 _22190_ (.A(_05087_),
    .B(_09140_),
    .Y(_01485_));
 sky130_fd_sc_hd__nor2_1 _22191_ (.A(_05095_),
    .B(_09140_),
    .Y(_01486_));
 sky130_fd_sc_hd__nor2_1 _22192_ (.A(_05102_),
    .B(_09140_),
    .Y(_01487_));
 sky130_fd_sc_hd__nor2_1 _22193_ (.A(_05112_),
    .B(_09140_),
    .Y(_01488_));
 sky130_fd_sc_hd__nor2_1 _22194_ (.A(_05121_),
    .B(_09140_),
    .Y(_01489_));
 sky130_fd_sc_hd__nor2_1 _22195_ (.A(_05128_),
    .B(_09140_),
    .Y(_01490_));
 sky130_fd_sc_hd__nor2_1 _22196_ (.A(_05137_),
    .B(_09140_),
    .Y(_01491_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_810 ();
 sky130_fd_sc_hd__nor2_1 _22198_ (.A(_05154_),
    .B(_09140_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_1 _22199_ (.A(_04992_),
    .B(_09140_),
    .Y(_01493_));
 sky130_fd_sc_hd__nor2_1 _22200_ (.A(_05167_),
    .B(_09140_),
    .Y(_01494_));
 sky130_fd_sc_hd__nor2_1 _22201_ (.A(_05175_),
    .B(_09140_),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_1 _22202_ (.A(_05184_),
    .B(_09140_),
    .Y(_01496_));
 sky130_fd_sc_hd__nor2_1 _22203_ (.A(_05196_),
    .B(_09140_),
    .Y(_01497_));
 sky130_fd_sc_hd__nor2_1 _22204_ (.A(_05206_),
    .B(_09140_),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_1 _22205_ (.A(_05214_),
    .B(_09140_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _22206_ (.A(_05224_),
    .B(_09140_),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_1 _22207_ (.A(_05236_),
    .B(_09140_),
    .Y(_01501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_809 ();
 sky130_fd_sc_hd__nor2_1 _22209_ (.A(_05243_),
    .B(_09140_),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _22210_ (.A(_05251_),
    .B(_09140_),
    .Y(_01503_));
 sky130_fd_sc_hd__nor2_1 _22211_ (.A(_04995_),
    .B(_09140_),
    .Y(_01504_));
 sky130_fd_sc_hd__nor2_1 _22212_ (.A(_05260_),
    .B(_09140_),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_1 _22213_ (.A(_05310_),
    .B(_09140_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_1 _22214_ (.A(_05003_),
    .B(_09140_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_1 _22215_ (.A(_05012_),
    .B(_09140_),
    .Y(_01508_));
 sky130_fd_sc_hd__nor2_1 _22216_ (.A(_05021_),
    .B(_09140_),
    .Y(_01509_));
 sky130_fd_sc_hd__nor2_1 _22217_ (.A(_05032_),
    .B(_09140_),
    .Y(_01510_));
 sky130_fd_sc_hd__nor2_1 _22218_ (.A(_05039_),
    .B(_09140_),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_1 _22219_ (.A(_05048_),
    .B(_09140_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_1 _22220_ (.A(_05055_),
    .B(_09140_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_8 _22221_ (.A(_09966_),
    .B(_06133_),
    .Y(_09144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_808 ();
 sky130_fd_sc_hd__nor2_1 _22223_ (.A(_05317_),
    .B(_09144_),
    .Y(_01514_));
 sky130_fd_sc_hd__nor2_1 _22224_ (.A(_05388_),
    .B(_09144_),
    .Y(_01515_));
 sky130_fd_sc_hd__nor2_1 _22225_ (.A(_05402_),
    .B(_09144_),
    .Y(_01516_));
 sky130_fd_sc_hd__nor2_1 _22226_ (.A(_05412_),
    .B(_09144_),
    .Y(_01517_));
 sky130_fd_sc_hd__nor2_1 _22227_ (.A(_05419_),
    .B(_09144_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor2_1 _22228_ (.A(_05426_),
    .B(_09144_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor2_1 _22229_ (.A(_05438_),
    .B(_09144_),
    .Y(_01520_));
 sky130_fd_sc_hd__nor2_1 _22230_ (.A(_05447_),
    .B(_09144_),
    .Y(_01521_));
 sky130_fd_sc_hd__nor2_1 _22231_ (.A(_05453_),
    .B(_09144_),
    .Y(_01522_));
 sky130_fd_sc_hd__nor2_1 _22232_ (.A(_05465_),
    .B(_09144_),
    .Y(_01523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_807 ();
 sky130_fd_sc_hd__nor2_1 _22234_ (.A(_05480_),
    .B(_09144_),
    .Y(_01524_));
 sky130_fd_sc_hd__nor2_1 _22235_ (.A(_05321_),
    .B(_09144_),
    .Y(_01525_));
 sky130_fd_sc_hd__nor2_1 _22236_ (.A(_05488_),
    .B(_09144_),
    .Y(_01526_));
 sky130_fd_sc_hd__nor2_1 _22237_ (.A(_05498_),
    .B(_09144_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _22238_ (.A(_05509_),
    .B(_09144_),
    .Y(_01528_));
 sky130_fd_sc_hd__nor2_1 _22239_ (.A(_05515_),
    .B(_09144_),
    .Y(_01529_));
 sky130_fd_sc_hd__nor2_1 _22240_ (.A(_05523_),
    .B(_09144_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _22241_ (.A(_05535_),
    .B(_09144_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _22242_ (.A(_05542_),
    .B(_09144_),
    .Y(_01532_));
 sky130_fd_sc_hd__nor2_1 _22243_ (.A(_05551_),
    .B(_09144_),
    .Y(_01533_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_806 ();
 sky130_fd_sc_hd__nor2_1 _22245_ (.A(_05559_),
    .B(_09144_),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _22246_ (.A(_05567_),
    .B(_09144_),
    .Y(_01535_));
 sky130_fd_sc_hd__nor2_1 _22247_ (.A(_05324_),
    .B(_09144_),
    .Y(_01536_));
 sky130_fd_sc_hd__nor2_1 _22248_ (.A(_05573_),
    .B(_09144_),
    .Y(_01537_));
 sky130_fd_sc_hd__nor2_1 _22249_ (.A(_05611_),
    .B(_09144_),
    .Y(_01538_));
 sky130_fd_sc_hd__nor2_1 _22250_ (.A(_05330_),
    .B(_09144_),
    .Y(_01539_));
 sky130_fd_sc_hd__nor2_1 _22251_ (.A(_05338_),
    .B(_09144_),
    .Y(_01540_));
 sky130_fd_sc_hd__nor2_1 _22252_ (.A(_05347_),
    .B(_09144_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _22253_ (.A(_05354_),
    .B(_09144_),
    .Y(_01542_));
 sky130_fd_sc_hd__nor2_1 _22254_ (.A(_05360_),
    .B(_09144_),
    .Y(_01543_));
 sky130_fd_sc_hd__nor2_1 _22255_ (.A(_05371_),
    .B(_09144_),
    .Y(_01544_));
 sky130_fd_sc_hd__nor2_1 _22256_ (.A(_05380_),
    .B(_09144_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_8 _22257_ (.A(_09921_),
    .B(_04982_),
    .Y(_09148_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_805 ();
 sky130_fd_sc_hd__nor2_1 _22259_ (.A(_04988_),
    .B(_09148_),
    .Y(_01546_));
 sky130_fd_sc_hd__nor2_1 _22260_ (.A(_05062_),
    .B(_09148_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_1 _22261_ (.A(_05077_),
    .B(_09148_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _22262_ (.A(_05087_),
    .B(_09148_),
    .Y(_01549_));
 sky130_fd_sc_hd__nor2_1 _22263_ (.A(_05095_),
    .B(_09148_),
    .Y(_01550_));
 sky130_fd_sc_hd__nor2_1 _22264_ (.A(_05102_),
    .B(_09148_),
    .Y(_01551_));
 sky130_fd_sc_hd__nor2_1 _22265_ (.A(_05112_),
    .B(_09148_),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _22266_ (.A(_05121_),
    .B(_09148_),
    .Y(_01553_));
 sky130_fd_sc_hd__nor2_1 _22267_ (.A(_05128_),
    .B(_09148_),
    .Y(_01554_));
 sky130_fd_sc_hd__nor2_1 _22268_ (.A(_05137_),
    .B(_09148_),
    .Y(_01555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_804 ();
 sky130_fd_sc_hd__nor2_1 _22270_ (.A(_05154_),
    .B(_09148_),
    .Y(_01556_));
 sky130_fd_sc_hd__nor2_1 _22271_ (.A(_04992_),
    .B(_09148_),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2_1 _22272_ (.A(_05167_),
    .B(_09148_),
    .Y(_01558_));
 sky130_fd_sc_hd__nor2_1 _22273_ (.A(_05175_),
    .B(_09148_),
    .Y(_01559_));
 sky130_fd_sc_hd__nor2_1 _22274_ (.A(_05184_),
    .B(_09148_),
    .Y(_01560_));
 sky130_fd_sc_hd__nor2_1 _22275_ (.A(_05196_),
    .B(_09148_),
    .Y(_01561_));
 sky130_fd_sc_hd__nor2_1 _22276_ (.A(_05206_),
    .B(_09148_),
    .Y(_01562_));
 sky130_fd_sc_hd__nor2_1 _22277_ (.A(_05214_),
    .B(_09148_),
    .Y(_01563_));
 sky130_fd_sc_hd__nor2_1 _22278_ (.A(_05224_),
    .B(_09148_),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_1 _22279_ (.A(_05236_),
    .B(_09148_),
    .Y(_01565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_803 ();
 sky130_fd_sc_hd__nor2_1 _22281_ (.A(_05243_),
    .B(_09148_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_1 _22282_ (.A(_05251_),
    .B(_09148_),
    .Y(_01567_));
 sky130_fd_sc_hd__nor2_1 _22283_ (.A(_04995_),
    .B(_09148_),
    .Y(_01568_));
 sky130_fd_sc_hd__nor2_1 _22284_ (.A(_05260_),
    .B(_09148_),
    .Y(_01569_));
 sky130_fd_sc_hd__nor2_1 _22285_ (.A(_05310_),
    .B(_09148_),
    .Y(_01570_));
 sky130_fd_sc_hd__nor2_1 _22286_ (.A(_05003_),
    .B(_09148_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_1 _22287_ (.A(_05012_),
    .B(_09148_),
    .Y(_01572_));
 sky130_fd_sc_hd__nor2_1 _22288_ (.A(_05021_),
    .B(_09148_),
    .Y(_01573_));
 sky130_fd_sc_hd__nor2_1 _22289_ (.A(_05032_),
    .B(_09148_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor2_1 _22290_ (.A(_05039_),
    .B(_09148_),
    .Y(_01575_));
 sky130_fd_sc_hd__nor2_1 _22291_ (.A(_05048_),
    .B(_09148_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _22292_ (.A(_05055_),
    .B(_09148_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand2_8 _22293_ (.A(_09972_),
    .B(_05313_),
    .Y(_09152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_802 ();
 sky130_fd_sc_hd__nor2_1 _22295_ (.A(_05317_),
    .B(_09152_),
    .Y(_01578_));
 sky130_fd_sc_hd__nor2_1 _22296_ (.A(_05388_),
    .B(_09152_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _22297_ (.A(_05402_),
    .B(_09152_),
    .Y(_01580_));
 sky130_fd_sc_hd__nor2_1 _22298_ (.A(_05412_),
    .B(_09152_),
    .Y(_01581_));
 sky130_fd_sc_hd__nor2_1 _22299_ (.A(_05419_),
    .B(_09152_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_1 _22300_ (.A(_05426_),
    .B(_09152_),
    .Y(_01583_));
 sky130_fd_sc_hd__nor2_1 _22301_ (.A(_05438_),
    .B(_09152_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _22302_ (.A(_05447_),
    .B(_09152_),
    .Y(_01585_));
 sky130_fd_sc_hd__nor2_1 _22303_ (.A(_05453_),
    .B(_09152_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor2_1 _22304_ (.A(_05465_),
    .B(_09152_),
    .Y(_01587_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_801 ();
 sky130_fd_sc_hd__nor2_1 _22306_ (.A(_05480_),
    .B(_09152_),
    .Y(_01588_));
 sky130_fd_sc_hd__nor2_1 _22307_ (.A(_05321_),
    .B(_09152_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_1 _22308_ (.A(_05488_),
    .B(_09152_),
    .Y(_01590_));
 sky130_fd_sc_hd__nor2_1 _22309_ (.A(_05498_),
    .B(_09152_),
    .Y(_01591_));
 sky130_fd_sc_hd__nor2_1 _22310_ (.A(_05509_),
    .B(_09152_),
    .Y(_01592_));
 sky130_fd_sc_hd__nor2_1 _22311_ (.A(_05515_),
    .B(_09152_),
    .Y(_01593_));
 sky130_fd_sc_hd__nor2_1 _22312_ (.A(_05523_),
    .B(_09152_),
    .Y(_01594_));
 sky130_fd_sc_hd__nor2_1 _22313_ (.A(_05535_),
    .B(_09152_),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_1 _22314_ (.A(_05542_),
    .B(_09152_),
    .Y(_01596_));
 sky130_fd_sc_hd__nor2_1 _22315_ (.A(_05551_),
    .B(_09152_),
    .Y(_01597_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_800 ();
 sky130_fd_sc_hd__nor2_1 _22317_ (.A(_05559_),
    .B(_09152_),
    .Y(_01598_));
 sky130_fd_sc_hd__nor2_1 _22318_ (.A(_05567_),
    .B(_09152_),
    .Y(_01599_));
 sky130_fd_sc_hd__nor2_1 _22319_ (.A(_05324_),
    .B(_09152_),
    .Y(_01600_));
 sky130_fd_sc_hd__nor2_1 _22320_ (.A(_05573_),
    .B(_09152_),
    .Y(_01601_));
 sky130_fd_sc_hd__nor2_1 _22321_ (.A(_05611_),
    .B(_09152_),
    .Y(_01602_));
 sky130_fd_sc_hd__nor2_1 _22322_ (.A(_05330_),
    .B(_09152_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _22323_ (.A(_05338_),
    .B(_09152_),
    .Y(_01604_));
 sky130_fd_sc_hd__nor2_1 _22324_ (.A(_05347_),
    .B(_09152_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _22325_ (.A(_05354_),
    .B(_09152_),
    .Y(_01606_));
 sky130_fd_sc_hd__nor2_1 _22326_ (.A(_05360_),
    .B(_09152_),
    .Y(_01607_));
 sky130_fd_sc_hd__nor2_1 _22327_ (.A(_05371_),
    .B(_09152_),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_1 _22328_ (.A(_05380_),
    .B(_09152_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_8 _22329_ (.A(_09921_),
    .B(_05614_),
    .Y(_09156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_799 ();
 sky130_fd_sc_hd__nor2_1 _22331_ (.A(_04988_),
    .B(_09156_),
    .Y(_01610_));
 sky130_fd_sc_hd__nor2_1 _22332_ (.A(_05062_),
    .B(_09156_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_1 _22333_ (.A(_05077_),
    .B(_09156_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_1 _22334_ (.A(_05087_),
    .B(_09156_),
    .Y(_01613_));
 sky130_fd_sc_hd__nor2_1 _22335_ (.A(_05095_),
    .B(_09156_),
    .Y(_01614_));
 sky130_fd_sc_hd__nor2_1 _22336_ (.A(_05102_),
    .B(_09156_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_1 _22337_ (.A(_05112_),
    .B(_09156_),
    .Y(_01616_));
 sky130_fd_sc_hd__nor2_1 _22338_ (.A(_05121_),
    .B(_09156_),
    .Y(_01617_));
 sky130_fd_sc_hd__nor2_1 _22339_ (.A(_05128_),
    .B(_09156_),
    .Y(_01618_));
 sky130_fd_sc_hd__nor2_1 _22340_ (.A(_05137_),
    .B(_09156_),
    .Y(_01619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_798 ();
 sky130_fd_sc_hd__nor2_1 _22342_ (.A(_05154_),
    .B(_09156_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _22343_ (.A(_04992_),
    .B(_09156_),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_1 _22344_ (.A(_05167_),
    .B(_09156_),
    .Y(_01622_));
 sky130_fd_sc_hd__nor2_1 _22345_ (.A(_05175_),
    .B(_09156_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_1 _22346_ (.A(_05184_),
    .B(_09156_),
    .Y(_01624_));
 sky130_fd_sc_hd__nor2_1 _22347_ (.A(_05196_),
    .B(_09156_),
    .Y(_01625_));
 sky130_fd_sc_hd__nor2_1 _22348_ (.A(_05206_),
    .B(_09156_),
    .Y(_01626_));
 sky130_fd_sc_hd__nor2_1 _22349_ (.A(_05214_),
    .B(_09156_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _22350_ (.A(_05224_),
    .B(_09156_),
    .Y(_01628_));
 sky130_fd_sc_hd__nor2_1 _22351_ (.A(_05236_),
    .B(_09156_),
    .Y(_01629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_797 ();
 sky130_fd_sc_hd__nor2_1 _22353_ (.A(_05243_),
    .B(_09156_),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_1 _22354_ (.A(_05251_),
    .B(_09156_),
    .Y(_01631_));
 sky130_fd_sc_hd__nor2_1 _22355_ (.A(_04995_),
    .B(_09156_),
    .Y(_01632_));
 sky130_fd_sc_hd__nor2_1 _22356_ (.A(_05260_),
    .B(_09156_),
    .Y(_01633_));
 sky130_fd_sc_hd__nor2_1 _22357_ (.A(_05310_),
    .B(_09156_),
    .Y(_01634_));
 sky130_fd_sc_hd__nor2_1 _22358_ (.A(_05003_),
    .B(_09156_),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_1 _22359_ (.A(_05012_),
    .B(_09156_),
    .Y(_01636_));
 sky130_fd_sc_hd__nor2_1 _22360_ (.A(_05021_),
    .B(_09156_),
    .Y(_01637_));
 sky130_fd_sc_hd__nor2_1 _22361_ (.A(_05032_),
    .B(_09156_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor2_1 _22362_ (.A(_05039_),
    .B(_09156_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_1 _22363_ (.A(_05048_),
    .B(_09156_),
    .Y(_01640_));
 sky130_fd_sc_hd__nor2_1 _22364_ (.A(_05055_),
    .B(_09156_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_8 _22365_ (.A(_09972_),
    .B(_05655_),
    .Y(_09160_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_796 ();
 sky130_fd_sc_hd__nor2_1 _22367_ (.A(_05317_),
    .B(_09160_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor2_1 _22368_ (.A(_05388_),
    .B(_09160_),
    .Y(_01643_));
 sky130_fd_sc_hd__nor2_1 _22369_ (.A(_05402_),
    .B(_09160_),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _22370_ (.A(_05412_),
    .B(_09160_),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_1 _22371_ (.A(_05419_),
    .B(_09160_),
    .Y(_01646_));
 sky130_fd_sc_hd__nor2_1 _22372_ (.A(_05426_),
    .B(_09160_),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_1 _22373_ (.A(_05438_),
    .B(_09160_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_1 _22374_ (.A(_05447_),
    .B(_09160_),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_1 _22375_ (.A(_05453_),
    .B(_09160_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _22376_ (.A(_05465_),
    .B(_09160_),
    .Y(_01651_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_795 ();
 sky130_fd_sc_hd__nor2_1 _22378_ (.A(_05480_),
    .B(_09160_),
    .Y(_01652_));
 sky130_fd_sc_hd__nor2_1 _22379_ (.A(_05321_),
    .B(_09160_),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _22380_ (.A(_05488_),
    .B(_09160_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_1 _22381_ (.A(_05498_),
    .B(_09160_),
    .Y(_01655_));
 sky130_fd_sc_hd__nor2_1 _22382_ (.A(_05509_),
    .B(_09160_),
    .Y(_01656_));
 sky130_fd_sc_hd__nor2_1 _22383_ (.A(_05515_),
    .B(_09160_),
    .Y(_01657_));
 sky130_fd_sc_hd__nor2_1 _22384_ (.A(_05523_),
    .B(_09160_),
    .Y(_01658_));
 sky130_fd_sc_hd__nor2_1 _22385_ (.A(_05535_),
    .B(_09160_),
    .Y(_01659_));
 sky130_fd_sc_hd__nor2_1 _22386_ (.A(_05542_),
    .B(_09160_),
    .Y(_01660_));
 sky130_fd_sc_hd__nor2_1 _22387_ (.A(_05551_),
    .B(_09160_),
    .Y(_01661_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_794 ();
 sky130_fd_sc_hd__nor2_1 _22389_ (.A(_05559_),
    .B(_09160_),
    .Y(_01662_));
 sky130_fd_sc_hd__nor2_1 _22390_ (.A(_05567_),
    .B(_09160_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor2_1 _22391_ (.A(_05324_),
    .B(_09160_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_1 _22392_ (.A(_05573_),
    .B(_09160_),
    .Y(_01665_));
 sky130_fd_sc_hd__nor2_1 _22393_ (.A(_05611_),
    .B(_09160_),
    .Y(_01666_));
 sky130_fd_sc_hd__nor2_1 _22394_ (.A(_05330_),
    .B(_09160_),
    .Y(_01667_));
 sky130_fd_sc_hd__nor2_1 _22395_ (.A(_05338_),
    .B(_09160_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _22396_ (.A(_05347_),
    .B(_09160_),
    .Y(_01669_));
 sky130_fd_sc_hd__nor2_1 _22397_ (.A(_05354_),
    .B(_09160_),
    .Y(_01670_));
 sky130_fd_sc_hd__nor2_1 _22398_ (.A(_05360_),
    .B(_09160_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_1 _22399_ (.A(_05371_),
    .B(_09160_),
    .Y(_01672_));
 sky130_fd_sc_hd__nor2_1 _22400_ (.A(_05380_),
    .B(_09160_),
    .Y(_01673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_793 ();
 sky130_fd_sc_hd__nand2_8 _22402_ (.A(_09921_),
    .B(_05696_),
    .Y(_09165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_792 ();
 sky130_fd_sc_hd__nor2_1 _22404_ (.A(_04988_),
    .B(_09165_),
    .Y(_01674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_791 ();
 sky130_fd_sc_hd__nor2_1 _22406_ (.A(_05062_),
    .B(_09165_),
    .Y(_01675_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_790 ();
 sky130_fd_sc_hd__nor2_1 _22408_ (.A(_05077_),
    .B(_09165_),
    .Y(_01676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_789 ();
 sky130_fd_sc_hd__nor2_1 _22410_ (.A(_05087_),
    .B(_09165_),
    .Y(_01677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_788 ();
 sky130_fd_sc_hd__nor2_1 _22412_ (.A(_05095_),
    .B(_09165_),
    .Y(_01678_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_787 ();
 sky130_fd_sc_hd__nor2_1 _22414_ (.A(_05102_),
    .B(_09165_),
    .Y(_01679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_786 ();
 sky130_fd_sc_hd__nor2_1 _22416_ (.A(_05112_),
    .B(_09165_),
    .Y(_01680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_785 ();
 sky130_fd_sc_hd__nor2_1 _22418_ (.A(_05121_),
    .B(_09165_),
    .Y(_01681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_784 ();
 sky130_fd_sc_hd__nor2_1 _22420_ (.A(_05128_),
    .B(_09165_),
    .Y(_01682_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_783 ();
 sky130_fd_sc_hd__nor2_1 _22422_ (.A(_05137_),
    .B(_09165_),
    .Y(_01683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_781 ();
 sky130_fd_sc_hd__nor2_1 _22425_ (.A(_05154_),
    .B(_09165_),
    .Y(_01684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_780 ();
 sky130_fd_sc_hd__nor2_1 _22427_ (.A(_04992_),
    .B(_09165_),
    .Y(_01685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_779 ();
 sky130_fd_sc_hd__nor2_1 _22429_ (.A(_05167_),
    .B(_09165_),
    .Y(_01686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_778 ();
 sky130_fd_sc_hd__nor2_1 _22431_ (.A(_05175_),
    .B(_09165_),
    .Y(_01687_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_777 ();
 sky130_fd_sc_hd__nor2_1 _22433_ (.A(_05184_),
    .B(_09165_),
    .Y(_01688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_776 ();
 sky130_fd_sc_hd__nor2_1 _22435_ (.A(_05196_),
    .B(_09165_),
    .Y(_01689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_775 ();
 sky130_fd_sc_hd__nor2_1 _22437_ (.A(_05206_),
    .B(_09165_),
    .Y(_01690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_774 ();
 sky130_fd_sc_hd__nor2_1 _22439_ (.A(_05214_),
    .B(_09165_),
    .Y(_01691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_773 ();
 sky130_fd_sc_hd__nor2_1 _22441_ (.A(_05224_),
    .B(_09165_),
    .Y(_01692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_772 ();
 sky130_fd_sc_hd__nor2_1 _22443_ (.A(_05236_),
    .B(_09165_),
    .Y(_01693_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_770 ();
 sky130_fd_sc_hd__nor2_1 _22446_ (.A(_05243_),
    .B(_09165_),
    .Y(_01694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_769 ();
 sky130_fd_sc_hd__nor2_1 _22448_ (.A(_05251_),
    .B(_09165_),
    .Y(_01695_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_768 ();
 sky130_fd_sc_hd__nor2_1 _22450_ (.A(_04995_),
    .B(_09165_),
    .Y(_01696_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_767 ();
 sky130_fd_sc_hd__nor2_1 _22452_ (.A(_05260_),
    .B(_09165_),
    .Y(_01697_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_766 ();
 sky130_fd_sc_hd__nor2_1 _22454_ (.A(_05310_),
    .B(_09165_),
    .Y(_01698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_765 ();
 sky130_fd_sc_hd__nor2_1 _22456_ (.A(_05003_),
    .B(_09165_),
    .Y(_01699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_764 ();
 sky130_fd_sc_hd__nor2_1 _22458_ (.A(_05012_),
    .B(_09165_),
    .Y(_01700_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_763 ();
 sky130_fd_sc_hd__nor2_1 _22460_ (.A(_05021_),
    .B(_09165_),
    .Y(_01701_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_762 ();
 sky130_fd_sc_hd__nor2_1 _22462_ (.A(_05032_),
    .B(_09165_),
    .Y(_01702_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_761 ();
 sky130_fd_sc_hd__nor2_1 _22464_ (.A(_05039_),
    .B(_09165_),
    .Y(_01703_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_760 ();
 sky130_fd_sc_hd__nor2_1 _22466_ (.A(_05048_),
    .B(_09165_),
    .Y(_01704_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_759 ();
 sky130_fd_sc_hd__nor2_1 _22468_ (.A(_05055_),
    .B(_09165_),
    .Y(_01705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_758 ();
 sky130_fd_sc_hd__nand2_8 _22470_ (.A(_09972_),
    .B(_05737_),
    .Y(_09201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_757 ();
 sky130_fd_sc_hd__nor2_1 _22472_ (.A(_05317_),
    .B(_09201_),
    .Y(_01706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_756 ();
 sky130_fd_sc_hd__nor2_1 _22474_ (.A(_05388_),
    .B(_09201_),
    .Y(_01707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_755 ();
 sky130_fd_sc_hd__nor2_1 _22476_ (.A(_05402_),
    .B(_09201_),
    .Y(_01708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_754 ();
 sky130_fd_sc_hd__nor2_1 _22478_ (.A(_05412_),
    .B(_09201_),
    .Y(_01709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_753 ();
 sky130_fd_sc_hd__nor2_1 _22480_ (.A(_05419_),
    .B(_09201_),
    .Y(_01710_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_752 ();
 sky130_fd_sc_hd__nor2_1 _22482_ (.A(_05426_),
    .B(_09201_),
    .Y(_01711_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_751 ();
 sky130_fd_sc_hd__nor2_1 _22484_ (.A(_05438_),
    .B(_09201_),
    .Y(_01712_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_750 ();
 sky130_fd_sc_hd__nor2_1 _22486_ (.A(_05447_),
    .B(_09201_),
    .Y(_01713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_749 ();
 sky130_fd_sc_hd__nor2_1 _22488_ (.A(_05453_),
    .B(_09201_),
    .Y(_01714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_748 ();
 sky130_fd_sc_hd__nor2_1 _22490_ (.A(_05465_),
    .B(_09201_),
    .Y(_01715_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_746 ();
 sky130_fd_sc_hd__nor2_1 _22493_ (.A(_05480_),
    .B(_09201_),
    .Y(_01716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_745 ();
 sky130_fd_sc_hd__nor2_1 _22495_ (.A(_05321_),
    .B(_09201_),
    .Y(_01717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_744 ();
 sky130_fd_sc_hd__nor2_1 _22497_ (.A(_05488_),
    .B(_09201_),
    .Y(_01718_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_743 ();
 sky130_fd_sc_hd__nor2_1 _22499_ (.A(_05498_),
    .B(_09201_),
    .Y(_01719_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_742 ();
 sky130_fd_sc_hd__nor2_1 _22501_ (.A(_05509_),
    .B(_09201_),
    .Y(_01720_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_741 ();
 sky130_fd_sc_hd__nor2_1 _22503_ (.A(_05515_),
    .B(_09201_),
    .Y(_01721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_740 ();
 sky130_fd_sc_hd__nor2_1 _22505_ (.A(_05523_),
    .B(_09201_),
    .Y(_01722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_739 ();
 sky130_fd_sc_hd__nor2_1 _22507_ (.A(_05535_),
    .B(_09201_),
    .Y(_01723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_738 ();
 sky130_fd_sc_hd__nor2_1 _22509_ (.A(_05542_),
    .B(_09201_),
    .Y(_01724_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_737 ();
 sky130_fd_sc_hd__nor2_1 _22511_ (.A(_05551_),
    .B(_09201_),
    .Y(_01725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_735 ();
 sky130_fd_sc_hd__nor2_1 _22514_ (.A(_05559_),
    .B(_09201_),
    .Y(_01726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_734 ();
 sky130_fd_sc_hd__nor2_1 _22516_ (.A(_05567_),
    .B(_09201_),
    .Y(_01727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_733 ();
 sky130_fd_sc_hd__nor2_1 _22518_ (.A(_05324_),
    .B(_09201_),
    .Y(_01728_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_732 ();
 sky130_fd_sc_hd__nor2_1 _22520_ (.A(_05573_),
    .B(_09201_),
    .Y(_01729_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_731 ();
 sky130_fd_sc_hd__nor2_1 _22522_ (.A(_05611_),
    .B(_09201_),
    .Y(_01730_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_730 ();
 sky130_fd_sc_hd__nor2_1 _22524_ (.A(_05330_),
    .B(_09201_),
    .Y(_01731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_729 ();
 sky130_fd_sc_hd__nor2_1 _22526_ (.A(_05338_),
    .B(_09201_),
    .Y(_01732_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_728 ();
 sky130_fd_sc_hd__nor2_1 _22528_ (.A(_05347_),
    .B(_09201_),
    .Y(_01733_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_727 ();
 sky130_fd_sc_hd__nor2_1 _22530_ (.A(_05354_),
    .B(_09201_),
    .Y(_01734_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_726 ();
 sky130_fd_sc_hd__nor2_1 _22532_ (.A(_05360_),
    .B(_09201_),
    .Y(_01735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_725 ();
 sky130_fd_sc_hd__nor2_1 _22534_ (.A(_05371_),
    .B(_09201_),
    .Y(_01736_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_724 ();
 sky130_fd_sc_hd__nor2_1 _22536_ (.A(_05380_),
    .B(_09201_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_8 _22537_ (.A(_09921_),
    .B(_05778_),
    .Y(_09236_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_723 ();
 sky130_fd_sc_hd__nor2_1 _22539_ (.A(_04988_),
    .B(_09236_),
    .Y(_01738_));
 sky130_fd_sc_hd__nor2_1 _22540_ (.A(_05062_),
    .B(_09236_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _22541_ (.A(_05077_),
    .B(_09236_),
    .Y(_01740_));
 sky130_fd_sc_hd__nor2_1 _22542_ (.A(_05087_),
    .B(_09236_),
    .Y(_01741_));
 sky130_fd_sc_hd__nor2_1 _22543_ (.A(_05095_),
    .B(_09236_),
    .Y(_01742_));
 sky130_fd_sc_hd__nor2_1 _22544_ (.A(_05102_),
    .B(_09236_),
    .Y(_01743_));
 sky130_fd_sc_hd__nor2_1 _22545_ (.A(_05112_),
    .B(_09236_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _22546_ (.A(_05121_),
    .B(_09236_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor2_1 _22547_ (.A(_05128_),
    .B(_09236_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _22548_ (.A(_05137_),
    .B(_09236_),
    .Y(_01747_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_722 ();
 sky130_fd_sc_hd__nor2_1 _22550_ (.A(_05154_),
    .B(_09236_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _22551_ (.A(_04992_),
    .B(_09236_),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_1 _22552_ (.A(_05167_),
    .B(_09236_),
    .Y(_01750_));
 sky130_fd_sc_hd__nor2_1 _22553_ (.A(_05175_),
    .B(_09236_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor2_1 _22554_ (.A(_05184_),
    .B(_09236_),
    .Y(_01752_));
 sky130_fd_sc_hd__nor2_1 _22555_ (.A(_05196_),
    .B(_09236_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_1 _22556_ (.A(_05206_),
    .B(_09236_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _22557_ (.A(_05214_),
    .B(_09236_),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_1 _22558_ (.A(_05224_),
    .B(_09236_),
    .Y(_01756_));
 sky130_fd_sc_hd__nor2_1 _22559_ (.A(_05236_),
    .B(_09236_),
    .Y(_01757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_721 ();
 sky130_fd_sc_hd__nor2_1 _22561_ (.A(_05243_),
    .B(_09236_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _22562_ (.A(_05251_),
    .B(_09236_),
    .Y(_01759_));
 sky130_fd_sc_hd__nor2_1 _22563_ (.A(_04995_),
    .B(_09236_),
    .Y(_01760_));
 sky130_fd_sc_hd__nor2_1 _22564_ (.A(_05260_),
    .B(_09236_),
    .Y(_01761_));
 sky130_fd_sc_hd__nor2_1 _22565_ (.A(_05310_),
    .B(_09236_),
    .Y(_01762_));
 sky130_fd_sc_hd__nor2_1 _22566_ (.A(_05003_),
    .B(_09236_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _22567_ (.A(_05012_),
    .B(_09236_),
    .Y(_01764_));
 sky130_fd_sc_hd__nor2_1 _22568_ (.A(_05021_),
    .B(_09236_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_1 _22569_ (.A(_05032_),
    .B(_09236_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor2_1 _22570_ (.A(_05039_),
    .B(_09236_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _22571_ (.A(_05048_),
    .B(_09236_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _22572_ (.A(_05055_),
    .B(_09236_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand3_4 _22573_ (.A(_13709_),
    .B(\count_2[5] ),
    .C(_05820_),
    .Y(_09240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_720 ();
 sky130_fd_sc_hd__nor2_1 _22575_ (.A(_05317_),
    .B(_09240_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor2_1 _22576_ (.A(_05388_),
    .B(_09240_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _22577_ (.A(_05402_),
    .B(_09240_),
    .Y(_01772_));
 sky130_fd_sc_hd__nor2_1 _22578_ (.A(_05412_),
    .B(_09240_),
    .Y(_01773_));
 sky130_fd_sc_hd__nor2_1 _22579_ (.A(_05419_),
    .B(_09240_),
    .Y(_01774_));
 sky130_fd_sc_hd__nor2_1 _22580_ (.A(_05426_),
    .B(_09240_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _22581_ (.A(_05438_),
    .B(_09240_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor2_1 _22582_ (.A(_05447_),
    .B(_09240_),
    .Y(_01777_));
 sky130_fd_sc_hd__nor2_1 _22583_ (.A(_05453_),
    .B(_09240_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _22584_ (.A(_05465_),
    .B(_09240_),
    .Y(_01779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_719 ();
 sky130_fd_sc_hd__nor2_1 _22586_ (.A(_05480_),
    .B(_09240_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _22587_ (.A(_05321_),
    .B(_09240_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _22588_ (.A(_05488_),
    .B(_09240_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor2_1 _22589_ (.A(_05498_),
    .B(_09240_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_1 _22590_ (.A(_05509_),
    .B(_09240_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _22591_ (.A(_05515_),
    .B(_09240_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _22592_ (.A(_05523_),
    .B(_09240_),
    .Y(_01786_));
 sky130_fd_sc_hd__nor2_1 _22593_ (.A(_05535_),
    .B(_09240_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _22594_ (.A(_05542_),
    .B(_09240_),
    .Y(_01788_));
 sky130_fd_sc_hd__nor2_1 _22595_ (.A(_05551_),
    .B(_09240_),
    .Y(_01789_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_718 ();
 sky130_fd_sc_hd__nor2_1 _22597_ (.A(_05559_),
    .B(_09240_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor2_1 _22598_ (.A(_05567_),
    .B(_09240_),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _22599_ (.A(_05324_),
    .B(_09240_),
    .Y(_01792_));
 sky130_fd_sc_hd__nor2_1 _22600_ (.A(_05573_),
    .B(_09240_),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _22601_ (.A(_05611_),
    .B(_09240_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _22602_ (.A(_05330_),
    .B(_09240_),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_1 _22603_ (.A(_05338_),
    .B(_09240_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _22604_ (.A(_05347_),
    .B(_09240_),
    .Y(_01797_));
 sky130_fd_sc_hd__nor2_1 _22605_ (.A(_05354_),
    .B(_09240_),
    .Y(_01798_));
 sky130_fd_sc_hd__nor2_1 _22606_ (.A(_05360_),
    .B(_09240_),
    .Y(_01799_));
 sky130_fd_sc_hd__nor2_1 _22607_ (.A(_05371_),
    .B(_09240_),
    .Y(_01800_));
 sky130_fd_sc_hd__nor2_1 _22608_ (.A(_05380_),
    .B(_09240_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_8 _22609_ (.A(_09926_),
    .B(_04982_),
    .Y(_09244_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_717 ();
 sky130_fd_sc_hd__nor2_1 _22611_ (.A(_04988_),
    .B(_09244_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _22612_ (.A(_05062_),
    .B(_09244_),
    .Y(_01803_));
 sky130_fd_sc_hd__nor2_1 _22613_ (.A(_05077_),
    .B(_09244_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _22614_ (.A(_05087_),
    .B(_09244_),
    .Y(_01805_));
 sky130_fd_sc_hd__nor2_1 _22615_ (.A(_05095_),
    .B(_09244_),
    .Y(_01806_));
 sky130_fd_sc_hd__nor2_1 _22616_ (.A(_05102_),
    .B(_09244_),
    .Y(_01807_));
 sky130_fd_sc_hd__nor2_1 _22617_ (.A(_05112_),
    .B(_09244_),
    .Y(_01808_));
 sky130_fd_sc_hd__nor2_1 _22618_ (.A(_05121_),
    .B(_09244_),
    .Y(_01809_));
 sky130_fd_sc_hd__nor2_1 _22619_ (.A(_05128_),
    .B(_09244_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _22620_ (.A(_05137_),
    .B(_09244_),
    .Y(_01811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_716 ();
 sky130_fd_sc_hd__nor2_1 _22622_ (.A(_05154_),
    .B(_09244_),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_1 _22623_ (.A(_04992_),
    .B(_09244_),
    .Y(_01813_));
 sky130_fd_sc_hd__nor2_1 _22624_ (.A(_05167_),
    .B(_09244_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_1 _22625_ (.A(_05175_),
    .B(_09244_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _22626_ (.A(_05184_),
    .B(_09244_),
    .Y(_01816_));
 sky130_fd_sc_hd__nor2_1 _22627_ (.A(_05196_),
    .B(_09244_),
    .Y(_01817_));
 sky130_fd_sc_hd__nor2_1 _22628_ (.A(_05206_),
    .B(_09244_),
    .Y(_01818_));
 sky130_fd_sc_hd__nor2_1 _22629_ (.A(_05214_),
    .B(_09244_),
    .Y(_01819_));
 sky130_fd_sc_hd__nor2_1 _22630_ (.A(_05224_),
    .B(_09244_),
    .Y(_01820_));
 sky130_fd_sc_hd__nor2_1 _22631_ (.A(_05236_),
    .B(_09244_),
    .Y(_01821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_715 ();
 sky130_fd_sc_hd__nor2_1 _22633_ (.A(_05243_),
    .B(_09244_),
    .Y(_01822_));
 sky130_fd_sc_hd__nor2_1 _22634_ (.A(_05251_),
    .B(_09244_),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_1 _22635_ (.A(_04995_),
    .B(_09244_),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _22636_ (.A(_05260_),
    .B(_09244_),
    .Y(_01825_));
 sky130_fd_sc_hd__nor2_1 _22637_ (.A(_05310_),
    .B(_09244_),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _22638_ (.A(_05003_),
    .B(_09244_),
    .Y(_01827_));
 sky130_fd_sc_hd__nor2_1 _22639_ (.A(_05012_),
    .B(_09244_),
    .Y(_01828_));
 sky130_fd_sc_hd__nor2_1 _22640_ (.A(_05021_),
    .B(_09244_),
    .Y(_01829_));
 sky130_fd_sc_hd__nor2_1 _22641_ (.A(_05032_),
    .B(_09244_),
    .Y(_01830_));
 sky130_fd_sc_hd__nor2_1 _22642_ (.A(_05039_),
    .B(_09244_),
    .Y(_01831_));
 sky130_fd_sc_hd__nor2_1 _22643_ (.A(_05048_),
    .B(_09244_),
    .Y(_01832_));
 sky130_fd_sc_hd__nor2_1 _22644_ (.A(_05055_),
    .B(_09244_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_8 _22645_ (.A(_09979_),
    .B(_05313_),
    .Y(_09248_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_714 ();
 sky130_fd_sc_hd__nor2_1 _22647_ (.A(_05317_),
    .B(_09248_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _22648_ (.A(_05388_),
    .B(_09248_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor2_1 _22649_ (.A(_05402_),
    .B(_09248_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _22650_ (.A(_05412_),
    .B(_09248_),
    .Y(_01837_));
 sky130_fd_sc_hd__nor2_1 _22651_ (.A(_05419_),
    .B(_09248_),
    .Y(_01838_));
 sky130_fd_sc_hd__nor2_1 _22652_ (.A(_05426_),
    .B(_09248_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _22653_ (.A(_05438_),
    .B(_09248_),
    .Y(_01840_));
 sky130_fd_sc_hd__nor2_1 _22654_ (.A(_05447_),
    .B(_09248_),
    .Y(_01841_));
 sky130_fd_sc_hd__nor2_1 _22655_ (.A(_05453_),
    .B(_09248_),
    .Y(_01842_));
 sky130_fd_sc_hd__nor2_1 _22656_ (.A(_05465_),
    .B(_09248_),
    .Y(_01843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_713 ();
 sky130_fd_sc_hd__nor2_1 _22658_ (.A(_05480_),
    .B(_09248_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _22659_ (.A(_05321_),
    .B(_09248_),
    .Y(_01845_));
 sky130_fd_sc_hd__nor2_1 _22660_ (.A(_05488_),
    .B(_09248_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_1 _22661_ (.A(_05498_),
    .B(_09248_),
    .Y(_01847_));
 sky130_fd_sc_hd__nor2_1 _22662_ (.A(_05509_),
    .B(_09248_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_1 _22663_ (.A(_05515_),
    .B(_09248_),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _22664_ (.A(_05523_),
    .B(_09248_),
    .Y(_01850_));
 sky130_fd_sc_hd__nor2_1 _22665_ (.A(_05535_),
    .B(_09248_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor2_1 _22666_ (.A(_05542_),
    .B(_09248_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _22667_ (.A(_05551_),
    .B(_09248_),
    .Y(_01853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_712 ();
 sky130_fd_sc_hd__nor2_1 _22669_ (.A(_05559_),
    .B(_09248_),
    .Y(_01854_));
 sky130_fd_sc_hd__nor2_1 _22670_ (.A(_05567_),
    .B(_09248_),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_1 _22671_ (.A(_05324_),
    .B(_09248_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _22672_ (.A(_05573_),
    .B(_09248_),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _22673_ (.A(_05611_),
    .B(_09248_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _22674_ (.A(_05330_),
    .B(_09248_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _22675_ (.A(_05338_),
    .B(_09248_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor2_1 _22676_ (.A(_05347_),
    .B(_09248_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _22677_ (.A(_05354_),
    .B(_09248_),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_1 _22678_ (.A(_05360_),
    .B(_09248_),
    .Y(_01863_));
 sky130_fd_sc_hd__nor2_1 _22679_ (.A(_05371_),
    .B(_09248_),
    .Y(_01864_));
 sky130_fd_sc_hd__nor2_1 _22680_ (.A(_05380_),
    .B(_09248_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_8 _22681_ (.A(_09926_),
    .B(_05614_),
    .Y(_09252_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_711 ();
 sky130_fd_sc_hd__nor2_1 _22683_ (.A(_04988_),
    .B(_09252_),
    .Y(_01866_));
 sky130_fd_sc_hd__nor2_1 _22684_ (.A(_05062_),
    .B(_09252_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor2_1 _22685_ (.A(_05077_),
    .B(_09252_),
    .Y(_01868_));
 sky130_fd_sc_hd__nor2_1 _22686_ (.A(_05087_),
    .B(_09252_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _22687_ (.A(_05095_),
    .B(_09252_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _22688_ (.A(_05102_),
    .B(_09252_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _22689_ (.A(_05112_),
    .B(_09252_),
    .Y(_01872_));
 sky130_fd_sc_hd__nor2_1 _22690_ (.A(_05121_),
    .B(_09252_),
    .Y(_01873_));
 sky130_fd_sc_hd__nor2_1 _22691_ (.A(_05128_),
    .B(_09252_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _22692_ (.A(_05137_),
    .B(_09252_),
    .Y(_01875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_710 ();
 sky130_fd_sc_hd__nor2_1 _22694_ (.A(_05154_),
    .B(_09252_),
    .Y(_01876_));
 sky130_fd_sc_hd__nor2_1 _22695_ (.A(_04992_),
    .B(_09252_),
    .Y(_01877_));
 sky130_fd_sc_hd__nor2_1 _22696_ (.A(_05167_),
    .B(_09252_),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _22697_ (.A(_05175_),
    .B(_09252_),
    .Y(_01879_));
 sky130_fd_sc_hd__nor2_1 _22698_ (.A(_05184_),
    .B(_09252_),
    .Y(_01880_));
 sky130_fd_sc_hd__nor2_1 _22699_ (.A(_05196_),
    .B(_09252_),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_1 _22700_ (.A(_05206_),
    .B(_09252_),
    .Y(_01882_));
 sky130_fd_sc_hd__nor2_1 _22701_ (.A(_05214_),
    .B(_09252_),
    .Y(_01883_));
 sky130_fd_sc_hd__nor2_1 _22702_ (.A(_05224_),
    .B(_09252_),
    .Y(_01884_));
 sky130_fd_sc_hd__nor2_1 _22703_ (.A(_05236_),
    .B(_09252_),
    .Y(_01885_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_709 ();
 sky130_fd_sc_hd__nor2_1 _22705_ (.A(_05243_),
    .B(_09252_),
    .Y(_01886_));
 sky130_fd_sc_hd__nor2_1 _22706_ (.A(_05251_),
    .B(_09252_),
    .Y(_01887_));
 sky130_fd_sc_hd__nor2_1 _22707_ (.A(_04995_),
    .B(_09252_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor2_1 _22708_ (.A(_05260_),
    .B(_09252_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor2_1 _22709_ (.A(_05310_),
    .B(_09252_),
    .Y(_01890_));
 sky130_fd_sc_hd__nor2_1 _22710_ (.A(_05003_),
    .B(_09252_),
    .Y(_01891_));
 sky130_fd_sc_hd__nor2_1 _22711_ (.A(_05012_),
    .B(_09252_),
    .Y(_01892_));
 sky130_fd_sc_hd__nor2_1 _22712_ (.A(_05021_),
    .B(_09252_),
    .Y(_01893_));
 sky130_fd_sc_hd__nor2_1 _22713_ (.A(_05032_),
    .B(_09252_),
    .Y(_01894_));
 sky130_fd_sc_hd__nor2_1 _22714_ (.A(_05039_),
    .B(_09252_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _22715_ (.A(_05048_),
    .B(_09252_),
    .Y(_01896_));
 sky130_fd_sc_hd__nor2_1 _22716_ (.A(_05055_),
    .B(_09252_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_8 _22717_ (.A(_09979_),
    .B(_05655_),
    .Y(_09256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_708 ();
 sky130_fd_sc_hd__nor2_1 _22719_ (.A(_05317_),
    .B(_09256_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _22720_ (.A(_05388_),
    .B(_09256_),
    .Y(_01899_));
 sky130_fd_sc_hd__nor2_1 _22721_ (.A(_05402_),
    .B(_09256_),
    .Y(_01900_));
 sky130_fd_sc_hd__nor2_1 _22722_ (.A(_05412_),
    .B(_09256_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _22723_ (.A(_05419_),
    .B(_09256_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _22724_ (.A(_05426_),
    .B(_09256_),
    .Y(_01903_));
 sky130_fd_sc_hd__nor2_1 _22725_ (.A(_05438_),
    .B(_09256_),
    .Y(_01904_));
 sky130_fd_sc_hd__nor2_1 _22726_ (.A(_05447_),
    .B(_09256_),
    .Y(_01905_));
 sky130_fd_sc_hd__nor2_1 _22727_ (.A(_05453_),
    .B(_09256_),
    .Y(_01906_));
 sky130_fd_sc_hd__nor2_1 _22728_ (.A(_05465_),
    .B(_09256_),
    .Y(_01907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_707 ();
 sky130_fd_sc_hd__nor2_1 _22730_ (.A(_05480_),
    .B(_09256_),
    .Y(_01908_));
 sky130_fd_sc_hd__nor2_1 _22731_ (.A(_05321_),
    .B(_09256_),
    .Y(_01909_));
 sky130_fd_sc_hd__nor2_1 _22732_ (.A(_05488_),
    .B(_09256_),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _22733_ (.A(_05498_),
    .B(_09256_),
    .Y(_01911_));
 sky130_fd_sc_hd__nor2_1 _22734_ (.A(_05509_),
    .B(_09256_),
    .Y(_01912_));
 sky130_fd_sc_hd__nor2_1 _22735_ (.A(_05515_),
    .B(_09256_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _22736_ (.A(_05523_),
    .B(_09256_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _22737_ (.A(_05535_),
    .B(_09256_),
    .Y(_01915_));
 sky130_fd_sc_hd__nor2_1 _22738_ (.A(_05542_),
    .B(_09256_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _22739_ (.A(_05551_),
    .B(_09256_),
    .Y(_01917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_706 ();
 sky130_fd_sc_hd__nor2_1 _22741_ (.A(_05559_),
    .B(_09256_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _22742_ (.A(_05567_),
    .B(_09256_),
    .Y(_01919_));
 sky130_fd_sc_hd__nor2_1 _22743_ (.A(_05324_),
    .B(_09256_),
    .Y(_01920_));
 sky130_fd_sc_hd__nor2_1 _22744_ (.A(_05573_),
    .B(_09256_),
    .Y(_01921_));
 sky130_fd_sc_hd__nor2_1 _22745_ (.A(_05611_),
    .B(_09256_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _22746_ (.A(_05330_),
    .B(_09256_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_1 _22747_ (.A(_05338_),
    .B(_09256_),
    .Y(_01924_));
 sky130_fd_sc_hd__nor2_1 _22748_ (.A(_05347_),
    .B(_09256_),
    .Y(_01925_));
 sky130_fd_sc_hd__nor2_1 _22749_ (.A(_05354_),
    .B(_09256_),
    .Y(_01926_));
 sky130_fd_sc_hd__nor2_1 _22750_ (.A(_05360_),
    .B(_09256_),
    .Y(_01927_));
 sky130_fd_sc_hd__nor2_1 _22751_ (.A(_05371_),
    .B(_09256_),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _22752_ (.A(_05380_),
    .B(_09256_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_8 _22753_ (.A(_09926_),
    .B(_05696_),
    .Y(_09260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_705 ();
 sky130_fd_sc_hd__nor2_1 _22755_ (.A(_04988_),
    .B(_09260_),
    .Y(_01930_));
 sky130_fd_sc_hd__nor2_1 _22756_ (.A(_05062_),
    .B(_09260_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _22757_ (.A(_05077_),
    .B(_09260_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_1 _22758_ (.A(_05087_),
    .B(_09260_),
    .Y(_01933_));
 sky130_fd_sc_hd__nor2_1 _22759_ (.A(_05095_),
    .B(_09260_),
    .Y(_01934_));
 sky130_fd_sc_hd__nor2_1 _22760_ (.A(_05102_),
    .B(_09260_),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_1 _22761_ (.A(_05112_),
    .B(_09260_),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _22762_ (.A(_05121_),
    .B(_09260_),
    .Y(_01937_));
 sky130_fd_sc_hd__nor2_1 _22763_ (.A(_05128_),
    .B(_09260_),
    .Y(_01938_));
 sky130_fd_sc_hd__nor2_1 _22764_ (.A(_05137_),
    .B(_09260_),
    .Y(_01939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_704 ();
 sky130_fd_sc_hd__nor2_1 _22766_ (.A(_05154_),
    .B(_09260_),
    .Y(_01940_));
 sky130_fd_sc_hd__nor2_1 _22767_ (.A(_04992_),
    .B(_09260_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor2_1 _22768_ (.A(_05167_),
    .B(_09260_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_1 _22769_ (.A(_05175_),
    .B(_09260_),
    .Y(_01943_));
 sky130_fd_sc_hd__nor2_1 _22770_ (.A(_05184_),
    .B(_09260_),
    .Y(_01944_));
 sky130_fd_sc_hd__nor2_1 _22771_ (.A(_05196_),
    .B(_09260_),
    .Y(_01945_));
 sky130_fd_sc_hd__nor2_1 _22772_ (.A(_05206_),
    .B(_09260_),
    .Y(_01946_));
 sky130_fd_sc_hd__nor2_1 _22773_ (.A(_05214_),
    .B(_09260_),
    .Y(_01947_));
 sky130_fd_sc_hd__nor2_1 _22774_ (.A(_05224_),
    .B(_09260_),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_1 _22775_ (.A(_05236_),
    .B(_09260_),
    .Y(_01949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_703 ();
 sky130_fd_sc_hd__nor2_1 _22777_ (.A(_05243_),
    .B(_09260_),
    .Y(_01950_));
 sky130_fd_sc_hd__nor2_1 _22778_ (.A(_05251_),
    .B(_09260_),
    .Y(_01951_));
 sky130_fd_sc_hd__nor2_1 _22779_ (.A(_04995_),
    .B(_09260_),
    .Y(_01952_));
 sky130_fd_sc_hd__nor2_1 _22780_ (.A(_05260_),
    .B(_09260_),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _22781_ (.A(_05310_),
    .B(_09260_),
    .Y(_01954_));
 sky130_fd_sc_hd__nor2_1 _22782_ (.A(_05003_),
    .B(_09260_),
    .Y(_01955_));
 sky130_fd_sc_hd__nor2_1 _22783_ (.A(_05012_),
    .B(_09260_),
    .Y(_01956_));
 sky130_fd_sc_hd__nor2_1 _22784_ (.A(_05021_),
    .B(_09260_),
    .Y(_01957_));
 sky130_fd_sc_hd__nor2_1 _22785_ (.A(_05032_),
    .B(_09260_),
    .Y(_01958_));
 sky130_fd_sc_hd__nor2_1 _22786_ (.A(_05039_),
    .B(_09260_),
    .Y(_01959_));
 sky130_fd_sc_hd__nor2_1 _22787_ (.A(_05048_),
    .B(_09260_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2_1 _22788_ (.A(_05055_),
    .B(_09260_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_8 _22789_ (.A(_09979_),
    .B(_05737_),
    .Y(_09264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_702 ();
 sky130_fd_sc_hd__nor2_1 _22791_ (.A(_05317_),
    .B(_09264_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _22792_ (.A(_05388_),
    .B(_09264_),
    .Y(_01963_));
 sky130_fd_sc_hd__nor2_1 _22793_ (.A(_05402_),
    .B(_09264_),
    .Y(_01964_));
 sky130_fd_sc_hd__nor2_1 _22794_ (.A(_05412_),
    .B(_09264_),
    .Y(_01965_));
 sky130_fd_sc_hd__nor2_1 _22795_ (.A(_05419_),
    .B(_09264_),
    .Y(_01966_));
 sky130_fd_sc_hd__nor2_1 _22796_ (.A(_05426_),
    .B(_09264_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _22797_ (.A(_05438_),
    .B(_09264_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor2_1 _22798_ (.A(_05447_),
    .B(_09264_),
    .Y(_01969_));
 sky130_fd_sc_hd__nor2_1 _22799_ (.A(_05453_),
    .B(_09264_),
    .Y(_01970_));
 sky130_fd_sc_hd__nor2_1 _22800_ (.A(_05465_),
    .B(_09264_),
    .Y(_01971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_701 ();
 sky130_fd_sc_hd__nor2_1 _22802_ (.A(_05480_),
    .B(_09264_),
    .Y(_01972_));
 sky130_fd_sc_hd__nor2_1 _22803_ (.A(_05321_),
    .B(_09264_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_1 _22804_ (.A(_05488_),
    .B(_09264_),
    .Y(_01974_));
 sky130_fd_sc_hd__nor2_1 _22805_ (.A(_05498_),
    .B(_09264_),
    .Y(_01975_));
 sky130_fd_sc_hd__nor2_1 _22806_ (.A(_05509_),
    .B(_09264_),
    .Y(_01976_));
 sky130_fd_sc_hd__nor2_1 _22807_ (.A(_05515_),
    .B(_09264_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_1 _22808_ (.A(_05523_),
    .B(_09264_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _22809_ (.A(_05535_),
    .B(_09264_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _22810_ (.A(_05542_),
    .B(_09264_),
    .Y(_01980_));
 sky130_fd_sc_hd__nor2_1 _22811_ (.A(_05551_),
    .B(_09264_),
    .Y(_01981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_700 ();
 sky130_fd_sc_hd__nor2_1 _22813_ (.A(_05559_),
    .B(_09264_),
    .Y(_01982_));
 sky130_fd_sc_hd__nor2_1 _22814_ (.A(_05567_),
    .B(_09264_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _22815_ (.A(_05324_),
    .B(_09264_),
    .Y(_01984_));
 sky130_fd_sc_hd__nor2_1 _22816_ (.A(_05573_),
    .B(_09264_),
    .Y(_01985_));
 sky130_fd_sc_hd__nor2_1 _22817_ (.A(_05611_),
    .B(_09264_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_1 _22818_ (.A(_05330_),
    .B(_09264_),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2_1 _22819_ (.A(_05338_),
    .B(_09264_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor2_1 _22820_ (.A(_05347_),
    .B(_09264_),
    .Y(_01989_));
 sky130_fd_sc_hd__nor2_1 _22821_ (.A(_05354_),
    .B(_09264_),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_1 _22822_ (.A(_05360_),
    .B(_09264_),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_1 _22823_ (.A(_05371_),
    .B(_09264_),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _22824_ (.A(_05380_),
    .B(_09264_),
    .Y(_01993_));
 sky130_fd_sc_hd__nand2_8 _22825_ (.A(_09926_),
    .B(_05778_),
    .Y(_09268_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_699 ();
 sky130_fd_sc_hd__nor2_1 _22827_ (.A(_04988_),
    .B(_09268_),
    .Y(_01994_));
 sky130_fd_sc_hd__nor2_1 _22828_ (.A(_05062_),
    .B(_09268_),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_1 _22829_ (.A(_05077_),
    .B(_09268_),
    .Y(_01996_));
 sky130_fd_sc_hd__nor2_1 _22830_ (.A(_05087_),
    .B(_09268_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _22831_ (.A(_05095_),
    .B(_09268_),
    .Y(_01998_));
 sky130_fd_sc_hd__nor2_1 _22832_ (.A(_05102_),
    .B(_09268_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor2_1 _22833_ (.A(_05112_),
    .B(_09268_),
    .Y(_02000_));
 sky130_fd_sc_hd__nor2_1 _22834_ (.A(_05121_),
    .B(_09268_),
    .Y(_02001_));
 sky130_fd_sc_hd__nor2_1 _22835_ (.A(_05128_),
    .B(_09268_),
    .Y(_02002_));
 sky130_fd_sc_hd__nor2_1 _22836_ (.A(_05137_),
    .B(_09268_),
    .Y(_02003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_698 ();
 sky130_fd_sc_hd__nor2_1 _22838_ (.A(_05154_),
    .B(_09268_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_1 _22839_ (.A(_04992_),
    .B(_09268_),
    .Y(_02005_));
 sky130_fd_sc_hd__nor2_1 _22840_ (.A(_05167_),
    .B(_09268_),
    .Y(_02006_));
 sky130_fd_sc_hd__nor2_1 _22841_ (.A(_05175_),
    .B(_09268_),
    .Y(_02007_));
 sky130_fd_sc_hd__nor2_1 _22842_ (.A(_05184_),
    .B(_09268_),
    .Y(_02008_));
 sky130_fd_sc_hd__nor2_1 _22843_ (.A(_05196_),
    .B(_09268_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _22844_ (.A(_05206_),
    .B(_09268_),
    .Y(_02010_));
 sky130_fd_sc_hd__nor2_1 _22845_ (.A(_05214_),
    .B(_09268_),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _22846_ (.A(_05224_),
    .B(_09268_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_1 _22847_ (.A(_05236_),
    .B(_09268_),
    .Y(_02013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_697 ();
 sky130_fd_sc_hd__nor2_1 _22849_ (.A(_05243_),
    .B(_09268_),
    .Y(_02014_));
 sky130_fd_sc_hd__nor2_1 _22850_ (.A(_05251_),
    .B(_09268_),
    .Y(_02015_));
 sky130_fd_sc_hd__nor2_1 _22851_ (.A(_04995_),
    .B(_09268_),
    .Y(_02016_));
 sky130_fd_sc_hd__nor2_1 _22852_ (.A(_05260_),
    .B(_09268_),
    .Y(_02017_));
 sky130_fd_sc_hd__nor2_1 _22853_ (.A(_05310_),
    .B(_09268_),
    .Y(_02018_));
 sky130_fd_sc_hd__nor2_1 _22854_ (.A(_05003_),
    .B(_09268_),
    .Y(_02019_));
 sky130_fd_sc_hd__nor2_1 _22855_ (.A(_05012_),
    .B(_09268_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _22856_ (.A(_05021_),
    .B(_09268_),
    .Y(_02021_));
 sky130_fd_sc_hd__nor2_1 _22857_ (.A(_05032_),
    .B(_09268_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_1 _22858_ (.A(_05039_),
    .B(_09268_),
    .Y(_02023_));
 sky130_fd_sc_hd__nor2_1 _22859_ (.A(_05048_),
    .B(_09268_),
    .Y(_02024_));
 sky130_fd_sc_hd__nor2_1 _22860_ (.A(_05055_),
    .B(_09268_),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_8 _22861_ (.A(_09979_),
    .B(_06133_),
    .Y(_09272_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_696 ();
 sky130_fd_sc_hd__nor2_1 _22863_ (.A(_05317_),
    .B(_09272_),
    .Y(_02026_));
 sky130_fd_sc_hd__nor2_1 _22864_ (.A(_05388_),
    .B(_09272_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _22865_ (.A(_05402_),
    .B(_09272_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _22866_ (.A(_05412_),
    .B(_09272_),
    .Y(_02029_));
 sky130_fd_sc_hd__nor2_1 _22867_ (.A(_05419_),
    .B(_09272_),
    .Y(_02030_));
 sky130_fd_sc_hd__nor2_1 _22868_ (.A(_05426_),
    .B(_09272_),
    .Y(_02031_));
 sky130_fd_sc_hd__nor2_1 _22869_ (.A(_05438_),
    .B(_09272_),
    .Y(_02032_));
 sky130_fd_sc_hd__nor2_1 _22870_ (.A(_05447_),
    .B(_09272_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_1 _22871_ (.A(_05453_),
    .B(_09272_),
    .Y(_02034_));
 sky130_fd_sc_hd__nor2_1 _22872_ (.A(_05465_),
    .B(_09272_),
    .Y(_02035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_695 ();
 sky130_fd_sc_hd__nor2_1 _22874_ (.A(_05480_),
    .B(_09272_),
    .Y(_02036_));
 sky130_fd_sc_hd__nor2_1 _22875_ (.A(_05321_),
    .B(_09272_),
    .Y(_02037_));
 sky130_fd_sc_hd__nor2_1 _22876_ (.A(_05488_),
    .B(_09272_),
    .Y(_02038_));
 sky130_fd_sc_hd__nor2_1 _22877_ (.A(_05498_),
    .B(_09272_),
    .Y(_02039_));
 sky130_fd_sc_hd__nor2_1 _22878_ (.A(_05509_),
    .B(_09272_),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _22879_ (.A(_05515_),
    .B(_09272_),
    .Y(_02041_));
 sky130_fd_sc_hd__nor2_1 _22880_ (.A(_05523_),
    .B(_09272_),
    .Y(_02042_));
 sky130_fd_sc_hd__nor2_1 _22881_ (.A(_05535_),
    .B(_09272_),
    .Y(_02043_));
 sky130_fd_sc_hd__nor2_1 _22882_ (.A(_05542_),
    .B(_09272_),
    .Y(_02044_));
 sky130_fd_sc_hd__nor2_1 _22883_ (.A(_05551_),
    .B(_09272_),
    .Y(_02045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_694 ();
 sky130_fd_sc_hd__nor2_1 _22885_ (.A(_05559_),
    .B(_09272_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_1 _22886_ (.A(_05567_),
    .B(_09272_),
    .Y(_02047_));
 sky130_fd_sc_hd__nor2_1 _22887_ (.A(_05324_),
    .B(_09272_),
    .Y(_02048_));
 sky130_fd_sc_hd__nor2_1 _22888_ (.A(_05573_),
    .B(_09272_),
    .Y(_02049_));
 sky130_fd_sc_hd__nor2_1 _22889_ (.A(_05611_),
    .B(_09272_),
    .Y(_02050_));
 sky130_fd_sc_hd__nor2_1 _22890_ (.A(_05330_),
    .B(_09272_),
    .Y(_02051_));
 sky130_fd_sc_hd__nor2_1 _22891_ (.A(_05338_),
    .B(_09272_),
    .Y(_02052_));
 sky130_fd_sc_hd__nor2_1 _22892_ (.A(_05347_),
    .B(_09272_),
    .Y(_02053_));
 sky130_fd_sc_hd__nor2_1 _22893_ (.A(_05354_),
    .B(_09272_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _22894_ (.A(_05360_),
    .B(_09272_),
    .Y(_02055_));
 sky130_fd_sc_hd__nor2_1 _22895_ (.A(_05371_),
    .B(_09272_),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_1 _22896_ (.A(_05380_),
    .B(_09272_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_8 _22897_ (.A(_09933_),
    .B(_04982_),
    .Y(_09276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_693 ();
 sky130_fd_sc_hd__nor2_1 _22899_ (.A(_04988_),
    .B(_09276_),
    .Y(_02058_));
 sky130_fd_sc_hd__nor2_1 _22900_ (.A(_05062_),
    .B(_09276_),
    .Y(_02059_));
 sky130_fd_sc_hd__nor2_1 _22901_ (.A(_05077_),
    .B(_09276_),
    .Y(_02060_));
 sky130_fd_sc_hd__nor2_1 _22902_ (.A(_05087_),
    .B(_09276_),
    .Y(_02061_));
 sky130_fd_sc_hd__nor2_1 _22903_ (.A(_05095_),
    .B(_09276_),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _22904_ (.A(_05102_),
    .B(_09276_),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_1 _22905_ (.A(_05112_),
    .B(_09276_),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _22906_ (.A(_05121_),
    .B(_09276_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor2_1 _22907_ (.A(_05128_),
    .B(_09276_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _22908_ (.A(_05137_),
    .B(_09276_),
    .Y(_02067_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_692 ();
 sky130_fd_sc_hd__nor2_1 _22910_ (.A(_05154_),
    .B(_09276_),
    .Y(_02068_));
 sky130_fd_sc_hd__nor2_1 _22911_ (.A(_04992_),
    .B(_09276_),
    .Y(_02069_));
 sky130_fd_sc_hd__nor2_1 _22912_ (.A(_05167_),
    .B(_09276_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_1 _22913_ (.A(_05175_),
    .B(_09276_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_1 _22914_ (.A(_05184_),
    .B(_09276_),
    .Y(_02072_));
 sky130_fd_sc_hd__nor2_1 _22915_ (.A(_05196_),
    .B(_09276_),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_1 _22916_ (.A(_05206_),
    .B(_09276_),
    .Y(_02074_));
 sky130_fd_sc_hd__nor2_1 _22917_ (.A(_05214_),
    .B(_09276_),
    .Y(_02075_));
 sky130_fd_sc_hd__nor2_1 _22918_ (.A(_05224_),
    .B(_09276_),
    .Y(_02076_));
 sky130_fd_sc_hd__nor2_1 _22919_ (.A(_05236_),
    .B(_09276_),
    .Y(_02077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_691 ();
 sky130_fd_sc_hd__nor2_1 _22921_ (.A(_05243_),
    .B(_09276_),
    .Y(_02078_));
 sky130_fd_sc_hd__nor2_1 _22922_ (.A(_05251_),
    .B(_09276_),
    .Y(_02079_));
 sky130_fd_sc_hd__nor2_1 _22923_ (.A(_04995_),
    .B(_09276_),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _22924_ (.A(_05260_),
    .B(_09276_),
    .Y(_02081_));
 sky130_fd_sc_hd__nor2_1 _22925_ (.A(_05310_),
    .B(_09276_),
    .Y(_02082_));
 sky130_fd_sc_hd__nor2_1 _22926_ (.A(_05003_),
    .B(_09276_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_1 _22927_ (.A(_05012_),
    .B(_09276_),
    .Y(_02084_));
 sky130_fd_sc_hd__nor2_1 _22928_ (.A(_05021_),
    .B(_09276_),
    .Y(_02085_));
 sky130_fd_sc_hd__nor2_1 _22929_ (.A(_05032_),
    .B(_09276_),
    .Y(_02086_));
 sky130_fd_sc_hd__nor2_1 _22930_ (.A(_05039_),
    .B(_09276_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor2_1 _22931_ (.A(_05048_),
    .B(_09276_),
    .Y(_02088_));
 sky130_fd_sc_hd__nor2_1 _22932_ (.A(_05055_),
    .B(_09276_),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_8 _22933_ (.A(_09986_),
    .B(_05313_),
    .Y(_09280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_690 ();
 sky130_fd_sc_hd__nor2_1 _22935_ (.A(_05317_),
    .B(_09280_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _22936_ (.A(_05388_),
    .B(_09280_),
    .Y(_02091_));
 sky130_fd_sc_hd__nor2_1 _22937_ (.A(_05402_),
    .B(_09280_),
    .Y(_02092_));
 sky130_fd_sc_hd__nor2_1 _22938_ (.A(_05412_),
    .B(_09280_),
    .Y(_02093_));
 sky130_fd_sc_hd__nor2_1 _22939_ (.A(_05419_),
    .B(_09280_),
    .Y(_02094_));
 sky130_fd_sc_hd__nor2_1 _22940_ (.A(_05426_),
    .B(_09280_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor2_1 _22941_ (.A(_05438_),
    .B(_09280_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_1 _22942_ (.A(_05447_),
    .B(_09280_),
    .Y(_02097_));
 sky130_fd_sc_hd__nor2_1 _22943_ (.A(_05453_),
    .B(_09280_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_1 _22944_ (.A(_05465_),
    .B(_09280_),
    .Y(_02099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_689 ();
 sky130_fd_sc_hd__nor2_1 _22946_ (.A(_05480_),
    .B(_09280_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_1 _22947_ (.A(_05321_),
    .B(_09280_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor2_1 _22948_ (.A(_05488_),
    .B(_09280_),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _22949_ (.A(_05498_),
    .B(_09280_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _22950_ (.A(_05509_),
    .B(_09280_),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _22951_ (.A(_05515_),
    .B(_09280_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _22952_ (.A(_05523_),
    .B(_09280_),
    .Y(_02106_));
 sky130_fd_sc_hd__nor2_1 _22953_ (.A(_05535_),
    .B(_09280_),
    .Y(_02107_));
 sky130_fd_sc_hd__nor2_1 _22954_ (.A(_05542_),
    .B(_09280_),
    .Y(_02108_));
 sky130_fd_sc_hd__nor2_1 _22955_ (.A(_05551_),
    .B(_09280_),
    .Y(_02109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_688 ();
 sky130_fd_sc_hd__nor2_1 _22957_ (.A(_05559_),
    .B(_09280_),
    .Y(_02110_));
 sky130_fd_sc_hd__nor2_1 _22958_ (.A(_05567_),
    .B(_09280_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor2_1 _22959_ (.A(_05324_),
    .B(_09280_),
    .Y(_02112_));
 sky130_fd_sc_hd__nor2_1 _22960_ (.A(_05573_),
    .B(_09280_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor2_1 _22961_ (.A(_05611_),
    .B(_09280_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _22962_ (.A(_05330_),
    .B(_09280_),
    .Y(_02115_));
 sky130_fd_sc_hd__nor2_1 _22963_ (.A(_05338_),
    .B(_09280_),
    .Y(_02116_));
 sky130_fd_sc_hd__nor2_1 _22964_ (.A(_05347_),
    .B(_09280_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _22965_ (.A(_05354_),
    .B(_09280_),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_1 _22966_ (.A(_05360_),
    .B(_09280_),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _22967_ (.A(_05371_),
    .B(_09280_),
    .Y(_02120_));
 sky130_fd_sc_hd__nor2_1 _22968_ (.A(_05380_),
    .B(_09280_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_8 _22969_ (.A(_09933_),
    .B(_05614_),
    .Y(_09284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_687 ();
 sky130_fd_sc_hd__nor2_1 _22971_ (.A(_04988_),
    .B(_09284_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _22972_ (.A(_05062_),
    .B(_09284_),
    .Y(_02123_));
 sky130_fd_sc_hd__nor2_1 _22973_ (.A(_05077_),
    .B(_09284_),
    .Y(_02124_));
 sky130_fd_sc_hd__nor2_1 _22974_ (.A(_05087_),
    .B(_09284_),
    .Y(_02125_));
 sky130_fd_sc_hd__nor2_1 _22975_ (.A(_05095_),
    .B(_09284_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor2_1 _22976_ (.A(_05102_),
    .B(_09284_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _22977_ (.A(_05112_),
    .B(_09284_),
    .Y(_02128_));
 sky130_fd_sc_hd__nor2_1 _22978_ (.A(_05121_),
    .B(_09284_),
    .Y(_02129_));
 sky130_fd_sc_hd__nor2_1 _22979_ (.A(_05128_),
    .B(_09284_),
    .Y(_02130_));
 sky130_fd_sc_hd__nor2_1 _22980_ (.A(_05137_),
    .B(_09284_),
    .Y(_02131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_686 ();
 sky130_fd_sc_hd__nor2_1 _22982_ (.A(_05154_),
    .B(_09284_),
    .Y(_02132_));
 sky130_fd_sc_hd__nor2_1 _22983_ (.A(_04992_),
    .B(_09284_),
    .Y(_02133_));
 sky130_fd_sc_hd__nor2_1 _22984_ (.A(_05167_),
    .B(_09284_),
    .Y(_02134_));
 sky130_fd_sc_hd__nor2_1 _22985_ (.A(_05175_),
    .B(_09284_),
    .Y(_02135_));
 sky130_fd_sc_hd__nor2_1 _22986_ (.A(_05184_),
    .B(_09284_),
    .Y(_02136_));
 sky130_fd_sc_hd__nor2_1 _22987_ (.A(_05196_),
    .B(_09284_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _22988_ (.A(_05206_),
    .B(_09284_),
    .Y(_02138_));
 sky130_fd_sc_hd__nor2_1 _22989_ (.A(_05214_),
    .B(_09284_),
    .Y(_02139_));
 sky130_fd_sc_hd__nor2_1 _22990_ (.A(_05224_),
    .B(_09284_),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2_1 _22991_ (.A(_05236_),
    .B(_09284_),
    .Y(_02141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_685 ();
 sky130_fd_sc_hd__nor2_1 _22993_ (.A(_05243_),
    .B(_09284_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _22994_ (.A(_05251_),
    .B(_09284_),
    .Y(_02143_));
 sky130_fd_sc_hd__nor2_1 _22995_ (.A(_04995_),
    .B(_09284_),
    .Y(_02144_));
 sky130_fd_sc_hd__nor2_1 _22996_ (.A(_05260_),
    .B(_09284_),
    .Y(_02145_));
 sky130_fd_sc_hd__nor2_1 _22997_ (.A(_05310_),
    .B(_09284_),
    .Y(_02146_));
 sky130_fd_sc_hd__nor2_1 _22998_ (.A(_05003_),
    .B(_09284_),
    .Y(_02147_));
 sky130_fd_sc_hd__nor2_1 _22999_ (.A(_05012_),
    .B(_09284_),
    .Y(_02148_));
 sky130_fd_sc_hd__nor2_1 _23000_ (.A(_05021_),
    .B(_09284_),
    .Y(_02149_));
 sky130_fd_sc_hd__nor2_1 _23001_ (.A(_05032_),
    .B(_09284_),
    .Y(_02150_));
 sky130_fd_sc_hd__nor2_1 _23002_ (.A(_05039_),
    .B(_09284_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_1 _23003_ (.A(_05048_),
    .B(_09284_),
    .Y(_02152_));
 sky130_fd_sc_hd__nor2_1 _23004_ (.A(_05055_),
    .B(_09284_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_8 _23005_ (.A(_09986_),
    .B(_05655_),
    .Y(_09288_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_684 ();
 sky130_fd_sc_hd__nor2_1 _23007_ (.A(_05317_),
    .B(_09288_),
    .Y(_02154_));
 sky130_fd_sc_hd__nor2_1 _23008_ (.A(_05388_),
    .B(_09288_),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _23009_ (.A(_05402_),
    .B(_09288_),
    .Y(_02156_));
 sky130_fd_sc_hd__nor2_1 _23010_ (.A(_05412_),
    .B(_09288_),
    .Y(_02157_));
 sky130_fd_sc_hd__nor2_1 _23011_ (.A(_05419_),
    .B(_09288_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _23012_ (.A(_05426_),
    .B(_09288_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _23013_ (.A(_05438_),
    .B(_09288_),
    .Y(_02160_));
 sky130_fd_sc_hd__nor2_1 _23014_ (.A(_05447_),
    .B(_09288_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_1 _23015_ (.A(_05453_),
    .B(_09288_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _23016_ (.A(_05465_),
    .B(_09288_),
    .Y(_02163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_683 ();
 sky130_fd_sc_hd__nor2_1 _23018_ (.A(_05480_),
    .B(_09288_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _23019_ (.A(_05321_),
    .B(_09288_),
    .Y(_02165_));
 sky130_fd_sc_hd__nor2_1 _23020_ (.A(_05488_),
    .B(_09288_),
    .Y(_02166_));
 sky130_fd_sc_hd__nor2_1 _23021_ (.A(_05498_),
    .B(_09288_),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _23022_ (.A(_05509_),
    .B(_09288_),
    .Y(_02168_));
 sky130_fd_sc_hd__nor2_1 _23023_ (.A(_05515_),
    .B(_09288_),
    .Y(_02169_));
 sky130_fd_sc_hd__nor2_1 _23024_ (.A(_05523_),
    .B(_09288_),
    .Y(_02170_));
 sky130_fd_sc_hd__nor2_1 _23025_ (.A(_05535_),
    .B(_09288_),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_1 _23026_ (.A(_05542_),
    .B(_09288_),
    .Y(_02172_));
 sky130_fd_sc_hd__nor2_1 _23027_ (.A(_05551_),
    .B(_09288_),
    .Y(_02173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_682 ();
 sky130_fd_sc_hd__nor2_1 _23029_ (.A(_05559_),
    .B(_09288_),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_1 _23030_ (.A(_05567_),
    .B(_09288_),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _23031_ (.A(_05324_),
    .B(_09288_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _23032_ (.A(_05573_),
    .B(_09288_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _23033_ (.A(_05611_),
    .B(_09288_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _23034_ (.A(_05330_),
    .B(_09288_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_1 _23035_ (.A(_05338_),
    .B(_09288_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _23036_ (.A(_05347_),
    .B(_09288_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_1 _23037_ (.A(_05354_),
    .B(_09288_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_1 _23038_ (.A(_05360_),
    .B(_09288_),
    .Y(_02183_));
 sky130_fd_sc_hd__nor2_1 _23039_ (.A(_05371_),
    .B(_09288_),
    .Y(_02184_));
 sky130_fd_sc_hd__nor2_1 _23040_ (.A(_05380_),
    .B(_09288_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand2_8 _23041_ (.A(_09933_),
    .B(_05696_),
    .Y(_09292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_681 ();
 sky130_fd_sc_hd__nor2_1 _23043_ (.A(_04988_),
    .B(_09292_),
    .Y(_02186_));
 sky130_fd_sc_hd__nor2_1 _23044_ (.A(_05062_),
    .B(_09292_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _23045_ (.A(_05077_),
    .B(_09292_),
    .Y(_02188_));
 sky130_fd_sc_hd__nor2_1 _23046_ (.A(_05087_),
    .B(_09292_),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _23047_ (.A(_05095_),
    .B(_09292_),
    .Y(_02190_));
 sky130_fd_sc_hd__nor2_1 _23048_ (.A(_05102_),
    .B(_09292_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _23049_ (.A(_05112_),
    .B(_09292_),
    .Y(_02192_));
 sky130_fd_sc_hd__nor2_1 _23050_ (.A(_05121_),
    .B(_09292_),
    .Y(_02193_));
 sky130_fd_sc_hd__nor2_1 _23051_ (.A(_05128_),
    .B(_09292_),
    .Y(_02194_));
 sky130_fd_sc_hd__nor2_1 _23052_ (.A(_05137_),
    .B(_09292_),
    .Y(_02195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_680 ();
 sky130_fd_sc_hd__nor2_1 _23054_ (.A(_05154_),
    .B(_09292_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _23055_ (.A(_04992_),
    .B(_09292_),
    .Y(_02197_));
 sky130_fd_sc_hd__nor2_1 _23056_ (.A(_05167_),
    .B(_09292_),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _23057_ (.A(_05175_),
    .B(_09292_),
    .Y(_02199_));
 sky130_fd_sc_hd__nor2_1 _23058_ (.A(_05184_),
    .B(_09292_),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_1 _23059_ (.A(_05196_),
    .B(_09292_),
    .Y(_02201_));
 sky130_fd_sc_hd__nor2_1 _23060_ (.A(_05206_),
    .B(_09292_),
    .Y(_02202_));
 sky130_fd_sc_hd__nor2_1 _23061_ (.A(_05214_),
    .B(_09292_),
    .Y(_02203_));
 sky130_fd_sc_hd__nor2_1 _23062_ (.A(_05224_),
    .B(_09292_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _23063_ (.A(_05236_),
    .B(_09292_),
    .Y(_02205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_679 ();
 sky130_fd_sc_hd__nor2_1 _23065_ (.A(_05243_),
    .B(_09292_),
    .Y(_02206_));
 sky130_fd_sc_hd__nor2_1 _23066_ (.A(_05251_),
    .B(_09292_),
    .Y(_02207_));
 sky130_fd_sc_hd__nor2_1 _23067_ (.A(_04995_),
    .B(_09292_),
    .Y(_02208_));
 sky130_fd_sc_hd__nor2_1 _23068_ (.A(_05260_),
    .B(_09292_),
    .Y(_02209_));
 sky130_fd_sc_hd__nor2_1 _23069_ (.A(_05310_),
    .B(_09292_),
    .Y(_02210_));
 sky130_fd_sc_hd__nor2_1 _23070_ (.A(_05003_),
    .B(_09292_),
    .Y(_02211_));
 sky130_fd_sc_hd__nor2_1 _23071_ (.A(_05012_),
    .B(_09292_),
    .Y(_02212_));
 sky130_fd_sc_hd__nor2_1 _23072_ (.A(_05021_),
    .B(_09292_),
    .Y(_02213_));
 sky130_fd_sc_hd__nor2_1 _23073_ (.A(_05032_),
    .B(_09292_),
    .Y(_02214_));
 sky130_fd_sc_hd__nor2_1 _23074_ (.A(_05039_),
    .B(_09292_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _23075_ (.A(_05048_),
    .B(_09292_),
    .Y(_02216_));
 sky130_fd_sc_hd__nor2_1 _23076_ (.A(_05055_),
    .B(_09292_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_8 _23077_ (.A(_09986_),
    .B(_05737_),
    .Y(_09296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_678 ();
 sky130_fd_sc_hd__nor2_1 _23079_ (.A(_05317_),
    .B(_09296_),
    .Y(_02218_));
 sky130_fd_sc_hd__nor2_1 _23080_ (.A(_05388_),
    .B(_09296_),
    .Y(_02219_));
 sky130_fd_sc_hd__nor2_1 _23081_ (.A(_05402_),
    .B(_09296_),
    .Y(_02220_));
 sky130_fd_sc_hd__nor2_1 _23082_ (.A(_05412_),
    .B(_09296_),
    .Y(_02221_));
 sky130_fd_sc_hd__nor2_1 _23083_ (.A(_05419_),
    .B(_09296_),
    .Y(_02222_));
 sky130_fd_sc_hd__nor2_1 _23084_ (.A(_05426_),
    .B(_09296_),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _23085_ (.A(_05438_),
    .B(_09296_),
    .Y(_02224_));
 sky130_fd_sc_hd__nor2_1 _23086_ (.A(_05447_),
    .B(_09296_),
    .Y(_02225_));
 sky130_fd_sc_hd__nor2_1 _23087_ (.A(_05453_),
    .B(_09296_),
    .Y(_02226_));
 sky130_fd_sc_hd__nor2_1 _23088_ (.A(_05465_),
    .B(_09296_),
    .Y(_02227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_677 ();
 sky130_fd_sc_hd__nor2_1 _23090_ (.A(_05480_),
    .B(_09296_),
    .Y(_02228_));
 sky130_fd_sc_hd__nor2_1 _23091_ (.A(_05321_),
    .B(_09296_),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _23092_ (.A(_05488_),
    .B(_09296_),
    .Y(_02230_));
 sky130_fd_sc_hd__nor2_1 _23093_ (.A(_05498_),
    .B(_09296_),
    .Y(_02231_));
 sky130_fd_sc_hd__nor2_1 _23094_ (.A(_05509_),
    .B(_09296_),
    .Y(_02232_));
 sky130_fd_sc_hd__nor2_1 _23095_ (.A(_05515_),
    .B(_09296_),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_1 _23096_ (.A(_05523_),
    .B(_09296_),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _23097_ (.A(_05535_),
    .B(_09296_),
    .Y(_02235_));
 sky130_fd_sc_hd__nor2_1 _23098_ (.A(_05542_),
    .B(_09296_),
    .Y(_02236_));
 sky130_fd_sc_hd__nor2_1 _23099_ (.A(_05551_),
    .B(_09296_),
    .Y(_02237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_676 ();
 sky130_fd_sc_hd__nor2_1 _23101_ (.A(_05559_),
    .B(_09296_),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_1 _23102_ (.A(_05567_),
    .B(_09296_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _23103_ (.A(_05324_),
    .B(_09296_),
    .Y(_02240_));
 sky130_fd_sc_hd__nor2_1 _23104_ (.A(_05573_),
    .B(_09296_),
    .Y(_02241_));
 sky130_fd_sc_hd__nor2_1 _23105_ (.A(_05611_),
    .B(_09296_),
    .Y(_02242_));
 sky130_fd_sc_hd__nor2_1 _23106_ (.A(_05330_),
    .B(_09296_),
    .Y(_02243_));
 sky130_fd_sc_hd__nor2_1 _23107_ (.A(_05338_),
    .B(_09296_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_1 _23108_ (.A(_05347_),
    .B(_09296_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _23109_ (.A(_05354_),
    .B(_09296_),
    .Y(_02246_));
 sky130_fd_sc_hd__nor2_1 _23110_ (.A(_05360_),
    .B(_09296_),
    .Y(_02247_));
 sky130_fd_sc_hd__nor2_1 _23111_ (.A(_05371_),
    .B(_09296_),
    .Y(_02248_));
 sky130_fd_sc_hd__nor2_1 _23112_ (.A(_05380_),
    .B(_09296_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_8 _23113_ (.A(_09933_),
    .B(_05778_),
    .Y(_09300_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_675 ();
 sky130_fd_sc_hd__nor2_1 _23115_ (.A(_04988_),
    .B(_09300_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _23116_ (.A(_05062_),
    .B(_09300_),
    .Y(_02251_));
 sky130_fd_sc_hd__nor2_1 _23117_ (.A(_05077_),
    .B(_09300_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor2_1 _23118_ (.A(_05087_),
    .B(_09300_),
    .Y(_02253_));
 sky130_fd_sc_hd__nor2_1 _23119_ (.A(_05095_),
    .B(_09300_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor2_1 _23120_ (.A(_05102_),
    .B(_09300_),
    .Y(_02255_));
 sky130_fd_sc_hd__nor2_1 _23121_ (.A(_05112_),
    .B(_09300_),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_1 _23122_ (.A(_05121_),
    .B(_09300_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _23123_ (.A(_05128_),
    .B(_09300_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _23124_ (.A(_05137_),
    .B(_09300_),
    .Y(_02259_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_674 ();
 sky130_fd_sc_hd__nor2_1 _23126_ (.A(_05154_),
    .B(_09300_),
    .Y(_02260_));
 sky130_fd_sc_hd__nor2_1 _23127_ (.A(_04992_),
    .B(_09300_),
    .Y(_02261_));
 sky130_fd_sc_hd__nor2_1 _23128_ (.A(_05167_),
    .B(_09300_),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_1 _23129_ (.A(_05175_),
    .B(_09300_),
    .Y(_02263_));
 sky130_fd_sc_hd__nor2_1 _23130_ (.A(_05184_),
    .B(_09300_),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _23131_ (.A(_05196_),
    .B(_09300_),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _23132_ (.A(_05206_),
    .B(_09300_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_1 _23133_ (.A(_05214_),
    .B(_09300_),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _23134_ (.A(_05224_),
    .B(_09300_),
    .Y(_02268_));
 sky130_fd_sc_hd__nor2_1 _23135_ (.A(_05236_),
    .B(_09300_),
    .Y(_02269_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_673 ();
 sky130_fd_sc_hd__nor2_1 _23137_ (.A(_05243_),
    .B(_09300_),
    .Y(_02270_));
 sky130_fd_sc_hd__nor2_1 _23138_ (.A(_05251_),
    .B(_09300_),
    .Y(_02271_));
 sky130_fd_sc_hd__nor2_1 _23139_ (.A(_04995_),
    .B(_09300_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _23140_ (.A(_05260_),
    .B(_09300_),
    .Y(_02273_));
 sky130_fd_sc_hd__nor2_1 _23141_ (.A(_05310_),
    .B(_09300_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _23142_ (.A(_05003_),
    .B(_09300_),
    .Y(_02275_));
 sky130_fd_sc_hd__nor2_1 _23143_ (.A(_05012_),
    .B(_09300_),
    .Y(_02276_));
 sky130_fd_sc_hd__nor2_1 _23144_ (.A(_05021_),
    .B(_09300_),
    .Y(_02277_));
 sky130_fd_sc_hd__nor2_1 _23145_ (.A(_05032_),
    .B(_09300_),
    .Y(_02278_));
 sky130_fd_sc_hd__nor2_1 _23146_ (.A(_05039_),
    .B(_09300_),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_1 _23147_ (.A(_05048_),
    .B(_09300_),
    .Y(_02280_));
 sky130_fd_sc_hd__nor2_1 _23148_ (.A(_05055_),
    .B(_09300_),
    .Y(_02281_));
 sky130_fd_sc_hd__or3_4 _23149_ (.A(net762),
    .B(_09977_),
    .C(_09955_),
    .X(_09304_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_671 ();
 sky130_fd_sc_hd__nor2_1 _23152_ (.A(_05317_),
    .B(_09304_),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2_1 _23153_ (.A(_05388_),
    .B(_09304_),
    .Y(_02283_));
 sky130_fd_sc_hd__nor2_1 _23154_ (.A(_05402_),
    .B(_09304_),
    .Y(_02284_));
 sky130_fd_sc_hd__nor2_1 _23155_ (.A(_05412_),
    .B(_09304_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _23156_ (.A(_05419_),
    .B(_09304_),
    .Y(_02286_));
 sky130_fd_sc_hd__nor2_1 _23157_ (.A(_05426_),
    .B(_09304_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_1 _23158_ (.A(_05438_),
    .B(_09304_),
    .Y(_02288_));
 sky130_fd_sc_hd__nor2_1 _23159_ (.A(_05447_),
    .B(_09304_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _23160_ (.A(_05453_),
    .B(_09304_),
    .Y(_02290_));
 sky130_fd_sc_hd__nor2_1 _23161_ (.A(_05465_),
    .B(_09304_),
    .Y(_02291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_670 ();
 sky130_fd_sc_hd__nor2_1 _23163_ (.A(_05480_),
    .B(_09304_),
    .Y(_02292_));
 sky130_fd_sc_hd__nor2_1 _23164_ (.A(_05321_),
    .B(_09304_),
    .Y(_02293_));
 sky130_fd_sc_hd__nor2_1 _23165_ (.A(_05488_),
    .B(_09304_),
    .Y(_02294_));
 sky130_fd_sc_hd__nor2_1 _23166_ (.A(_05498_),
    .B(_09304_),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_1 _23167_ (.A(_05509_),
    .B(_09304_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor2_1 _23168_ (.A(_05515_),
    .B(_09304_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _23169_ (.A(_05523_),
    .B(_09304_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _23170_ (.A(_05535_),
    .B(_09304_),
    .Y(_02299_));
 sky130_fd_sc_hd__nor2_1 _23171_ (.A(_05542_),
    .B(_09304_),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _23172_ (.A(_05551_),
    .B(_09304_),
    .Y(_02301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_669 ();
 sky130_fd_sc_hd__nor2_1 _23174_ (.A(_05559_),
    .B(_09304_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _23175_ (.A(_05567_),
    .B(_09304_),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _23176_ (.A(_05324_),
    .B(_09304_),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _23177_ (.A(_05573_),
    .B(_09304_),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _23178_ (.A(_05611_),
    .B(_09304_),
    .Y(_02306_));
 sky130_fd_sc_hd__nor2_1 _23179_ (.A(_05330_),
    .B(_09304_),
    .Y(_02307_));
 sky130_fd_sc_hd__nor2_1 _23180_ (.A(_05338_),
    .B(_09304_),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2_1 _23181_ (.A(_05347_),
    .B(_09304_),
    .Y(_02309_));
 sky130_fd_sc_hd__nor2_1 _23182_ (.A(_05354_),
    .B(_09304_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor2_1 _23183_ (.A(_05360_),
    .B(_09304_),
    .Y(_02311_));
 sky130_fd_sc_hd__nor2_1 _23184_ (.A(_05371_),
    .B(_09304_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _23185_ (.A(_05380_),
    .B(_09304_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_8 _23186_ (.A(_09940_),
    .B(_04982_),
    .Y(_09309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_668 ();
 sky130_fd_sc_hd__nor2_1 _23188_ (.A(_04988_),
    .B(_09309_),
    .Y(_02314_));
 sky130_fd_sc_hd__nor2_1 _23189_ (.A(_05062_),
    .B(_09309_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _23190_ (.A(_05077_),
    .B(_09309_),
    .Y(_02316_));
 sky130_fd_sc_hd__nor2_1 _23191_ (.A(_05087_),
    .B(_09309_),
    .Y(_02317_));
 sky130_fd_sc_hd__nor2_1 _23192_ (.A(_05095_),
    .B(_09309_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_1 _23193_ (.A(_05102_),
    .B(_09309_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _23194_ (.A(_05112_),
    .B(_09309_),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _23195_ (.A(_05121_),
    .B(_09309_),
    .Y(_02321_));
 sky130_fd_sc_hd__nor2_1 _23196_ (.A(_05128_),
    .B(_09309_),
    .Y(_02322_));
 sky130_fd_sc_hd__nor2_1 _23197_ (.A(_05137_),
    .B(_09309_),
    .Y(_02323_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_667 ();
 sky130_fd_sc_hd__nor2_1 _23199_ (.A(_05154_),
    .B(_09309_),
    .Y(_02324_));
 sky130_fd_sc_hd__nor2_1 _23200_ (.A(_04992_),
    .B(_09309_),
    .Y(_02325_));
 sky130_fd_sc_hd__nor2_1 _23201_ (.A(_05167_),
    .B(_09309_),
    .Y(_02326_));
 sky130_fd_sc_hd__nor2_1 _23202_ (.A(_05175_),
    .B(_09309_),
    .Y(_02327_));
 sky130_fd_sc_hd__nor2_1 _23203_ (.A(_05184_),
    .B(_09309_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_1 _23204_ (.A(_05196_),
    .B(_09309_),
    .Y(_02329_));
 sky130_fd_sc_hd__nor2_1 _23205_ (.A(_05206_),
    .B(_09309_),
    .Y(_02330_));
 sky130_fd_sc_hd__nor2_1 _23206_ (.A(_05214_),
    .B(_09309_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_1 _23207_ (.A(_05224_),
    .B(_09309_),
    .Y(_02332_));
 sky130_fd_sc_hd__nor2_1 _23208_ (.A(_05236_),
    .B(_09309_),
    .Y(_02333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_666 ();
 sky130_fd_sc_hd__nor2_1 _23210_ (.A(_05243_),
    .B(_09309_),
    .Y(_02334_));
 sky130_fd_sc_hd__nor2_1 _23211_ (.A(_05251_),
    .B(_09309_),
    .Y(_02335_));
 sky130_fd_sc_hd__nor2_1 _23212_ (.A(_04995_),
    .B(_09309_),
    .Y(_02336_));
 sky130_fd_sc_hd__nor2_1 _23213_ (.A(_05260_),
    .B(_09309_),
    .Y(_02337_));
 sky130_fd_sc_hd__nor2_1 _23214_ (.A(_05310_),
    .B(_09309_),
    .Y(_02338_));
 sky130_fd_sc_hd__nor2_1 _23215_ (.A(_05003_),
    .B(_09309_),
    .Y(_02339_));
 sky130_fd_sc_hd__nor2_1 _23216_ (.A(_05012_),
    .B(_09309_),
    .Y(_02340_));
 sky130_fd_sc_hd__nor2_1 _23217_ (.A(_05021_),
    .B(_09309_),
    .Y(_02341_));
 sky130_fd_sc_hd__nor2_1 _23218_ (.A(_05032_),
    .B(_09309_),
    .Y(_02342_));
 sky130_fd_sc_hd__nor2_1 _23219_ (.A(_05039_),
    .B(_09309_),
    .Y(_02343_));
 sky130_fd_sc_hd__nor2_1 _23220_ (.A(_05048_),
    .B(_09309_),
    .Y(_02344_));
 sky130_fd_sc_hd__nor2_1 _23221_ (.A(_05055_),
    .B(_09309_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand2_8 _23222_ (.A(_09991_),
    .B(_05313_),
    .Y(_09313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_665 ();
 sky130_fd_sc_hd__nor2_1 _23224_ (.A(_05317_),
    .B(_09313_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _23225_ (.A(_05388_),
    .B(_09313_),
    .Y(_02347_));
 sky130_fd_sc_hd__nor2_1 _23226_ (.A(_05402_),
    .B(_09313_),
    .Y(_02348_));
 sky130_fd_sc_hd__nor2_1 _23227_ (.A(_05412_),
    .B(_09313_),
    .Y(_02349_));
 sky130_fd_sc_hd__nor2_1 _23228_ (.A(_05419_),
    .B(_09313_),
    .Y(_02350_));
 sky130_fd_sc_hd__nor2_1 _23229_ (.A(_05426_),
    .B(_09313_),
    .Y(_02351_));
 sky130_fd_sc_hd__nor2_1 _23230_ (.A(_05438_),
    .B(_09313_),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_1 _23231_ (.A(_05447_),
    .B(_09313_),
    .Y(_02353_));
 sky130_fd_sc_hd__nor2_1 _23232_ (.A(_05453_),
    .B(_09313_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _23233_ (.A(_05465_),
    .B(_09313_),
    .Y(_02355_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_664 ();
 sky130_fd_sc_hd__nor2_1 _23235_ (.A(_05480_),
    .B(_09313_),
    .Y(_02356_));
 sky130_fd_sc_hd__nor2_1 _23236_ (.A(_05321_),
    .B(_09313_),
    .Y(_02357_));
 sky130_fd_sc_hd__nor2_1 _23237_ (.A(_05488_),
    .B(_09313_),
    .Y(_02358_));
 sky130_fd_sc_hd__nor2_1 _23238_ (.A(_05498_),
    .B(_09313_),
    .Y(_02359_));
 sky130_fd_sc_hd__nor2_1 _23239_ (.A(_05509_),
    .B(_09313_),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_1 _23240_ (.A(_05515_),
    .B(_09313_),
    .Y(_02361_));
 sky130_fd_sc_hd__nor2_1 _23241_ (.A(_05523_),
    .B(_09313_),
    .Y(_02362_));
 sky130_fd_sc_hd__nor2_1 _23242_ (.A(_05535_),
    .B(_09313_),
    .Y(_02363_));
 sky130_fd_sc_hd__nor2_1 _23243_ (.A(_05542_),
    .B(_09313_),
    .Y(_02364_));
 sky130_fd_sc_hd__nor2_1 _23244_ (.A(_05551_),
    .B(_09313_),
    .Y(_02365_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_663 ();
 sky130_fd_sc_hd__nor2_1 _23246_ (.A(_05559_),
    .B(_09313_),
    .Y(_02366_));
 sky130_fd_sc_hd__nor2_1 _23247_ (.A(_05567_),
    .B(_09313_),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_1 _23248_ (.A(_05324_),
    .B(_09313_),
    .Y(_02368_));
 sky130_fd_sc_hd__nor2_1 _23249_ (.A(_05573_),
    .B(_09313_),
    .Y(_02369_));
 sky130_fd_sc_hd__nor2_1 _23250_ (.A(_05611_),
    .B(_09313_),
    .Y(_02370_));
 sky130_fd_sc_hd__nor2_1 _23251_ (.A(_05330_),
    .B(_09313_),
    .Y(_02371_));
 sky130_fd_sc_hd__nor2_1 _23252_ (.A(_05338_),
    .B(_09313_),
    .Y(_02372_));
 sky130_fd_sc_hd__nor2_1 _23253_ (.A(_05347_),
    .B(_09313_),
    .Y(_02373_));
 sky130_fd_sc_hd__nor2_1 _23254_ (.A(_05354_),
    .B(_09313_),
    .Y(_02374_));
 sky130_fd_sc_hd__nor2_1 _23255_ (.A(_05360_),
    .B(_09313_),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2_1 _23256_ (.A(_05371_),
    .B(_09313_),
    .Y(_02376_));
 sky130_fd_sc_hd__nor2_1 _23257_ (.A(_05380_),
    .B(_09313_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_8 _23258_ (.A(_09940_),
    .B(_05614_),
    .Y(_09317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_662 ();
 sky130_fd_sc_hd__nor2_1 _23260_ (.A(_04988_),
    .B(_09317_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _23261_ (.A(_05062_),
    .B(_09317_),
    .Y(_02379_));
 sky130_fd_sc_hd__nor2_1 _23262_ (.A(_05077_),
    .B(_09317_),
    .Y(_02380_));
 sky130_fd_sc_hd__nor2_1 _23263_ (.A(_05087_),
    .B(_09317_),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_1 _23264_ (.A(_05095_),
    .B(_09317_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor2_1 _23265_ (.A(_05102_),
    .B(_09317_),
    .Y(_02383_));
 sky130_fd_sc_hd__nor2_1 _23266_ (.A(_05112_),
    .B(_09317_),
    .Y(_02384_));
 sky130_fd_sc_hd__nor2_1 _23267_ (.A(_05121_),
    .B(_09317_),
    .Y(_02385_));
 sky130_fd_sc_hd__nor2_1 _23268_ (.A(_05128_),
    .B(_09317_),
    .Y(_02386_));
 sky130_fd_sc_hd__nor2_1 _23269_ (.A(_05137_),
    .B(_09317_),
    .Y(_02387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_661 ();
 sky130_fd_sc_hd__nor2_1 _23271_ (.A(_05154_),
    .B(_09317_),
    .Y(_02388_));
 sky130_fd_sc_hd__nor2_1 _23272_ (.A(_04992_),
    .B(_09317_),
    .Y(_02389_));
 sky130_fd_sc_hd__nor2_1 _23273_ (.A(_05167_),
    .B(_09317_),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_1 _23274_ (.A(_05175_),
    .B(_09317_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_1 _23275_ (.A(_05184_),
    .B(_09317_),
    .Y(_02392_));
 sky130_fd_sc_hd__nor2_1 _23276_ (.A(_05196_),
    .B(_09317_),
    .Y(_02393_));
 sky130_fd_sc_hd__nor2_1 _23277_ (.A(_05206_),
    .B(_09317_),
    .Y(_02394_));
 sky130_fd_sc_hd__nor2_1 _23278_ (.A(_05214_),
    .B(_09317_),
    .Y(_02395_));
 sky130_fd_sc_hd__nor2_1 _23279_ (.A(_05224_),
    .B(_09317_),
    .Y(_02396_));
 sky130_fd_sc_hd__nor2_1 _23280_ (.A(_05236_),
    .B(_09317_),
    .Y(_02397_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_660 ();
 sky130_fd_sc_hd__nor2_1 _23282_ (.A(_05243_),
    .B(_09317_),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _23283_ (.A(_05251_),
    .B(_09317_),
    .Y(_02399_));
 sky130_fd_sc_hd__nor2_1 _23284_ (.A(_04995_),
    .B(_09317_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _23285_ (.A(_05260_),
    .B(_09317_),
    .Y(_02401_));
 sky130_fd_sc_hd__nor2_1 _23286_ (.A(_05310_),
    .B(_09317_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_1 _23287_ (.A(_05003_),
    .B(_09317_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _23288_ (.A(_05012_),
    .B(_09317_),
    .Y(_02404_));
 sky130_fd_sc_hd__nor2_1 _23289_ (.A(_05021_),
    .B(_09317_),
    .Y(_02405_));
 sky130_fd_sc_hd__nor2_1 _23290_ (.A(_05032_),
    .B(_09317_),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _23291_ (.A(_05039_),
    .B(_09317_),
    .Y(_02407_));
 sky130_fd_sc_hd__nor2_1 _23292_ (.A(_05048_),
    .B(_09317_),
    .Y(_02408_));
 sky130_fd_sc_hd__nor2_1 _23293_ (.A(_05055_),
    .B(_09317_),
    .Y(_02409_));
 sky130_fd_sc_hd__nand2_8 _23294_ (.A(_09991_),
    .B(_05655_),
    .Y(_09321_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_659 ();
 sky130_fd_sc_hd__nor2_1 _23296_ (.A(_05317_),
    .B(_09321_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor2_1 _23297_ (.A(_05388_),
    .B(_09321_),
    .Y(_02411_));
 sky130_fd_sc_hd__nor2_1 _23298_ (.A(_05402_),
    .B(_09321_),
    .Y(_02412_));
 sky130_fd_sc_hd__nor2_1 _23299_ (.A(_05412_),
    .B(_09321_),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _23300_ (.A(_05419_),
    .B(_09321_),
    .Y(_02414_));
 sky130_fd_sc_hd__nor2_1 _23301_ (.A(_05426_),
    .B(_09321_),
    .Y(_02415_));
 sky130_fd_sc_hd__nor2_1 _23302_ (.A(_05438_),
    .B(_09321_),
    .Y(_02416_));
 sky130_fd_sc_hd__nor2_1 _23303_ (.A(_05447_),
    .B(_09321_),
    .Y(_02417_));
 sky130_fd_sc_hd__nor2_1 _23304_ (.A(_05453_),
    .B(_09321_),
    .Y(_02418_));
 sky130_fd_sc_hd__nor2_1 _23305_ (.A(_05465_),
    .B(_09321_),
    .Y(_02419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_658 ();
 sky130_fd_sc_hd__nor2_1 _23307_ (.A(_05480_),
    .B(_09321_),
    .Y(_02420_));
 sky130_fd_sc_hd__nor2_1 _23308_ (.A(_05321_),
    .B(_09321_),
    .Y(_02421_));
 sky130_fd_sc_hd__nor2_1 _23309_ (.A(_05488_),
    .B(_09321_),
    .Y(_02422_));
 sky130_fd_sc_hd__nor2_1 _23310_ (.A(_05498_),
    .B(_09321_),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_1 _23311_ (.A(_05509_),
    .B(_09321_),
    .Y(_02424_));
 sky130_fd_sc_hd__nor2_1 _23312_ (.A(_05515_),
    .B(_09321_),
    .Y(_02425_));
 sky130_fd_sc_hd__nor2_1 _23313_ (.A(_05523_),
    .B(_09321_),
    .Y(_02426_));
 sky130_fd_sc_hd__nor2_1 _23314_ (.A(_05535_),
    .B(_09321_),
    .Y(_02427_));
 sky130_fd_sc_hd__nor2_1 _23315_ (.A(_05542_),
    .B(_09321_),
    .Y(_02428_));
 sky130_fd_sc_hd__nor2_1 _23316_ (.A(_05551_),
    .B(_09321_),
    .Y(_02429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_657 ();
 sky130_fd_sc_hd__nor2_1 _23318_ (.A(_05559_),
    .B(_09321_),
    .Y(_02430_));
 sky130_fd_sc_hd__nor2_1 _23319_ (.A(_05567_),
    .B(_09321_),
    .Y(_02431_));
 sky130_fd_sc_hd__nor2_1 _23320_ (.A(_05324_),
    .B(_09321_),
    .Y(_02432_));
 sky130_fd_sc_hd__nor2_1 _23321_ (.A(_05573_),
    .B(_09321_),
    .Y(_02433_));
 sky130_fd_sc_hd__nor2_1 _23322_ (.A(_05611_),
    .B(_09321_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_1 _23323_ (.A(_05330_),
    .B(_09321_),
    .Y(_02435_));
 sky130_fd_sc_hd__nor2_1 _23324_ (.A(_05338_),
    .B(_09321_),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _23325_ (.A(_05347_),
    .B(_09321_),
    .Y(_02437_));
 sky130_fd_sc_hd__nor2_1 _23326_ (.A(_05354_),
    .B(_09321_),
    .Y(_02438_));
 sky130_fd_sc_hd__nor2_1 _23327_ (.A(_05360_),
    .B(_09321_),
    .Y(_02439_));
 sky130_fd_sc_hd__nor2_1 _23328_ (.A(_05371_),
    .B(_09321_),
    .Y(_02440_));
 sky130_fd_sc_hd__nor2_1 _23329_ (.A(_05380_),
    .B(_09321_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_8 _23330_ (.A(_09940_),
    .B(_05696_),
    .Y(_09325_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_656 ();
 sky130_fd_sc_hd__nor2_1 _23332_ (.A(_04988_),
    .B(_09325_),
    .Y(_02442_));
 sky130_fd_sc_hd__nor2_1 _23333_ (.A(_05062_),
    .B(_09325_),
    .Y(_02443_));
 sky130_fd_sc_hd__nor2_1 _23334_ (.A(_05077_),
    .B(_09325_),
    .Y(_02444_));
 sky130_fd_sc_hd__nor2_1 _23335_ (.A(_05087_),
    .B(_09325_),
    .Y(_02445_));
 sky130_fd_sc_hd__nor2_1 _23336_ (.A(_05095_),
    .B(_09325_),
    .Y(_02446_));
 sky130_fd_sc_hd__nor2_1 _23337_ (.A(_05102_),
    .B(_09325_),
    .Y(_02447_));
 sky130_fd_sc_hd__nor2_1 _23338_ (.A(_05112_),
    .B(_09325_),
    .Y(_02448_));
 sky130_fd_sc_hd__nor2_1 _23339_ (.A(_05121_),
    .B(_09325_),
    .Y(_02449_));
 sky130_fd_sc_hd__nor2_1 _23340_ (.A(_05128_),
    .B(_09325_),
    .Y(_02450_));
 sky130_fd_sc_hd__nor2_1 _23341_ (.A(_05137_),
    .B(_09325_),
    .Y(_02451_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_655 ();
 sky130_fd_sc_hd__nor2_1 _23343_ (.A(_05154_),
    .B(_09325_),
    .Y(_02452_));
 sky130_fd_sc_hd__nor2_1 _23344_ (.A(_04992_),
    .B(_09325_),
    .Y(_02453_));
 sky130_fd_sc_hd__nor2_1 _23345_ (.A(_05167_),
    .B(_09325_),
    .Y(_02454_));
 sky130_fd_sc_hd__nor2_1 _23346_ (.A(_05175_),
    .B(_09325_),
    .Y(_02455_));
 sky130_fd_sc_hd__nor2_1 _23347_ (.A(_05184_),
    .B(_09325_),
    .Y(_02456_));
 sky130_fd_sc_hd__nor2_1 _23348_ (.A(_05196_),
    .B(_09325_),
    .Y(_02457_));
 sky130_fd_sc_hd__nor2_1 _23349_ (.A(_05206_),
    .B(_09325_),
    .Y(_02458_));
 sky130_fd_sc_hd__nor2_1 _23350_ (.A(_05214_),
    .B(_09325_),
    .Y(_02459_));
 sky130_fd_sc_hd__nor2_1 _23351_ (.A(_05224_),
    .B(_09325_),
    .Y(_02460_));
 sky130_fd_sc_hd__nor2_1 _23352_ (.A(_05236_),
    .B(_09325_),
    .Y(_02461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_654 ();
 sky130_fd_sc_hd__nor2_1 _23354_ (.A(_05243_),
    .B(_09325_),
    .Y(_02462_));
 sky130_fd_sc_hd__nor2_1 _23355_ (.A(_05251_),
    .B(_09325_),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _23356_ (.A(_04995_),
    .B(_09325_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor2_1 _23357_ (.A(_05260_),
    .B(_09325_),
    .Y(_02465_));
 sky130_fd_sc_hd__nor2_1 _23358_ (.A(_05310_),
    .B(_09325_),
    .Y(_02466_));
 sky130_fd_sc_hd__nor2_1 _23359_ (.A(_05003_),
    .B(_09325_),
    .Y(_02467_));
 sky130_fd_sc_hd__nor2_1 _23360_ (.A(_05012_),
    .B(_09325_),
    .Y(_02468_));
 sky130_fd_sc_hd__nor2_1 _23361_ (.A(_05021_),
    .B(_09325_),
    .Y(_02469_));
 sky130_fd_sc_hd__nor2_1 _23362_ (.A(_05032_),
    .B(_09325_),
    .Y(_02470_));
 sky130_fd_sc_hd__nor2_1 _23363_ (.A(_05039_),
    .B(_09325_),
    .Y(_02471_));
 sky130_fd_sc_hd__nor2_1 _23364_ (.A(_05048_),
    .B(_09325_),
    .Y(_02472_));
 sky130_fd_sc_hd__nor2_1 _23365_ (.A(_05055_),
    .B(_09325_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand2_8 _23366_ (.A(_09991_),
    .B(_05737_),
    .Y(_09329_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_653 ();
 sky130_fd_sc_hd__nor2_1 _23368_ (.A(_05317_),
    .B(_09329_),
    .Y(_02474_));
 sky130_fd_sc_hd__nor2_1 _23369_ (.A(_05388_),
    .B(_09329_),
    .Y(_02475_));
 sky130_fd_sc_hd__nor2_1 _23370_ (.A(_05402_),
    .B(_09329_),
    .Y(_02476_));
 sky130_fd_sc_hd__nor2_1 _23371_ (.A(_05412_),
    .B(_09329_),
    .Y(_02477_));
 sky130_fd_sc_hd__nor2_1 _23372_ (.A(_05419_),
    .B(_09329_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_1 _23373_ (.A(_05426_),
    .B(_09329_),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _23374_ (.A(_05438_),
    .B(_09329_),
    .Y(_02480_));
 sky130_fd_sc_hd__nor2_1 _23375_ (.A(_05447_),
    .B(_09329_),
    .Y(_02481_));
 sky130_fd_sc_hd__nor2_1 _23376_ (.A(_05453_),
    .B(_09329_),
    .Y(_02482_));
 sky130_fd_sc_hd__nor2_1 _23377_ (.A(_05465_),
    .B(_09329_),
    .Y(_02483_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_652 ();
 sky130_fd_sc_hd__nor2_1 _23379_ (.A(_05480_),
    .B(_09329_),
    .Y(_02484_));
 sky130_fd_sc_hd__nor2_1 _23380_ (.A(_05321_),
    .B(_09329_),
    .Y(_02485_));
 sky130_fd_sc_hd__nor2_1 _23381_ (.A(_05488_),
    .B(_09329_),
    .Y(_02486_));
 sky130_fd_sc_hd__nor2_1 _23382_ (.A(_05498_),
    .B(_09329_),
    .Y(_02487_));
 sky130_fd_sc_hd__nor2_1 _23383_ (.A(_05509_),
    .B(_09329_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_1 _23384_ (.A(_05515_),
    .B(_09329_),
    .Y(_02489_));
 sky130_fd_sc_hd__nor2_1 _23385_ (.A(_05523_),
    .B(_09329_),
    .Y(_02490_));
 sky130_fd_sc_hd__nor2_1 _23386_ (.A(_05535_),
    .B(_09329_),
    .Y(_02491_));
 sky130_fd_sc_hd__nor2_1 _23387_ (.A(_05542_),
    .B(_09329_),
    .Y(_02492_));
 sky130_fd_sc_hd__nor2_1 _23388_ (.A(_05551_),
    .B(_09329_),
    .Y(_02493_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_651 ();
 sky130_fd_sc_hd__nor2_1 _23390_ (.A(_05559_),
    .B(_09329_),
    .Y(_02494_));
 sky130_fd_sc_hd__nor2_1 _23391_ (.A(_05567_),
    .B(_09329_),
    .Y(_02495_));
 sky130_fd_sc_hd__nor2_1 _23392_ (.A(_05324_),
    .B(_09329_),
    .Y(_02496_));
 sky130_fd_sc_hd__nor2_1 _23393_ (.A(_05573_),
    .B(_09329_),
    .Y(_02497_));
 sky130_fd_sc_hd__nor2_1 _23394_ (.A(_05611_),
    .B(_09329_),
    .Y(_02498_));
 sky130_fd_sc_hd__nor2_1 _23395_ (.A(_05330_),
    .B(_09329_),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_1 _23396_ (.A(_05338_),
    .B(_09329_),
    .Y(_02500_));
 sky130_fd_sc_hd__nor2_1 _23397_ (.A(_05347_),
    .B(_09329_),
    .Y(_02501_));
 sky130_fd_sc_hd__nor2_1 _23398_ (.A(_05354_),
    .B(_09329_),
    .Y(_02502_));
 sky130_fd_sc_hd__nor2_1 _23399_ (.A(_05360_),
    .B(_09329_),
    .Y(_02503_));
 sky130_fd_sc_hd__nor2_1 _23400_ (.A(_05371_),
    .B(_09329_),
    .Y(_02504_));
 sky130_fd_sc_hd__nor2_1 _23401_ (.A(_05380_),
    .B(_09329_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_8 _23402_ (.A(_09940_),
    .B(_05778_),
    .Y(_09333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_650 ();
 sky130_fd_sc_hd__nor2_1 _23404_ (.A(_04988_),
    .B(_09333_),
    .Y(_02506_));
 sky130_fd_sc_hd__nor2_1 _23405_ (.A(_05062_),
    .B(_09333_),
    .Y(_02507_));
 sky130_fd_sc_hd__nor2_1 _23406_ (.A(_05077_),
    .B(_09333_),
    .Y(_02508_));
 sky130_fd_sc_hd__nor2_1 _23407_ (.A(_05087_),
    .B(_09333_),
    .Y(_02509_));
 sky130_fd_sc_hd__nor2_1 _23408_ (.A(_05095_),
    .B(_09333_),
    .Y(_02510_));
 sky130_fd_sc_hd__nor2_1 _23409_ (.A(_05102_),
    .B(_09333_),
    .Y(_02511_));
 sky130_fd_sc_hd__nor2_1 _23410_ (.A(_05112_),
    .B(_09333_),
    .Y(_02512_));
 sky130_fd_sc_hd__nor2_1 _23411_ (.A(_05121_),
    .B(_09333_),
    .Y(_02513_));
 sky130_fd_sc_hd__nor2_1 _23412_ (.A(_05128_),
    .B(_09333_),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _23413_ (.A(_05137_),
    .B(_09333_),
    .Y(_02515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_649 ();
 sky130_fd_sc_hd__nor2_1 _23415_ (.A(_05154_),
    .B(_09333_),
    .Y(_02516_));
 sky130_fd_sc_hd__nor2_1 _23416_ (.A(_04992_),
    .B(_09333_),
    .Y(_02517_));
 sky130_fd_sc_hd__nor2_1 _23417_ (.A(_05167_),
    .B(_09333_),
    .Y(_02518_));
 sky130_fd_sc_hd__nor2_1 _23418_ (.A(_05175_),
    .B(_09333_),
    .Y(_02519_));
 sky130_fd_sc_hd__nor2_1 _23419_ (.A(_05184_),
    .B(_09333_),
    .Y(_02520_));
 sky130_fd_sc_hd__nor2_1 _23420_ (.A(_05196_),
    .B(_09333_),
    .Y(_02521_));
 sky130_fd_sc_hd__nor2_1 _23421_ (.A(_05206_),
    .B(_09333_),
    .Y(_02522_));
 sky130_fd_sc_hd__nor2_1 _23422_ (.A(_05214_),
    .B(_09333_),
    .Y(_02523_));
 sky130_fd_sc_hd__nor2_1 _23423_ (.A(_05224_),
    .B(_09333_),
    .Y(_02524_));
 sky130_fd_sc_hd__nor2_1 _23424_ (.A(_05236_),
    .B(_09333_),
    .Y(_02525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_648 ();
 sky130_fd_sc_hd__nor2_1 _23426_ (.A(_05243_),
    .B(_09333_),
    .Y(_02526_));
 sky130_fd_sc_hd__nor2_1 _23427_ (.A(_05251_),
    .B(_09333_),
    .Y(_02527_));
 sky130_fd_sc_hd__nor2_1 _23428_ (.A(_04995_),
    .B(_09333_),
    .Y(_02528_));
 sky130_fd_sc_hd__nor2_1 _23429_ (.A(_05260_),
    .B(_09333_),
    .Y(_02529_));
 sky130_fd_sc_hd__nor2_1 _23430_ (.A(_05310_),
    .B(_09333_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_1 _23431_ (.A(_05003_),
    .B(_09333_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_1 _23432_ (.A(_05012_),
    .B(_09333_),
    .Y(_02532_));
 sky130_fd_sc_hd__nor2_1 _23433_ (.A(_05021_),
    .B(_09333_),
    .Y(_02533_));
 sky130_fd_sc_hd__nor2_1 _23434_ (.A(_05032_),
    .B(_09333_),
    .Y(_02534_));
 sky130_fd_sc_hd__nor2_1 _23435_ (.A(_05039_),
    .B(_09333_),
    .Y(_02535_));
 sky130_fd_sc_hd__nor2_1 _23436_ (.A(_05048_),
    .B(_09333_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor2_1 _23437_ (.A(_05055_),
    .B(_09333_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2b_4 _23438_ (.A_N(_09889_),
    .B(_09893_),
    .Y(_09337_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_647 ();
 sky130_fd_sc_hd__nor2_1 _23440_ (.A(_05317_),
    .B(_09337_),
    .Y(_02538_));
 sky130_fd_sc_hd__nor2_1 _23441_ (.A(_05388_),
    .B(_09337_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor2_1 _23442_ (.A(_05402_),
    .B(_09337_),
    .Y(_02540_));
 sky130_fd_sc_hd__nor2_1 _23443_ (.A(_05412_),
    .B(_09337_),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _23444_ (.A(_05419_),
    .B(_09337_),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_1 _23445_ (.A(_05426_),
    .B(_09337_),
    .Y(_02543_));
 sky130_fd_sc_hd__nor2_1 _23446_ (.A(_05438_),
    .B(_09337_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _23447_ (.A(_05447_),
    .B(_09337_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _23448_ (.A(_05453_),
    .B(_09337_),
    .Y(_02546_));
 sky130_fd_sc_hd__nor2_1 _23449_ (.A(_05465_),
    .B(_09337_),
    .Y(_02547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_646 ();
 sky130_fd_sc_hd__nor2_1 _23451_ (.A(_05480_),
    .B(_09337_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor2_1 _23452_ (.A(_05321_),
    .B(_09337_),
    .Y(_02549_));
 sky130_fd_sc_hd__nor2_1 _23453_ (.A(_05488_),
    .B(_09337_),
    .Y(_02550_));
 sky130_fd_sc_hd__nor2_1 _23454_ (.A(_05498_),
    .B(_09337_),
    .Y(_02551_));
 sky130_fd_sc_hd__nor2_1 _23455_ (.A(_05509_),
    .B(_09337_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _23456_ (.A(_05515_),
    .B(_09337_),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _23457_ (.A(_05523_),
    .B(_09337_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_1 _23458_ (.A(_05535_),
    .B(_09337_),
    .Y(_02555_));
 sky130_fd_sc_hd__nor2_1 _23459_ (.A(_05542_),
    .B(_09337_),
    .Y(_02556_));
 sky130_fd_sc_hd__nor2_1 _23460_ (.A(_05551_),
    .B(_09337_),
    .Y(_02557_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_645 ();
 sky130_fd_sc_hd__nor2_1 _23462_ (.A(_05559_),
    .B(_09337_),
    .Y(_02558_));
 sky130_fd_sc_hd__nor2_1 _23463_ (.A(_05567_),
    .B(_09337_),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2_1 _23464_ (.A(_05324_),
    .B(_09337_),
    .Y(_02560_));
 sky130_fd_sc_hd__nor2_1 _23465_ (.A(_05573_),
    .B(_09337_),
    .Y(_02561_));
 sky130_fd_sc_hd__nor2_1 _23466_ (.A(_05611_),
    .B(_09337_),
    .Y(_02562_));
 sky130_fd_sc_hd__nor2_1 _23467_ (.A(_05330_),
    .B(_09337_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_1 _23468_ (.A(_05338_),
    .B(_09337_),
    .Y(_02564_));
 sky130_fd_sc_hd__nor2_1 _23469_ (.A(_05347_),
    .B(_09337_),
    .Y(_02565_));
 sky130_fd_sc_hd__nor2_1 _23470_ (.A(_05354_),
    .B(_09337_),
    .Y(_02566_));
 sky130_fd_sc_hd__nor2_1 _23471_ (.A(_05360_),
    .B(_09337_),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_1 _23472_ (.A(_05371_),
    .B(_09337_),
    .Y(_02568_));
 sky130_fd_sc_hd__nor2_1 _23473_ (.A(_05380_),
    .B(_09337_),
    .Y(_02569_));
 sky130_fd_sc_hd__nor2b_2 _23474_ (.A(net520),
    .B_N(\hash.CA2.b_dash[0] ),
    .Y(\hash.CA1.d[0] ));
 sky130_fd_sc_hd__inv_1 _23475_ (.A(_13741_),
    .Y(_09341_));
 sky130_fd_sc_hd__inv_1 _23476_ (.A(_13733_),
    .Y(_09342_));
 sky130_fd_sc_hd__inv_1 _23477_ (.A(_13725_),
    .Y(_09343_));
 sky130_fd_sc_hd__nor2b_1 _23478_ (.A(_13053_),
    .B_N(_13722_),
    .Y(_09344_));
 sky130_fd_sc_hd__o21ai_1 _23479_ (.A1(_13721_),
    .A2(_09344_),
    .B1(_13726_),
    .Y(_09345_));
 sky130_fd_sc_hd__a21boi_2 _23480_ (.A1(_09345_),
    .A2(_09343_),
    .B1_N(_13730_),
    .Y(_09346_));
 sky130_fd_sc_hd__o21ai_2 _23481_ (.A1(_09346_),
    .A2(_13729_),
    .B1(_13734_),
    .Y(_09347_));
 sky130_fd_sc_hd__inv_1 _23482_ (.A(_13738_),
    .Y(_09348_));
 sky130_fd_sc_hd__a21oi_2 _23483_ (.A1(_09347_),
    .A2(_09342_),
    .B1(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__o21ai_2 _23484_ (.A1(_09349_),
    .A2(_13737_),
    .B1(_13742_),
    .Y(_09350_));
 sky130_fd_sc_hd__nand2_1 _23485_ (.A(_13746_),
    .B(_13750_),
    .Y(_09351_));
 sky130_fd_sc_hd__a21oi_4 _23486_ (.A1(_09350_),
    .A2(_09341_),
    .B1(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__a21o_1 _23487_ (.A1(_13750_),
    .A2(_13745_),
    .B1(_13749_),
    .X(_09353_));
 sky130_fd_sc_hd__nor2_1 _23488_ (.A(_09352_),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__xnor2_1 _23489_ (.A(_13754_),
    .B(_09354_),
    .Y(\hash.CA1.p1[10] ));
 sky130_fd_sc_hd__inv_1 _23490_ (.A(_13750_),
    .Y(_09355_));
 sky130_fd_sc_hd__inv_1 _23491_ (.A(_13726_),
    .Y(_09356_));
 sky130_fd_sc_hd__a21o_1 _23492_ (.A1(_14375_),
    .A2(_13718_),
    .B1(_13717_),
    .X(_09357_));
 sky130_fd_sc_hd__a21oi_1 _23493_ (.A1(_13722_),
    .A2(_09357_),
    .B1(_13721_),
    .Y(_09358_));
 sky130_fd_sc_hd__nor2_1 _23494_ (.A(_13725_),
    .B(_13729_),
    .Y(_09359_));
 sky130_fd_sc_hd__o21ai_1 _23495_ (.A1(_09356_),
    .A2(_09358_),
    .B1(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__o21a_1 _23496_ (.A1(_13730_),
    .A2(_13729_),
    .B1(_13734_),
    .X(_09361_));
 sky130_fd_sc_hd__a21oi_2 _23497_ (.A1(_09360_),
    .A2(_09361_),
    .B1(_13733_),
    .Y(_09362_));
 sky130_fd_sc_hd__nand2_1 _23498_ (.A(_13738_),
    .B(_13742_),
    .Y(_09363_));
 sky130_fd_sc_hd__a21oi_1 _23499_ (.A1(_13742_),
    .A2(_13737_),
    .B1(_13741_),
    .Y(_09364_));
 sky130_fd_sc_hd__o21ai_2 _23500_ (.A1(_09362_),
    .A2(_09363_),
    .B1(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__a21oi_4 _23501_ (.A1(_09365_),
    .A2(_13746_),
    .B1(_13745_),
    .Y(_09366_));
 sky130_fd_sc_hd__o21bai_1 _23502_ (.A1(_09355_),
    .A2(_09366_),
    .B1_N(_13749_),
    .Y(_09367_));
 sky130_fd_sc_hd__a21oi_1 _23503_ (.A1(_13754_),
    .A2(_09367_),
    .B1(_13753_),
    .Y(_09368_));
 sky130_fd_sc_hd__xnor2_1 _23504_ (.A(_13758_),
    .B(_09368_),
    .Y(\hash.CA1.p1[11] ));
 sky130_fd_sc_hd__o21ai_0 _23505_ (.A1(_09352_),
    .A2(_09353_),
    .B1(_13754_),
    .Y(_09369_));
 sky130_fd_sc_hd__nand2b_1 _23506_ (.A_N(_13753_),
    .B(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__a21oi_1 _23507_ (.A1(_13758_),
    .A2(_09370_),
    .B1(_13757_),
    .Y(_09371_));
 sky130_fd_sc_hd__xnor2_1 _23508_ (.A(_13762_),
    .B(_09371_),
    .Y(\hash.CA1.p1[12] ));
 sky130_fd_sc_hd__o2111ai_1 _23509_ (.A1(_13758_),
    .A2(_13757_),
    .B1(_13762_),
    .C1(_13750_),
    .D1(_13754_),
    .Y(_09372_));
 sky130_fd_sc_hd__a21o_1 _23510_ (.A1(_13754_),
    .A2(_13749_),
    .B1(_13753_),
    .X(_09373_));
 sky130_fd_sc_hd__a21o_1 _23511_ (.A1(_13758_),
    .A2(_09373_),
    .B1(_13757_),
    .X(_09374_));
 sky130_fd_sc_hd__a21oi_1 _23512_ (.A1(_13762_),
    .A2(_09374_),
    .B1(_13761_),
    .Y(_09375_));
 sky130_fd_sc_hd__o21a_4 _23513_ (.A1(_09372_),
    .A2(_09366_),
    .B1(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__xnor2_1 _23514_ (.A(_13766_),
    .B(_09376_),
    .Y(\hash.CA1.p1[13] ));
 sky130_fd_sc_hd__nand3_2 _23515_ (.A(_13754_),
    .B(_13758_),
    .C(_13762_),
    .Y(_09377_));
 sky130_fd_sc_hd__nor2_1 _23516_ (.A(_09354_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__inv_1 _23517_ (.A(_13766_),
    .Y(_09379_));
 sky130_fd_sc_hd__a21o_1 _23518_ (.A1(_13758_),
    .A2(_13753_),
    .B1(_13757_),
    .X(_09380_));
 sky130_fd_sc_hd__a21oi_1 _23519_ (.A1(_13762_),
    .A2(_09380_),
    .B1(_13761_),
    .Y(_09381_));
 sky130_fd_sc_hd__o21bai_1 _23520_ (.A1(_09379_),
    .A2(_09381_),
    .B1_N(_13765_),
    .Y(_09382_));
 sky130_fd_sc_hd__a21oi_1 _23521_ (.A1(_13766_),
    .A2(_09378_),
    .B1(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__xnor2_1 _23522_ (.A(_13770_),
    .B(_09383_),
    .Y(\hash.CA1.p1[14] ));
 sky130_fd_sc_hd__o21bai_1 _23523_ (.A1(_09379_),
    .A2(_09376_),
    .B1_N(_13765_),
    .Y(_09384_));
 sky130_fd_sc_hd__a21oi_1 _23524_ (.A1(_13770_),
    .A2(_09384_),
    .B1(_13769_),
    .Y(_09385_));
 sky130_fd_sc_hd__xnor2_1 _23525_ (.A(_13774_),
    .B(_09385_),
    .Y(\hash.CA1.p1[15] ));
 sky130_fd_sc_hd__nand3_2 _23526_ (.A(_13766_),
    .B(_13770_),
    .C(_13774_),
    .Y(_09386_));
 sky130_fd_sc_hd__a21o_1 _23527_ (.A1(_13770_),
    .A2(_09382_),
    .B1(_13769_),
    .X(_09387_));
 sky130_fd_sc_hd__a21oi_1 _23528_ (.A1(_13774_),
    .A2(_09387_),
    .B1(_13773_),
    .Y(_09388_));
 sky130_fd_sc_hd__o31ai_2 _23529_ (.A1(_09354_),
    .A2(_09377_),
    .A3(_09386_),
    .B1(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__xor2_1 _23530_ (.A(_13778_),
    .B(_09389_),
    .X(\hash.CA1.p1[16] ));
 sky130_fd_sc_hd__a21o_1 _23531_ (.A1(_13770_),
    .A2(_13765_),
    .B1(_13769_),
    .X(_09390_));
 sky130_fd_sc_hd__a21oi_2 _23532_ (.A1(_13774_),
    .A2(_09390_),
    .B1(_13773_),
    .Y(_09391_));
 sky130_fd_sc_hd__o21ai_1 _23533_ (.A1(_09376_),
    .A2(_09386_),
    .B1(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__a21oi_1 _23534_ (.A1(_13778_),
    .A2(_09392_),
    .B1(_13777_),
    .Y(_09393_));
 sky130_fd_sc_hd__xnor2_1 _23535_ (.A(_13782_),
    .B(_09393_),
    .Y(\hash.CA1.p1[17] ));
 sky130_fd_sc_hd__a21o_1 _23536_ (.A1(_13778_),
    .A2(_09389_),
    .B1(_13777_),
    .X(_09394_));
 sky130_fd_sc_hd__a21oi_1 _23537_ (.A1(_13782_),
    .A2(_09394_),
    .B1(_13781_),
    .Y(_09395_));
 sky130_fd_sc_hd__xnor2_1 _23538_ (.A(_13786_),
    .B(_09395_),
    .Y(\hash.CA1.p1[18] ));
 sky130_fd_sc_hd__and3_1 _23539_ (.A(_13778_),
    .B(_13782_),
    .C(_13786_),
    .X(_09396_));
 sky130_fd_sc_hd__a21o_1 _23540_ (.A1(_13782_),
    .A2(_13777_),
    .B1(_13781_),
    .X(_09397_));
 sky130_fd_sc_hd__a21o_1 _23541_ (.A1(_13786_),
    .A2(_09397_),
    .B1(_13785_),
    .X(_09398_));
 sky130_fd_sc_hd__a21oi_1 _23542_ (.A1(_09392_),
    .A2(_09396_),
    .B1(_09398_),
    .Y(_09399_));
 sky130_fd_sc_hd__xnor2_1 _23543_ (.A(_13790_),
    .B(_09399_),
    .Y(\hash.CA1.p1[19] ));
 sky130_fd_sc_hd__nand3_2 _23544_ (.A(_13778_),
    .B(_13782_),
    .C(_13786_),
    .Y(_09400_));
 sky130_fd_sc_hd__nor2_1 _23545_ (.A(_09388_),
    .B(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__nor2_2 _23546_ (.A(_09398_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__nor3_2 _23547_ (.A(_09377_),
    .B(_09386_),
    .C(_09400_),
    .Y(_09403_));
 sky130_fd_sc_hd__o21ai_4 _23548_ (.A1(_09353_),
    .A2(_09352_),
    .B1(_09403_),
    .Y(_09404_));
 sky130_fd_sc_hd__a21boi_0 _23549_ (.A1(_09402_),
    .A2(_09404_),
    .B1_N(_13790_),
    .Y(_09405_));
 sky130_fd_sc_hd__nor2_1 _23550_ (.A(_13789_),
    .B(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__xnor2_1 _23551_ (.A(_13794_),
    .B(_09406_),
    .Y(\hash.CA1.p1[20] ));
 sky130_fd_sc_hd__nor2_1 _23552_ (.A(_09386_),
    .B(_09400_),
    .Y(_09407_));
 sky130_fd_sc_hd__nand2_1 _23553_ (.A(_13790_),
    .B(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_1 _23554_ (.A(_13790_),
    .B(_09396_),
    .Y(_09409_));
 sky130_fd_sc_hd__a2bb2oi_1 _23555_ (.A1_N(_09391_),
    .A2_N(_09409_),
    .B1(_09398_),
    .B2(_13790_),
    .Y(_09410_));
 sky130_fd_sc_hd__inv_1 _23556_ (.A(_13789_),
    .Y(_09411_));
 sky130_fd_sc_hd__o211ai_1 _23557_ (.A1(_09376_),
    .A2(_09408_),
    .B1(_09410_),
    .C1(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__a21oi_1 _23558_ (.A1(_13794_),
    .A2(_09412_),
    .B1(_13793_),
    .Y(_09413_));
 sky130_fd_sc_hd__xnor2_1 _23559_ (.A(_13798_),
    .B(_09413_),
    .Y(\hash.CA1.p1[21] ));
 sky130_fd_sc_hd__nor3_2 _23560_ (.A(_13789_),
    .B(_13793_),
    .C(_13797_),
    .Y(_09414_));
 sky130_fd_sc_hd__o21ai_0 _23561_ (.A1(_13794_),
    .A2(_13793_),
    .B1(_13798_),
    .Y(_09415_));
 sky130_fd_sc_hd__nand2b_1 _23562_ (.A_N(_13797_),
    .B(_09415_),
    .Y(_09416_));
 sky130_fd_sc_hd__o41ai_2 _23563_ (.A1(_13790_),
    .A2(_13789_),
    .A3(_13793_),
    .A4(_13797_),
    .B1(_09416_),
    .Y(_09417_));
 sky130_fd_sc_hd__a31oi_4 _23564_ (.A1(_09404_),
    .A2(_09402_),
    .A3(_09414_),
    .B1(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__xor2_1 _23565_ (.A(_13802_),
    .B(_09418_),
    .X(\hash.CA1.p1[22] ));
 sky130_fd_sc_hd__o211ai_2 _23566_ (.A1(_09408_),
    .A2(_09376_),
    .B1(_09410_),
    .C1(_09414_),
    .Y(_09419_));
 sky130_fd_sc_hd__a31o_1 _23567_ (.A1(_09416_),
    .A2(_09419_),
    .A3(_13802_),
    .B1(_13801_),
    .X(_09420_));
 sky130_fd_sc_hd__xor2_1 _23568_ (.A(_13806_),
    .B(_09420_),
    .X(\hash.CA1.p1[23] ));
 sky130_fd_sc_hd__a21o_1 _23569_ (.A1(_13802_),
    .A2(_09418_),
    .B1(_13801_),
    .X(_09421_));
 sky130_fd_sc_hd__a21oi_1 _23570_ (.A1(_13806_),
    .A2(_09421_),
    .B1(_13805_),
    .Y(_09422_));
 sky130_fd_sc_hd__xnor2_1 _23571_ (.A(_13810_),
    .B(_09422_),
    .Y(\hash.CA1.p1[24] ));
 sky130_fd_sc_hd__a21o_1 _23572_ (.A1(_13806_),
    .A2(_09420_),
    .B1(_13805_),
    .X(_09423_));
 sky130_fd_sc_hd__a21oi_1 _23573_ (.A1(_13810_),
    .A2(_09423_),
    .B1(_13809_),
    .Y(_09424_));
 sky130_fd_sc_hd__xnor2_1 _23574_ (.A(_13814_),
    .B(_09424_),
    .Y(\hash.CA1.p1[25] ));
 sky130_fd_sc_hd__inv_1 _23575_ (.A(_13809_),
    .Y(_09425_));
 sky130_fd_sc_hd__and3_1 _23576_ (.A(_13802_),
    .B(_13806_),
    .C(_13810_),
    .X(_09426_));
 sky130_fd_sc_hd__nand2_1 _23577_ (.A(_13810_),
    .B(_13805_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand3_1 _23578_ (.A(_13806_),
    .B(_13810_),
    .C(_13801_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand2_1 _23579_ (.A(_09427_),
    .B(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__a21oi_1 _23580_ (.A1(_09418_),
    .A2(_09426_),
    .B1(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__nand2_1 _23581_ (.A(_09425_),
    .B(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__a21oi_1 _23582_ (.A1(_13814_),
    .A2(_09431_),
    .B1(_13813_),
    .Y(_09432_));
 sky130_fd_sc_hd__xnor2_1 _23583_ (.A(_13818_),
    .B(_09432_),
    .Y(\hash.CA1.p1[26] ));
 sky130_fd_sc_hd__nand2_1 _23584_ (.A(_13806_),
    .B(_13810_),
    .Y(_09433_));
 sky130_fd_sc_hd__nand2_1 _23585_ (.A(_13814_),
    .B(_13818_),
    .Y(_09434_));
 sky130_fd_sc_hd__nor2_1 _23586_ (.A(_09433_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__a21oi_1 _23587_ (.A1(_09425_),
    .A2(_09427_),
    .B1(_09434_),
    .Y(_09436_));
 sky130_fd_sc_hd__a21oi_2 _23588_ (.A1(_09420_),
    .A2(_09435_),
    .B1(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__a21oi_2 _23589_ (.A1(_13818_),
    .A2(_13813_),
    .B1(_13817_),
    .Y(_09438_));
 sky130_fd_sc_hd__nand2_1 _23590_ (.A(_09437_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__xor2_1 _23591_ (.A(_13822_),
    .B(_09439_),
    .X(\hash.CA1.p1[27] ));
 sky130_fd_sc_hd__nor2_1 _23592_ (.A(_13809_),
    .B(_13821_),
    .Y(_09440_));
 sky130_fd_sc_hd__nand2_1 _23593_ (.A(_09438_),
    .B(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__a211o_1 _23594_ (.A1(_09426_),
    .A2(_09418_),
    .B1(_09429_),
    .C1(_09441_),
    .X(_09442_));
 sky130_fd_sc_hd__a21oi_1 _23595_ (.A1(_13814_),
    .A2(_13818_),
    .B1(_13821_),
    .Y(_09443_));
 sky130_fd_sc_hd__nor2_1 _23596_ (.A(_13822_),
    .B(_13821_),
    .Y(_09444_));
 sky130_fd_sc_hd__a21oi_1 _23597_ (.A1(_09438_),
    .A2(_09443_),
    .B1(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__nand2_1 _23598_ (.A(_09442_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__xnor2_1 _23599_ (.A(_13826_),
    .B(_09446_),
    .Y(\hash.CA1.p1[28] ));
 sky130_fd_sc_hd__nor2_1 _23600_ (.A(_13821_),
    .B(_13825_),
    .Y(_09447_));
 sky130_fd_sc_hd__nor3_1 _23601_ (.A(_13822_),
    .B(_13821_),
    .C(_13825_),
    .Y(_09448_));
 sky130_fd_sc_hd__nor2_1 _23602_ (.A(_13826_),
    .B(_13825_),
    .Y(_09449_));
 sky130_fd_sc_hd__a311o_1 _23603_ (.A1(_09437_),
    .A2(_09438_),
    .A3(_09447_),
    .B1(_09448_),
    .C1(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__xnor2_1 _23604_ (.A(_13830_),
    .B(_09450_),
    .Y(\hash.CA1.p1[29] ));
 sky130_fd_sc_hd__xnor2_1 _23605_ (.A(_13053_),
    .B(_13722_),
    .Y(\hash.CA1.p1[2] ));
 sky130_fd_sc_hd__a31o_1 _23606_ (.A1(_13826_),
    .A2(_09442_),
    .A3(_09445_),
    .B1(_13825_),
    .X(_09451_));
 sky130_fd_sc_hd__a21oi_2 _23607_ (.A1(_13830_),
    .A2(_09451_),
    .B1(_13829_),
    .Y(_09452_));
 sky130_fd_sc_hd__xnor2_1 _23608_ (.A(_09452_),
    .B(_13834_),
    .Y(\hash.CA1.p1[30] ));
 sky130_fd_sc_hd__xor2_2 _23609_ (.A(_13409_),
    .B(_06337_),
    .X(_09453_));
 sky130_fd_sc_hd__xnor2_4 _23610_ (.A(_06251_),
    .B(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__or4b_1 _23611_ (.A(net521),
    .B(_06460_),
    .C(_09454_),
    .D_N(\hash.CA2.b_dash[31] ),
    .X(_09455_));
 sky130_fd_sc_hd__o32a_1 _23612_ (.A1(net521),
    .A2(_06459_),
    .A3(_09454_),
    .B1(_09455_),
    .B2(_06458_),
    .X(_09456_));
 sky130_fd_sc_hd__nor4_1 _23613_ (.A(net521),
    .B(\hash.CA2.b_dash[31] ),
    .C(_06460_),
    .D(_09454_),
    .Y(_09457_));
 sky130_fd_sc_hd__nand2_1 _23614_ (.A(_06458_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__nor2_2 _23615_ (.A(net521),
    .B(\hash.CA2.b_dash[31] ),
    .Y(_09459_));
 sky130_fd_sc_hd__nand4b_1 _23616_ (.A_N(_06458_),
    .B(_06459_),
    .C(_09454_),
    .D(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__and4_1 _23617_ (.A(net519),
    .B(\hash.CA2.b_dash[31] ),
    .C(_06459_),
    .D(_09454_),
    .X(_09461_));
 sky130_fd_sc_hd__a32oi_1 _23618_ (.A1(net519),
    .A2(_06460_),
    .A3(_09454_),
    .B1(_09461_),
    .B2(_06458_),
    .Y(_09462_));
 sky130_fd_sc_hd__nand4_1 _23619_ (.A(_09456_),
    .B(_09458_),
    .C(_09460_),
    .D(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__nand2_1 _23620_ (.A(_13830_),
    .B(_13834_),
    .Y(_09464_));
 sky130_fd_sc_hd__a21oi_1 _23621_ (.A1(_13834_),
    .A2(_13829_),
    .B1(_13833_),
    .Y(_09465_));
 sky130_fd_sc_hd__o21ai_2 _23622_ (.A1(_09450_),
    .A2(_09464_),
    .B1(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__xnor2_1 _23623_ (.A(_09466_),
    .B(_09463_),
    .Y(\hash.CA1.p1[31] ));
 sky130_fd_sc_hd__xnor2_1 _23624_ (.A(_13726_),
    .B(_09358_),
    .Y(\hash.CA1.p1[3] ));
 sky130_fd_sc_hd__nand2_1 _23625_ (.A(_09343_),
    .B(_09345_),
    .Y(_09467_));
 sky130_fd_sc_hd__nor2_1 _23626_ (.A(_13730_),
    .B(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__nor2_1 _23627_ (.A(_09346_),
    .B(_09468_),
    .Y(\hash.CA1.p1[4] ));
 sky130_fd_sc_hd__o21ai_0 _23628_ (.A1(_09356_),
    .A2(_09358_),
    .B1(_09343_),
    .Y(_09469_));
 sky130_fd_sc_hd__a211oi_1 _23629_ (.A1(_13730_),
    .A2(_09469_),
    .B1(_13729_),
    .C1(_13734_),
    .Y(_09470_));
 sky130_fd_sc_hd__a21oi_1 _23630_ (.A1(_09360_),
    .A2(_09361_),
    .B1(_09470_),
    .Y(\hash.CA1.p1[5] ));
 sky130_fd_sc_hd__and3_1 _23631_ (.A(_09348_),
    .B(_09342_),
    .C(_09347_),
    .X(_09471_));
 sky130_fd_sc_hd__nor2_1 _23632_ (.A(_09349_),
    .B(_09471_),
    .Y(\hash.CA1.p1[6] ));
 sky130_fd_sc_hd__o21bai_1 _23633_ (.A1(_09348_),
    .A2(_09362_),
    .B1_N(_13737_),
    .Y(_09472_));
 sky130_fd_sc_hd__xor2_1 _23634_ (.A(_13742_),
    .B(_09472_),
    .X(\hash.CA1.p1[7] ));
 sky130_fd_sc_hd__nand2_1 _23635_ (.A(_09341_),
    .B(_09350_),
    .Y(_09473_));
 sky130_fd_sc_hd__xor2_1 _23636_ (.A(_13746_),
    .B(_09473_),
    .X(\hash.CA1.p1[8] ));
 sky130_fd_sc_hd__xnor2_1 _23637_ (.A(_13750_),
    .B(_09366_),
    .Y(\hash.CA1.p1[9] ));
 sky130_fd_sc_hd__or3_1 _23638_ (.A(_14313_),
    .B(_14317_),
    .C(_14321_),
    .X(_09474_));
 sky130_fd_sc_hd__inv_1 _23639_ (.A(_14310_),
    .Y(_09475_));
 sky130_fd_sc_hd__a21o_1 _23640_ (.A1(_14378_),
    .A2(_14302_),
    .B1(_14301_),
    .X(_09476_));
 sky130_fd_sc_hd__a21oi_2 _23641_ (.A1(_14306_),
    .A2(_09476_),
    .B1(_14305_),
    .Y(_09477_));
 sky130_fd_sc_hd__inv_1 _23642_ (.A(_14309_),
    .Y(_09478_));
 sky130_fd_sc_hd__o21ai_2 _23643_ (.A1(_09475_),
    .A2(_09477_),
    .B1(_09478_),
    .Y(_09479_));
 sky130_fd_sc_hd__and2_0 _23644_ (.A(_14314_),
    .B(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__nor2_1 _23645_ (.A(_09474_),
    .B(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__o21a_1 _23646_ (.A1(_14318_),
    .A2(_14317_),
    .B1(_14322_),
    .X(_09482_));
 sky130_fd_sc_hd__o21ai_4 _23647_ (.A1(_14321_),
    .A2(_09482_),
    .B1(_14326_),
    .Y(_09483_));
 sky130_fd_sc_hd__o21bai_1 _23648_ (.A1(_09481_),
    .A2(_09483_),
    .B1_N(_14325_),
    .Y(_09484_));
 sky130_fd_sc_hd__a21oi_1 _23649_ (.A1(_14329_),
    .A2(_09484_),
    .B1(_14328_),
    .Y(_09485_));
 sky130_fd_sc_hd__xnor2_1 _23650_ (.A(_14331_),
    .B(_09485_),
    .Y(\hash.CA1.p2[10] ));
 sky130_fd_sc_hd__nand2_4 _23651_ (.A(_14331_),
    .B(_14329_),
    .Y(_09486_));
 sky130_fd_sc_hd__nor2b_1 _23652_ (.A(_13055_),
    .B_N(_14306_),
    .Y(_09487_));
 sky130_fd_sc_hd__o21ai_1 _23653_ (.A1(_14305_),
    .A2(_09487_),
    .B1(_14310_),
    .Y(_09488_));
 sky130_fd_sc_hd__a21boi_2 _23654_ (.A1(_09478_),
    .A2(_09488_),
    .B1_N(_14314_),
    .Y(_09489_));
 sky130_fd_sc_hd__nor2_2 _23655_ (.A(_09474_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__a21o_1 _23656_ (.A1(_14329_),
    .A2(_14325_),
    .B1(_14328_),
    .X(_09491_));
 sky130_fd_sc_hd__a21oi_4 _23657_ (.A1(_14331_),
    .A2(_09491_),
    .B1(_14330_),
    .Y(_09492_));
 sky130_fd_sc_hd__o31ai_1 _23658_ (.A1(_09483_),
    .A2(_09486_),
    .A3(_09490_),
    .B1(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__xor2_1 _23659_ (.A(_14333_),
    .B(_09493_),
    .X(\hash.CA1.p2[11] ));
 sky130_fd_sc_hd__nand2b_1 _23660_ (.A_N(_09474_),
    .B(_09492_),
    .Y(_09494_));
 sky130_fd_sc_hd__a21oi_2 _23661_ (.A1(_14314_),
    .A2(_09479_),
    .B1(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__o21ai_2 _23662_ (.A1(_09486_),
    .A2(_09483_),
    .B1(_09492_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand2_1 _23663_ (.A(_14333_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__o21bai_1 _23664_ (.A1(_09495_),
    .A2(_09497_),
    .B1_N(_14332_),
    .Y(_09498_));
 sky130_fd_sc_hd__xor2_2 _23665_ (.A(_14335_),
    .B(_09498_),
    .X(\hash.CA1.p2[12] ));
 sky130_fd_sc_hd__nand2_1 _23666_ (.A(_14333_),
    .B(_14335_),
    .Y(_09499_));
 sky130_fd_sc_hd__nor2b_1 _23667_ (.A(_09492_),
    .B_N(_14333_),
    .Y(_09500_));
 sky130_fd_sc_hd__o21ai_2 _23668_ (.A1(_14332_),
    .A2(_09500_),
    .B1(_14335_),
    .Y(_09501_));
 sky130_fd_sc_hd__o41ai_4 _23669_ (.A1(_09483_),
    .A2(_09499_),
    .A3(_09490_),
    .A4(_09486_),
    .B1(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__nor2_1 _23670_ (.A(_14334_),
    .B(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__xnor2_1 _23671_ (.A(_14337_),
    .B(_09503_),
    .Y(\hash.CA1.p2[13] ));
 sky130_fd_sc_hd__nand2_1 _23672_ (.A(_14335_),
    .B(_14337_),
    .Y(_09504_));
 sky130_fd_sc_hd__a21o_1 _23673_ (.A1(_14335_),
    .A2(_14332_),
    .B1(_14334_),
    .X(_09505_));
 sky130_fd_sc_hd__nand2_1 _23674_ (.A(_14337_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__o31a_2 _23675_ (.A1(_09495_),
    .A2(_09504_),
    .A3(_09497_),
    .B1(_09506_),
    .X(_09507_));
 sky130_fd_sc_hd__nand2b_1 _23676_ (.A_N(_14336_),
    .B(_09507_),
    .Y(_09508_));
 sky130_fd_sc_hd__xor2_1 _23677_ (.A(_14339_),
    .B(_09508_),
    .X(\hash.CA1.p2[14] ));
 sky130_fd_sc_hd__nor3_1 _23678_ (.A(_14337_),
    .B(_14336_),
    .C(_14338_),
    .Y(_09509_));
 sky130_fd_sc_hd__nor2_1 _23679_ (.A(_14339_),
    .B(_14338_),
    .Y(_09510_));
 sky130_fd_sc_hd__nor2_2 _23680_ (.A(_09509_),
    .B(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__o41ai_4 _23681_ (.A1(_14334_),
    .A2(_14336_),
    .A3(_14338_),
    .A4(_09502_),
    .B1(_09511_),
    .Y(_09512_));
 sky130_fd_sc_hd__xnor2_1 _23682_ (.A(_14341_),
    .B(_09512_),
    .Y(\hash.CA1.p2[15] ));
 sky130_fd_sc_hd__nor3_1 _23683_ (.A(_14336_),
    .B(_14338_),
    .C(_14340_),
    .Y(_09513_));
 sky130_fd_sc_hd__inv_1 _23684_ (.A(_14341_),
    .Y(_09514_));
 sky130_fd_sc_hd__o21ba_1 _23685_ (.A1(_09514_),
    .A2(_09510_),
    .B1_N(_14340_),
    .X(_09515_));
 sky130_fd_sc_hd__a21oi_4 _23686_ (.A1(_09513_),
    .A2(_09507_),
    .B1(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__xor2_1 _23687_ (.A(_14343_),
    .B(_09516_),
    .X(\hash.CA1.p2[16] ));
 sky130_fd_sc_hd__o21bai_1 _23688_ (.A1(_09514_),
    .A2(_09512_),
    .B1_N(_14340_),
    .Y(_09517_));
 sky130_fd_sc_hd__a21oi_1 _23689_ (.A1(_14343_),
    .A2(_09517_),
    .B1(_14342_),
    .Y(_09518_));
 sky130_fd_sc_hd__xnor2_1 _23690_ (.A(_14345_),
    .B(_09518_),
    .Y(\hash.CA1.p2[17] ));
 sky130_fd_sc_hd__a21o_1 _23691_ (.A1(_14343_),
    .A2(_09516_),
    .B1(_14342_),
    .X(_09519_));
 sky130_fd_sc_hd__a21oi_1 _23692_ (.A1(_14345_),
    .A2(_09519_),
    .B1(_14344_),
    .Y(_09520_));
 sky130_fd_sc_hd__xnor2_1 _23693_ (.A(_14347_),
    .B(_09520_),
    .Y(\hash.CA1.p2[18] ));
 sky130_fd_sc_hd__nand3_1 _23694_ (.A(_14341_),
    .B(_14343_),
    .C(_14345_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand2_1 _23695_ (.A(_14345_),
    .B(_14342_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand3_1 _23696_ (.A(_14343_),
    .B(_14345_),
    .C(_14340_),
    .Y(_09523_));
 sky130_fd_sc_hd__o211a_1 _23697_ (.A1(_09512_),
    .A2(_09521_),
    .B1(_09522_),
    .C1(_09523_),
    .X(_09524_));
 sky130_fd_sc_hd__nand2b_1 _23698_ (.A_N(_14344_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__a21oi_1 _23699_ (.A1(_14347_),
    .A2(_09525_),
    .B1(_14346_),
    .Y(_09526_));
 sky130_fd_sc_hd__xnor2_1 _23700_ (.A(_14349_),
    .B(_09526_),
    .Y(\hash.CA1.p2[19] ));
 sky130_fd_sc_hd__o21a_1 _23701_ (.A1(_14343_),
    .A2(_14342_),
    .B1(_14345_),
    .X(_09527_));
 sky130_fd_sc_hd__o211ai_1 _23702_ (.A1(_14344_),
    .A2(_09527_),
    .B1(_14347_),
    .C1(_14349_),
    .Y(_09528_));
 sky130_fd_sc_hd__nand2b_1 _23703_ (.A_N(_14344_),
    .B(_09522_),
    .Y(_09529_));
 sky130_fd_sc_hd__nor2_1 _23704_ (.A(_09516_),
    .B(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__a21oi_1 _23705_ (.A1(_14349_),
    .A2(_14346_),
    .B1(_14348_),
    .Y(_09531_));
 sky130_fd_sc_hd__o21ai_0 _23706_ (.A1(_09528_),
    .A2(_09530_),
    .B1(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__xor2_1 _23707_ (.A(_14351_),
    .B(_09532_),
    .X(\hash.CA1.p2[20] ));
 sky130_fd_sc_hd__nand3_1 _23708_ (.A(_14347_),
    .B(_14349_),
    .C(_14351_),
    .Y(_09533_));
 sky130_fd_sc_hd__a21o_1 _23709_ (.A1(_14347_),
    .A2(_14344_),
    .B1(_14346_),
    .X(_09534_));
 sky130_fd_sc_hd__a21o_1 _23710_ (.A1(_14349_),
    .A2(_09534_),
    .B1(_14348_),
    .X(_09535_));
 sky130_fd_sc_hd__a21oi_2 _23711_ (.A1(_14351_),
    .A2(_09535_),
    .B1(_14350_),
    .Y(_09536_));
 sky130_fd_sc_hd__o21ai_0 _23712_ (.A1(_09524_),
    .A2(_09533_),
    .B1(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__xor2_1 _23713_ (.A(_14353_),
    .B(_09537_),
    .X(\hash.CA1.p2[21] ));
 sky130_fd_sc_hd__nor4b_4 _23714_ (.A(_14350_),
    .B(_09529_),
    .C(_09516_),
    .D_N(_09531_),
    .Y(_09538_));
 sky130_fd_sc_hd__nand3b_1 _23715_ (.A_N(_14350_),
    .B(_09528_),
    .C(_09531_),
    .Y(_09539_));
 sky130_fd_sc_hd__o21ai_1 _23716_ (.A1(_14351_),
    .A2(_14350_),
    .B1(_09539_),
    .Y(_09540_));
 sky130_fd_sc_hd__nor2_1 _23717_ (.A(_09538_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__a21oi_1 _23718_ (.A1(_14353_),
    .A2(_09541_),
    .B1(_14352_),
    .Y(_09542_));
 sky130_fd_sc_hd__xnor2_1 _23719_ (.A(_14355_),
    .B(_09542_),
    .Y(\hash.CA1.p2[22] ));
 sky130_fd_sc_hd__nand2_1 _23720_ (.A(_14353_),
    .B(_14355_),
    .Y(_09543_));
 sky130_fd_sc_hd__nor2_1 _23721_ (.A(_09536_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__a21oi_2 _23722_ (.A1(_14355_),
    .A2(_14352_),
    .B1(_09544_),
    .Y(_09545_));
 sky130_fd_sc_hd__o31ai_1 _23723_ (.A1(_09524_),
    .A2(_09533_),
    .A3(_09543_),
    .B1(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__nor2_1 _23724_ (.A(_14354_),
    .B(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__xnor2_1 _23725_ (.A(_14357_),
    .B(_09547_),
    .Y(\hash.CA1.p2[23] ));
 sky130_fd_sc_hd__or4b_4 _23726_ (.A(_09543_),
    .B(_09540_),
    .C(_09538_),
    .D_N(_14357_),
    .X(_09548_));
 sky130_fd_sc_hd__and3_1 _23727_ (.A(_14355_),
    .B(_14357_),
    .C(_14352_),
    .X(_09549_));
 sky130_fd_sc_hd__a21oi_1 _23728_ (.A1(_14357_),
    .A2(_14354_),
    .B1(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__and3b_1 _23729_ (.A_N(_14356_),
    .B(_09548_),
    .C(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__xnor2_1 _23730_ (.A(_14359_),
    .B(_09551_),
    .Y(\hash.CA1.p2[24] ));
 sky130_fd_sc_hd__nor3_1 _23731_ (.A(_14354_),
    .B(_14356_),
    .C(_14358_),
    .Y(_09552_));
 sky130_fd_sc_hd__o311ai_2 _23732_ (.A1(_09524_),
    .A2(_09533_),
    .A3(_09543_),
    .B1(_09545_),
    .C1(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__or2_0 _23733_ (.A(_14359_),
    .B(_14358_),
    .X(_09554_));
 sky130_fd_sc_hd__o311a_4 _23734_ (.A1(_14357_),
    .A2(_14356_),
    .A3(_14358_),
    .B1(_09554_),
    .C1(_09553_),
    .X(_09555_));
 sky130_fd_sc_hd__xor2_1 _23735_ (.A(_14361_),
    .B(_09555_),
    .X(\hash.CA1.p2[25] ));
 sky130_fd_sc_hd__nor3_1 _23736_ (.A(_14356_),
    .B(_14358_),
    .C(_14360_),
    .Y(_09556_));
 sky130_fd_sc_hd__a21oi_1 _23737_ (.A1(_14361_),
    .A2(_09554_),
    .B1(_14360_),
    .Y(_09557_));
 sky130_fd_sc_hd__a31oi_4 _23738_ (.A1(_09556_),
    .A2(_09550_),
    .A3(_09548_),
    .B1(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__xor2_1 _23739_ (.A(_14363_),
    .B(_09558_),
    .X(\hash.CA1.p2[26] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_644 ();
 sky130_fd_sc_hd__a21o_1 _23741_ (.A1(_09555_),
    .A2(_14361_),
    .B1(_14360_),
    .X(_09560_));
 sky130_fd_sc_hd__a21oi_2 _23742_ (.A1(_09560_),
    .A2(_14363_),
    .B1(_14362_),
    .Y(_09561_));
 sky130_fd_sc_hd__xnor2_1 _23743_ (.A(_14365_),
    .B(_09561_),
    .Y(\hash.CA1.p2[27] ));
 sky130_fd_sc_hd__a21o_1 _23744_ (.A1(_09558_),
    .A2(_14363_),
    .B1(_14362_),
    .X(_09562_));
 sky130_fd_sc_hd__a21oi_2 _23745_ (.A1(_09562_),
    .A2(_14365_),
    .B1(_14364_),
    .Y(_09563_));
 sky130_fd_sc_hd__xnor2_1 _23746_ (.A(_09563_),
    .B(_14367_),
    .Y(\hash.CA1.p2[28] ));
 sky130_fd_sc_hd__nand2_1 _23747_ (.A(_14365_),
    .B(_14362_),
    .Y(_09564_));
 sky130_fd_sc_hd__nand3_1 _23748_ (.A(_14363_),
    .B(_14365_),
    .C(_14360_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand2_1 _23749_ (.A(_09564_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__a41oi_2 _23750_ (.A1(_14361_),
    .A2(_14363_),
    .A3(_14365_),
    .A4(_09555_),
    .B1(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand2b_1 _23751_ (.A_N(_14364_),
    .B(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__a21oi_2 _23752_ (.A1(_09568_),
    .A2(_14367_),
    .B1(_14366_),
    .Y(_09569_));
 sky130_fd_sc_hd__xnor2_1 _23753_ (.A(_09569_),
    .B(_14369_),
    .Y(\hash.CA1.p2[29] ));
 sky130_fd_sc_hd__nand4_1 _23754_ (.A(_09558_),
    .B(_14365_),
    .C(_14367_),
    .D(_14363_),
    .Y(_09570_));
 sky130_fd_sc_hd__nand2_1 _23755_ (.A(_14367_),
    .B(_14364_),
    .Y(_09571_));
 sky130_fd_sc_hd__nand3_1 _23756_ (.A(_14365_),
    .B(_14367_),
    .C(_14362_),
    .Y(_09572_));
 sky130_fd_sc_hd__nand4b_1 _23757_ (.A_N(_14366_),
    .B(_09571_),
    .C(_09570_),
    .D(_09572_),
    .Y(_09573_));
 sky130_fd_sc_hd__a21oi_2 _23758_ (.A1(_09573_),
    .A2(_14369_),
    .B1(_14368_),
    .Y(_09574_));
 sky130_fd_sc_hd__xnor2_1 _23759_ (.A(_14372_),
    .B(_09574_),
    .Y(\hash.CA1.p2[30] ));
 sky130_fd_sc_hd__nand2_1 _23760_ (.A(_14367_),
    .B(_14369_),
    .Y(_09575_));
 sky130_fd_sc_hd__nand2b_1 _23761_ (.A_N(_14366_),
    .B(_09571_),
    .Y(_09576_));
 sky130_fd_sc_hd__a21oi_1 _23762_ (.A1(_14369_),
    .A2(_09576_),
    .B1(_14368_),
    .Y(_09577_));
 sky130_fd_sc_hd__o21ai_1 _23763_ (.A1(_09567_),
    .A2(_09575_),
    .B1(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__a21oi_2 _23764_ (.A1(_09578_),
    .A2(_14372_),
    .B1(_14371_),
    .Y(_09579_));
 sky130_fd_sc_hd__nor2b_1 _23765_ (.A(net522),
    .B_N(\hash.CA2.S1.X[31] ),
    .Y(_09580_));
 sky130_fd_sc_hd__mux2i_2 _23766_ (.A0(_06602_),
    .A1(_09580_),
    .S(_06921_),
    .Y(_09581_));
 sky130_fd_sc_hd__nand2_1 _23767_ (.A(_14295_),
    .B(_07333_),
    .Y(_09582_));
 sky130_fd_sc_hd__a21oi_1 _23768_ (.A1(_14295_),
    .A2(_07338_),
    .B1(_14294_),
    .Y(_09583_));
 sky130_fd_sc_hd__o21ai_1 _23769_ (.A1(_07302_),
    .A2(_09582_),
    .B1(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__nor2_1 _23770_ (.A(net522),
    .B(\hash.CA2.f_dash[31] ),
    .Y(_09585_));
 sky130_fd_sc_hd__mux2i_1 _23771_ (.A0(_06546_),
    .A1(_09585_),
    .S(_06769_),
    .Y(_09586_));
 sky130_fd_sc_hd__xor2_4 _23772_ (.A(\hash.CA1.w_i1[31] ),
    .B(\hash.CA1.k_i1[31] ),
    .X(_09587_));
 sky130_fd_sc_hd__xnor2_1 _23773_ (.A(_06707_),
    .B(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__xnor2_1 _23774_ (.A(_09586_),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__xnor2_1 _23775_ (.A(\hash.CA1.S1.X[24] ),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__xor2_1 _23776_ (.A(_09584_),
    .B(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__a21o_1 _23777_ (.A1(_14272_),
    .A2(_14262_),
    .B1(_14271_),
    .X(_09592_));
 sky130_fd_sc_hd__a21oi_1 _23778_ (.A1(_14282_),
    .A2(_09592_),
    .B1(_14281_),
    .Y(_09593_));
 sky130_fd_sc_hd__nor2_1 _23779_ (.A(_14253_),
    .B(_14290_),
    .Y(_09594_));
 sky130_fd_sc_hd__nand2_1 _23780_ (.A(_09593_),
    .B(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__a31oi_1 _23781_ (.A1(_14263_),
    .A2(_14272_),
    .A3(_14282_),
    .B1(_14290_),
    .Y(_09596_));
 sky130_fd_sc_hd__nand2_1 _23782_ (.A(_09593_),
    .B(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__o221ai_4 _23783_ (.A1(_14291_),
    .A2(_14290_),
    .B1(_07306_),
    .B2(_09595_),
    .C1(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__xnor2_1 _23784_ (.A(_09591_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__xnor2_2 _23785_ (.A(_09581_),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__xnor2_1 _23786_ (.A(_13048_),
    .B(_13044_),
    .Y(_09601_));
 sky130_fd_sc_hd__xnor2_1 _23787_ (.A(_09459_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__xnor2_1 _23788_ (.A(_09600_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__xnor2_1 _23789_ (.A(_09579_),
    .B(_09603_),
    .Y(\hash.CA1.p2[31] ));
 sky130_fd_sc_hd__xnor2_1 _23790_ (.A(_13055_),
    .B(_14306_),
    .Y(\hash.CA1.p2[3] ));
 sky130_fd_sc_hd__xnor2_1 _23791_ (.A(_14310_),
    .B(_09477_),
    .Y(\hash.CA1.p2[4] ));
 sky130_fd_sc_hd__nand2_1 _23792_ (.A(_09478_),
    .B(_09488_),
    .Y(_09604_));
 sky130_fd_sc_hd__nor2_1 _23793_ (.A(_14314_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nor2_1 _23794_ (.A(_09489_),
    .B(_09605_),
    .Y(\hash.CA1.p2[5] ));
 sky130_fd_sc_hd__nor2_1 _23795_ (.A(_14313_),
    .B(_09480_),
    .Y(_09606_));
 sky130_fd_sc_hd__xnor2_1 _23796_ (.A(_14318_),
    .B(_09606_),
    .Y(\hash.CA1.p2[6] ));
 sky130_fd_sc_hd__o21a_1 _23797_ (.A1(_14313_),
    .A2(_09489_),
    .B1(_14318_),
    .X(_09607_));
 sky130_fd_sc_hd__nor2_1 _23798_ (.A(_14317_),
    .B(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__xnor2_1 _23799_ (.A(_14322_),
    .B(_09608_),
    .Y(\hash.CA1.p2[7] ));
 sky130_fd_sc_hd__nor2_1 _23800_ (.A(_14321_),
    .B(_09482_),
    .Y(_09609_));
 sky130_fd_sc_hd__nor2_1 _23801_ (.A(_09481_),
    .B(_09609_),
    .Y(_09610_));
 sky130_fd_sc_hd__xor2_1 _23802_ (.A(_14326_),
    .B(_09610_),
    .X(\hash.CA1.p2[8] ));
 sky130_fd_sc_hd__nor2_1 _23803_ (.A(_09483_),
    .B(_09490_),
    .Y(_09611_));
 sky130_fd_sc_hd__nor2_1 _23804_ (.A(_14325_),
    .B(_09611_),
    .Y(_09612_));
 sky130_fd_sc_hd__xnor2_1 _23805_ (.A(_14329_),
    .B(_09612_),
    .Y(\hash.CA1.p2[9] ));
 sky130_fd_sc_hd__inv_1 _23806_ (.A(_14107_),
    .Y(_09613_));
 sky130_fd_sc_hd__inv_1 _23807_ (.A(_14081_),
    .Y(_09614_));
 sky130_fd_sc_hd__inv_1 _23808_ (.A(_14064_),
    .Y(_09615_));
 sky130_fd_sc_hd__a21o_1 _23809_ (.A1(_14379_),
    .A2(_14045_),
    .B1(_14044_),
    .X(_09616_));
 sky130_fd_sc_hd__a21oi_1 _23810_ (.A1(_14054_),
    .A2(_09616_),
    .B1(_14053_),
    .Y(_09617_));
 sky130_fd_sc_hd__inv_1 _23811_ (.A(_14063_),
    .Y(_09618_));
 sky130_fd_sc_hd__o21ai_1 _23812_ (.A1(_09615_),
    .A2(_09617_),
    .B1(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__a21oi_4 _23813_ (.A1(_14073_),
    .A2(_09619_),
    .B1(_14072_),
    .Y(_09620_));
 sky130_fd_sc_hd__inv_1 _23814_ (.A(_14080_),
    .Y(_09621_));
 sky130_fd_sc_hd__o21ai_1 _23815_ (.A1(_09614_),
    .A2(_09620_),
    .B1(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__a21oi_4 _23816_ (.A1(_14089_),
    .A2(_09622_),
    .B1(_14088_),
    .Y(_09623_));
 sky130_fd_sc_hd__nor2b_1 _23817_ (.A(_09623_),
    .B_N(_14098_),
    .Y(_09624_));
 sky130_fd_sc_hd__nor2_1 _23818_ (.A(_14097_),
    .B(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__nor2_1 _23819_ (.A(_09613_),
    .B(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__nor2_1 _23820_ (.A(_14106_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__xnor2_2 _23821_ (.A(_14116_),
    .B(_09627_),
    .Y(\hash.CA1.p3[10] ));
 sky130_fd_sc_hd__nor2b_1 _23822_ (.A(_13062_),
    .B_N(_14054_),
    .Y(_09628_));
 sky130_fd_sc_hd__o21ai_1 _23823_ (.A1(_14053_),
    .A2(_09628_),
    .B1(_14064_),
    .Y(_09629_));
 sky130_fd_sc_hd__a21boi_2 _23824_ (.A1(_09618_),
    .A2(_09629_),
    .B1_N(_14073_),
    .Y(_09630_));
 sky130_fd_sc_hd__o211ai_4 _23825_ (.A1(_14072_),
    .A2(_09630_),
    .B1(_14081_),
    .C1(_14089_),
    .Y(_09631_));
 sky130_fd_sc_hd__a21oi_2 _23826_ (.A1(_14089_),
    .A2(_14080_),
    .B1(_14088_),
    .Y(_09632_));
 sky130_fd_sc_hd__nand2_1 _23827_ (.A(_09631_),
    .B(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__a21oi_1 _23828_ (.A1(_14098_),
    .A2(_09633_),
    .B1(_14097_),
    .Y(_09634_));
 sky130_fd_sc_hd__o21bai_1 _23829_ (.A1(_09613_),
    .A2(_09634_),
    .B1_N(_14106_),
    .Y(_09635_));
 sky130_fd_sc_hd__a21oi_1 _23830_ (.A1(_14116_),
    .A2(_09635_),
    .B1(_14115_),
    .Y(_09636_));
 sky130_fd_sc_hd__xnor2_1 _23831_ (.A(_14126_),
    .B(_09636_),
    .Y(\hash.CA1.p3[11] ));
 sky130_fd_sc_hd__o21ai_0 _23832_ (.A1(_14106_),
    .A2(_09626_),
    .B1(_14116_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand2b_1 _23833_ (.A_N(_14115_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__a21oi_1 _23834_ (.A1(_14126_),
    .A2(_09638_),
    .B1(_14125_),
    .Y(_09639_));
 sky130_fd_sc_hd__xnor2_2 _23835_ (.A(_14135_),
    .B(_09639_),
    .Y(\hash.CA1.p3[12] ));
 sky130_fd_sc_hd__a21o_1 _23836_ (.A1(_14107_),
    .A2(_14097_),
    .B1(_14106_),
    .X(_09640_));
 sky130_fd_sc_hd__a21o_1 _23837_ (.A1(_14116_),
    .A2(_09640_),
    .B1(_14115_),
    .X(_09641_));
 sky130_fd_sc_hd__a21oi_4 _23838_ (.A1(_14126_),
    .A2(_09641_),
    .B1(_14125_),
    .Y(_09642_));
 sky130_fd_sc_hd__nand4_4 _23839_ (.A(_14116_),
    .B(_14126_),
    .C(_14098_),
    .D(_14107_),
    .Y(_09643_));
 sky130_fd_sc_hd__nand2b_1 _23840_ (.A_N(_09643_),
    .B(_09633_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand2_1 _23841_ (.A(_09642_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__a21oi_1 _23842_ (.A1(_14135_),
    .A2(_09645_),
    .B1(_14134_),
    .Y(_09646_));
 sky130_fd_sc_hd__xnor2_2 _23843_ (.A(_14143_),
    .B(_09646_),
    .Y(\hash.CA1.p3[13] ));
 sky130_fd_sc_hd__o21ai_0 _23844_ (.A1(_14135_),
    .A2(_14134_),
    .B1(_14143_),
    .Y(_09647_));
 sky130_fd_sc_hd__nand2b_1 _23845_ (.A_N(_14142_),
    .B(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__a21oi_1 _23846_ (.A1(_14143_),
    .A2(_14134_),
    .B1(_14142_),
    .Y(_09649_));
 sky130_fd_sc_hd__o211ai_1 _23847_ (.A1(_09623_),
    .A2(_09643_),
    .B1(_09649_),
    .C1(_09642_),
    .Y(_09650_));
 sky130_fd_sc_hd__nand2_1 _23848_ (.A(_09648_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__xnor2_1 _23849_ (.A(_14152_),
    .B(_09651_),
    .Y(\hash.CA1.p3[14] ));
 sky130_fd_sc_hd__o21ai_0 _23850_ (.A1(_14143_),
    .A2(_14142_),
    .B1(_14152_),
    .Y(_09652_));
 sky130_fd_sc_hd__nand2b_1 _23851_ (.A_N(_14151_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__nor3_4 _23852_ (.A(_14134_),
    .B(_14142_),
    .C(_14151_),
    .Y(_09654_));
 sky130_fd_sc_hd__nand4_4 _23853_ (.A(_09654_),
    .B(_09632_),
    .C(_09642_),
    .D(_09631_),
    .Y(_09655_));
 sky130_fd_sc_hd__nor4_2 _23854_ (.A(_14135_),
    .B(_14134_),
    .C(_14142_),
    .D(_14151_),
    .Y(_09656_));
 sky130_fd_sc_hd__a31oi_4 _23855_ (.A1(_09642_),
    .A2(_09643_),
    .A3(_09654_),
    .B1(_09656_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand3_4 _23856_ (.A(_09653_),
    .B(_09655_),
    .C(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__xnor2_2 _23857_ (.A(_14162_),
    .B(_09658_),
    .Y(\hash.CA1.p3[15] ));
 sky130_fd_sc_hd__inv_1 _23858_ (.A(_14088_),
    .Y(_09659_));
 sky130_fd_sc_hd__o211ai_4 _23859_ (.A1(_09614_),
    .A2(_09620_),
    .B1(_09659_),
    .C1(_09621_),
    .Y(_09660_));
 sky130_fd_sc_hd__nor2_2 _23860_ (.A(_14089_),
    .B(_14088_),
    .Y(_09661_));
 sky130_fd_sc_hd__nor2_1 _23861_ (.A(_09643_),
    .B(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__and3_2 _23862_ (.A(_14152_),
    .B(_09648_),
    .C(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__nand2_1 _23863_ (.A(_14152_),
    .B(_09648_),
    .Y(_09664_));
 sky130_fd_sc_hd__a21oi_2 _23864_ (.A1(_09642_),
    .A2(_09649_),
    .B1(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__a211o_1 _23865_ (.A1(_09660_),
    .A2(_09663_),
    .B1(_09665_),
    .C1(_14151_),
    .X(_09666_));
 sky130_fd_sc_hd__a21oi_1 _23866_ (.A1(_14162_),
    .A2(_09666_),
    .B1(_14161_),
    .Y(_09667_));
 sky130_fd_sc_hd__xnor2_1 _23867_ (.A(_14171_),
    .B(_09667_),
    .Y(\hash.CA1.p3[16] ));
 sky130_fd_sc_hd__inv_1 _23868_ (.A(_14162_),
    .Y(_09668_));
 sky130_fd_sc_hd__o21bai_4 _23869_ (.A1(_09668_),
    .A2(_09658_),
    .B1_N(_14161_),
    .Y(_09669_));
 sky130_fd_sc_hd__a21oi_2 _23870_ (.A1(_14171_),
    .A2(_09669_),
    .B1(_14170_),
    .Y(_09670_));
 sky130_fd_sc_hd__xnor2_1 _23871_ (.A(_14179_),
    .B(_09670_),
    .Y(\hash.CA1.p3[17] ));
 sky130_fd_sc_hd__inv_1 _23872_ (.A(_14179_),
    .Y(_09671_));
 sky130_fd_sc_hd__or3_4 _23873_ (.A(_14161_),
    .B(_14151_),
    .C(_14170_),
    .X(_09672_));
 sky130_fd_sc_hd__a211oi_4 _23874_ (.A1(_09660_),
    .A2(_09663_),
    .B1(_09672_),
    .C1(_09665_),
    .Y(_09673_));
 sky130_fd_sc_hd__or2_0 _23875_ (.A(_14162_),
    .B(_14161_),
    .X(_09674_));
 sky130_fd_sc_hd__a21oi_1 _23876_ (.A1(_14171_),
    .A2(_09674_),
    .B1(_14170_),
    .Y(_09675_));
 sky130_fd_sc_hd__nor3_1 _23877_ (.A(_09671_),
    .B(_09673_),
    .C(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__nor2_1 _23878_ (.A(_14178_),
    .B(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__xnor2_1 _23879_ (.A(_14187_),
    .B(_09677_),
    .Y(\hash.CA1.p3[18] ));
 sky130_fd_sc_hd__o21bai_1 _23880_ (.A1(_09671_),
    .A2(_09670_),
    .B1_N(_14178_),
    .Y(_09678_));
 sky130_fd_sc_hd__a21oi_1 _23881_ (.A1(_09678_),
    .A2(_14187_),
    .B1(_14186_),
    .Y(_09679_));
 sky130_fd_sc_hd__xnor2_1 _23882_ (.A(_14195_),
    .B(_09679_),
    .Y(\hash.CA1.p3[19] ));
 sky130_fd_sc_hd__nand3_1 _23883_ (.A(_14179_),
    .B(_14187_),
    .C(_14195_),
    .Y(_09680_));
 sky130_fd_sc_hd__nor3_2 _23884_ (.A(_09680_),
    .B(_09675_),
    .C(_09673_),
    .Y(_09681_));
 sky130_fd_sc_hd__and3_1 _23885_ (.A(_14187_),
    .B(_14195_),
    .C(_14178_),
    .X(_09682_));
 sky130_fd_sc_hd__a2111oi_4 _23886_ (.A1(_14195_),
    .A2(_14186_),
    .B1(_14194_),
    .C1(_09681_),
    .D1(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__xnor2_1 _23887_ (.A(_14203_),
    .B(_09683_),
    .Y(\hash.CA1.p3[20] ));
 sky130_fd_sc_hd__inv_1 _23888_ (.A(_14171_),
    .Y(_09684_));
 sky130_fd_sc_hd__o21a_1 _23889_ (.A1(_14179_),
    .A2(_14178_),
    .B1(_14187_),
    .X(_09685_));
 sky130_fd_sc_hd__o211ai_2 _23890_ (.A1(_09685_),
    .A2(_14186_),
    .B1(_14195_),
    .C1(_14203_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand3_2 _23891_ (.A(_14162_),
    .B(_14212_),
    .C(_09653_),
    .Y(_09687_));
 sky130_fd_sc_hd__nor3_1 _23892_ (.A(_09684_),
    .B(_09687_),
    .C(_09686_),
    .Y(_09688_));
 sky130_fd_sc_hd__a2111oi_4 _23893_ (.A1(_14171_),
    .A2(_14161_),
    .B1(_14170_),
    .C1(_14178_),
    .D1(_14186_),
    .Y(_09689_));
 sky130_fd_sc_hd__a21oi_2 _23894_ (.A1(_14203_),
    .A2(_14194_),
    .B1(_14202_),
    .Y(_09690_));
 sky130_fd_sc_hd__o21ai_2 _23895_ (.A1(_09689_),
    .A2(_09686_),
    .B1(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__a32o_2 _23896_ (.A1(_09688_),
    .A2(_09657_),
    .A3(_09655_),
    .B1(_09691_),
    .B2(_14212_),
    .X(_09692_));
 sky130_fd_sc_hd__nor4_1 _23897_ (.A(_09668_),
    .B(_09684_),
    .C(_09658_),
    .D(_09686_),
    .Y(_09693_));
 sky130_fd_sc_hd__nor3_1 _23898_ (.A(_14212_),
    .B(_09691_),
    .C(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__nor2_1 _23899_ (.A(_09692_),
    .B(_09694_),
    .Y(\hash.CA1.p3[21] ));
 sky130_fd_sc_hd__inv_1 _23900_ (.A(_14203_),
    .Y(_09695_));
 sky130_fd_sc_hd__o21bai_4 _23901_ (.A1(_09695_),
    .A2(_09683_),
    .B1_N(_14202_),
    .Y(_09696_));
 sky130_fd_sc_hd__a21oi_2 _23902_ (.A1(_09696_),
    .A2(_14212_),
    .B1(_14211_),
    .Y(_09697_));
 sky130_fd_sc_hd__xnor2_1 _23903_ (.A(_14222_),
    .B(_09697_),
    .Y(\hash.CA1.p3[22] ));
 sky130_fd_sc_hd__inv_1 _23904_ (.A(_14222_),
    .Y(_09698_));
 sky130_fd_sc_hd__nor2_1 _23905_ (.A(_14211_),
    .B(_09692_),
    .Y(_09699_));
 sky130_fd_sc_hd__nor2_1 _23906_ (.A(_09698_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__nor2_1 _23907_ (.A(_14221_),
    .B(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__xnor2_1 _23908_ (.A(_14232_),
    .B(_09701_),
    .Y(\hash.CA1.p3[23] ));
 sky130_fd_sc_hd__o21bai_1 _23909_ (.A1(_09698_),
    .A2(_09697_),
    .B1_N(_14221_),
    .Y(_09702_));
 sky130_fd_sc_hd__a21oi_1 _23910_ (.A1(_09702_),
    .A2(_14232_),
    .B1(_14231_),
    .Y(_09703_));
 sky130_fd_sc_hd__xnor2_1 _23911_ (.A(_09703_),
    .B(_14242_),
    .Y(\hash.CA1.p3[24] ));
 sky130_fd_sc_hd__or4_4 _23912_ (.A(_14211_),
    .B(_14221_),
    .C(_14231_),
    .D(_09692_),
    .X(_09704_));
 sky130_fd_sc_hd__nor2_1 _23913_ (.A(_14232_),
    .B(_14231_),
    .Y(_09705_));
 sky130_fd_sc_hd__nor3_1 _23914_ (.A(_14222_),
    .B(_14221_),
    .C(_14231_),
    .Y(_09706_));
 sky130_fd_sc_hd__nor2_1 _23915_ (.A(_09705_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__a31oi_1 _23916_ (.A1(_14242_),
    .A2(_09704_),
    .A3(_09707_),
    .B1(_14241_),
    .Y(_09708_));
 sky130_fd_sc_hd__xnor2_1 _23917_ (.A(_14252_),
    .B(_09708_),
    .Y(\hash.CA1.p3[25] ));
 sky130_fd_sc_hd__and3_1 _23918_ (.A(_14212_),
    .B(_14222_),
    .C(_14242_),
    .X(_09709_));
 sky130_fd_sc_hd__nand4_4 _23919_ (.A(_14232_),
    .B(_14252_),
    .C(_09696_),
    .D(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__a21oi_1 _23920_ (.A1(_14222_),
    .A2(_14211_),
    .B1(_14221_),
    .Y(_09711_));
 sky130_fd_sc_hd__nor2b_2 _23921_ (.A(_09711_),
    .B_N(_14232_),
    .Y(_09712_));
 sky130_fd_sc_hd__o21ai_1 _23922_ (.A1(_09712_),
    .A2(_14231_),
    .B1(_14242_),
    .Y(_09713_));
 sky130_fd_sc_hd__nand2b_1 _23923_ (.A_N(_14241_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__a21oi_4 _23924_ (.A1(_09714_),
    .A2(_14252_),
    .B1(_14251_),
    .Y(_09715_));
 sky130_fd_sc_hd__nand2_2 _23925_ (.A(_09710_),
    .B(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__xor2_1 _23926_ (.A(_14261_),
    .B(_09716_),
    .X(\hash.CA1.p3[26] ));
 sky130_fd_sc_hd__a311oi_2 _23927_ (.A1(_14242_),
    .A2(_09704_),
    .A3(_09707_),
    .B1(_14241_),
    .C1(_14251_),
    .Y(_09717_));
 sky130_fd_sc_hd__o21ai_0 _23928_ (.A1(_14252_),
    .A2(_14251_),
    .B1(_14261_),
    .Y(_09718_));
 sky130_fd_sc_hd__nor2_2 _23929_ (.A(_09718_),
    .B(_09717_),
    .Y(_09719_));
 sky130_fd_sc_hd__nor2_1 _23930_ (.A(_09719_),
    .B(_14260_),
    .Y(_09720_));
 sky130_fd_sc_hd__xnor2_1 _23931_ (.A(_14270_),
    .B(_09720_),
    .Y(\hash.CA1.p3[27] ));
 sky130_fd_sc_hd__inv_1 _23932_ (.A(_14280_),
    .Y(_09721_));
 sky130_fd_sc_hd__nor2_1 _23933_ (.A(_14260_),
    .B(_14269_),
    .Y(_09722_));
 sky130_fd_sc_hd__nor3_1 _23934_ (.A(_14261_),
    .B(_14260_),
    .C(_14269_),
    .Y(_09723_));
 sky130_fd_sc_hd__nor2_1 _23935_ (.A(_14270_),
    .B(_14269_),
    .Y(_09724_));
 sky130_fd_sc_hd__a311oi_4 _23936_ (.A1(_09715_),
    .A2(_09710_),
    .A3(_09722_),
    .B1(_09723_),
    .C1(_09724_),
    .Y(_09725_));
 sky130_fd_sc_hd__xnor2_1 _23937_ (.A(_09721_),
    .B(_09725_),
    .Y(\hash.CA1.p3[28] ));
 sky130_fd_sc_hd__or3_1 _23938_ (.A(_14260_),
    .B(_14269_),
    .C(_14279_),
    .X(_09726_));
 sky130_fd_sc_hd__o21bai_1 _23939_ (.A1(_09721_),
    .A2(_09724_),
    .B1_N(_14279_),
    .Y(_09727_));
 sky130_fd_sc_hd__o21ai_1 _23940_ (.A1(_09719_),
    .A2(_09726_),
    .B1(_09727_),
    .Y(_09728_));
 sky130_fd_sc_hd__xnor2_1 _23941_ (.A(_09728_),
    .B(_14289_),
    .Y(\hash.CA1.p3[29] ));
 sky130_fd_sc_hd__nand4b_1 _23942_ (.A_N(_14298_),
    .B(_09725_),
    .C(_14280_),
    .D(_14289_),
    .Y(_09729_));
 sky130_fd_sc_hd__or4b_4 _23943_ (.A(_09725_),
    .B(_14288_),
    .C(_14279_),
    .D_N(_14298_),
    .X(_09730_));
 sky130_fd_sc_hd__nor2_1 _23944_ (.A(_14279_),
    .B(_14288_),
    .Y(_09731_));
 sky130_fd_sc_hd__nor3b_1 _23945_ (.A(_14289_),
    .B(_14288_),
    .C_N(_14298_),
    .Y(_09732_));
 sky130_fd_sc_hd__inv_1 _23946_ (.A(_14288_),
    .Y(_09733_));
 sky130_fd_sc_hd__nand3b_1 _23947_ (.A_N(_14298_),
    .B(_14279_),
    .C(_14289_),
    .Y(_09734_));
 sky130_fd_sc_hd__o21ai_0 _23948_ (.A1(_14298_),
    .A2(_09733_),
    .B1(_09734_),
    .Y(_09735_));
 sky130_fd_sc_hd__a311oi_1 _23949_ (.A1(_09721_),
    .A2(_14298_),
    .A3(_09731_),
    .B1(_09732_),
    .C1(_09735_),
    .Y(_09736_));
 sky130_fd_sc_hd__nand3_2 _23950_ (.A(_09730_),
    .B(_09729_),
    .C(_09736_),
    .Y(\hash.CA1.p3[30] ));
 sky130_fd_sc_hd__o211a_1 _23951_ (.A1(_09726_),
    .A2(_09719_),
    .B1(_09727_),
    .C1(_14289_),
    .X(_09737_));
 sky130_fd_sc_hd__nor2b_1 _23952_ (.A(_12822_),
    .B_N(_14298_),
    .Y(_09738_));
 sky130_fd_sc_hd__nor4b_2 _23953_ (.A(_14288_),
    .B(_14297_),
    .C(_09737_),
    .D_N(_12822_),
    .Y(_09739_));
 sky130_fd_sc_hd__a21oi_1 _23954_ (.A1(_14298_),
    .A2(_14288_),
    .B1(_14297_),
    .Y(_09740_));
 sky130_fd_sc_hd__nor2_1 _23955_ (.A(_14298_),
    .B(_14297_),
    .Y(_09741_));
 sky130_fd_sc_hd__nand2_1 _23956_ (.A(_12822_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__o21ai_0 _23957_ (.A1(_12822_),
    .A2(_09740_),
    .B1(_09742_),
    .Y(_09743_));
 sky130_fd_sc_hd__a211oi_2 _23958_ (.A1(_09737_),
    .A2(_09738_),
    .B1(_09743_),
    .C1(_09739_),
    .Y(_09744_));
 sky130_fd_sc_hd__xnor2_1 _23959_ (.A(_09600_),
    .B(_09744_),
    .Y(\hash.CA1.p3[31] ));
 sky130_fd_sc_hd__xnor2_1 _23960_ (.A(_13062_),
    .B(_14054_),
    .Y(\hash.CA1.p3[3] ));
 sky130_fd_sc_hd__xnor2_1 _23961_ (.A(_14064_),
    .B(_09617_),
    .Y(\hash.CA1.p3[4] ));
 sky130_fd_sc_hd__nand2_1 _23962_ (.A(_09618_),
    .B(_09629_),
    .Y(_09745_));
 sky130_fd_sc_hd__nor2_1 _23963_ (.A(_14073_),
    .B(_09745_),
    .Y(_09746_));
 sky130_fd_sc_hd__nor2_1 _23964_ (.A(_09630_),
    .B(_09746_),
    .Y(\hash.CA1.p3[5] ));
 sky130_fd_sc_hd__xnor2_2 _23965_ (.A(_14081_),
    .B(_09620_),
    .Y(\hash.CA1.p3[6] ));
 sky130_fd_sc_hd__o21ai_0 _23966_ (.A1(_14072_),
    .A2(_09630_),
    .B1(_14081_),
    .Y(_09747_));
 sky130_fd_sc_hd__nand2_1 _23967_ (.A(_09621_),
    .B(_09747_),
    .Y(_09748_));
 sky130_fd_sc_hd__xor2_2 _23968_ (.A(_14089_),
    .B(_09748_),
    .X(\hash.CA1.p3[7] ));
 sky130_fd_sc_hd__xnor2_2 _23969_ (.A(_14098_),
    .B(_09623_),
    .Y(\hash.CA1.p3[8] ));
 sky130_fd_sc_hd__xnor2_2 _23970_ (.A(_14107_),
    .B(_09634_),
    .Y(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__inv_1 _23971_ (.A(_08256_),
    .Y(_09749_));
 sky130_fd_sc_hd__o211ai_2 _23972_ (.A1(_08219_),
    .A2(_08241_),
    .B1(_08243_),
    .C1(_08255_),
    .Y(_09750_));
 sky130_fd_sc_hd__a31oi_4 _23973_ (.A1(_14012_),
    .A2(_09749_),
    .A3(_09750_),
    .B1(_14011_),
    .Y(_09751_));
 sky130_fd_sc_hd__xor2_1 _23974_ (.A(\hash.CA1.k_i2[31] ),
    .B(_12666_),
    .X(_09752_));
 sky130_fd_sc_hd__xnor2_1 _23975_ (.A(_06602_),
    .B(_09752_),
    .Y(_09753_));
 sky130_fd_sc_hd__xnor2_2 _23976_ (.A(\hash.CA1.w_i2[31] ),
    .B(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__xnor2_4 _23977_ (.A(_09751_),
    .B(_09754_),
    .Y(\hash.CA1.p4[31] ));
 sky130_fd_sc_hd__a21o_1 _23978_ (.A1(_13880_),
    .A2(_13872_),
    .B1(_13879_),
    .X(_09755_));
 sky130_fd_sc_hd__a21oi_1 _23979_ (.A1(_13886_),
    .A2(_09755_),
    .B1(_13885_),
    .Y(_09756_));
 sky130_fd_sc_hd__inv_1 _23980_ (.A(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__nor2b_1 _23981_ (.A(_13065_),
    .B_N(_13843_),
    .Y(_09758_));
 sky130_fd_sc_hd__o21a_1 _23982_ (.A1(_13842_),
    .A2(_09758_),
    .B1(_13849_),
    .X(_09759_));
 sky130_fd_sc_hd__o21ai_1 _23983_ (.A1(_13848_),
    .A2(_09759_),
    .B1(_13855_),
    .Y(_09760_));
 sky130_fd_sc_hd__nor3_1 _23984_ (.A(_13854_),
    .B(_13860_),
    .C(_13866_),
    .Y(_09761_));
 sky130_fd_sc_hd__o21a_1 _23985_ (.A1(_13861_),
    .A2(_13860_),
    .B1(_13867_),
    .X(_09762_));
 sky130_fd_sc_hd__o21a_1 _23986_ (.A1(_13866_),
    .A2(_09762_),
    .B1(_13873_),
    .X(_09763_));
 sky130_fd_sc_hd__nand3_1 _23987_ (.A(_13880_),
    .B(_13886_),
    .C(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__a21oi_1 _23988_ (.A1(_09760_),
    .A2(_09761_),
    .B1(_09764_),
    .Y(_09765_));
 sky130_fd_sc_hd__nor2_1 _23989_ (.A(_09757_),
    .B(_09765_),
    .Y(_09766_));
 sky130_fd_sc_hd__xnor2_1 _23990_ (.A(_13891_),
    .B(_09766_),
    .Y(\hash.CA1.p5[10] ));
 sky130_fd_sc_hd__inv_1 _23991_ (.A(_13849_),
    .Y(_09767_));
 sky130_fd_sc_hd__a21o_1 _23992_ (.A1(_13066_),
    .A2(_13838_),
    .B1(_13837_),
    .X(_09768_));
 sky130_fd_sc_hd__a21oi_1 _23993_ (.A1(_13843_),
    .A2(_09768_),
    .B1(_13842_),
    .Y(_09769_));
 sky130_fd_sc_hd__o21bai_1 _23994_ (.A1(_09767_),
    .A2(_09769_),
    .B1_N(_13848_),
    .Y(_09770_));
 sky130_fd_sc_hd__a21boi_2 _23995_ (.A1(_13855_),
    .A2(_09770_),
    .B1_N(_09761_),
    .Y(_09771_));
 sky130_fd_sc_hd__o21ai_0 _23996_ (.A1(_09764_),
    .A2(_09771_),
    .B1(_09756_),
    .Y(_09772_));
 sky130_fd_sc_hd__a21oi_1 _23997_ (.A1(_13891_),
    .A2(_09772_),
    .B1(_13890_),
    .Y(_09773_));
 sky130_fd_sc_hd__xnor2_1 _23998_ (.A(_13897_),
    .B(_09773_),
    .Y(\hash.CA1.p5[11] ));
 sky130_fd_sc_hd__inv_1 _23999_ (.A(_13890_),
    .Y(_09774_));
 sky130_fd_sc_hd__o21ai_1 _24000_ (.A1(_09757_),
    .A2(_09765_),
    .B1(_13891_),
    .Y(_09775_));
 sky130_fd_sc_hd__nand2_1 _24001_ (.A(_09774_),
    .B(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__a21oi_1 _24002_ (.A1(_13897_),
    .A2(_09776_),
    .B1(_13896_),
    .Y(_09777_));
 sky130_fd_sc_hd__xnor2_1 _24003_ (.A(_13904_),
    .B(_09777_),
    .Y(\hash.CA1.p5[12] ));
 sky130_fd_sc_hd__nand2_1 _24004_ (.A(_13891_),
    .B(_13897_),
    .Y(_09778_));
 sky130_fd_sc_hd__nor2_1 _24005_ (.A(_09756_),
    .B(_09778_),
    .Y(_09779_));
 sky130_fd_sc_hd__a211oi_1 _24006_ (.A1(_13897_),
    .A2(_13890_),
    .B1(_13896_),
    .C1(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__o31ai_1 _24007_ (.A1(_09764_),
    .A2(_09771_),
    .A3(_09778_),
    .B1(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__a21oi_1 _24008_ (.A1(_13904_),
    .A2(_09781_),
    .B1(_13903_),
    .Y(_09782_));
 sky130_fd_sc_hd__xnor2_1 _24009_ (.A(_13910_),
    .B(_09782_),
    .Y(\hash.CA1.p5[13] ));
 sky130_fd_sc_hd__nor2_1 _24010_ (.A(_13896_),
    .B(_13903_),
    .Y(_09783_));
 sky130_fd_sc_hd__o21a_1 _24011_ (.A1(_13897_),
    .A2(_13896_),
    .B1(_13904_),
    .X(_09784_));
 sky130_fd_sc_hd__o21ai_0 _24012_ (.A1(_13903_),
    .A2(_09784_),
    .B1(_13910_),
    .Y(_09785_));
 sky130_fd_sc_hd__a31o_2 _24013_ (.A1(_09774_),
    .A2(_09775_),
    .A3(_09783_),
    .B1(_09785_),
    .X(_09786_));
 sky130_fd_sc_hd__nand2b_1 _24014_ (.A_N(_13909_),
    .B(_09786_),
    .Y(_09787_));
 sky130_fd_sc_hd__xor2_1 _24015_ (.A(_13916_),
    .B(_09787_),
    .X(\hash.CA1.p5[14] ));
 sky130_fd_sc_hd__inv_1 _24016_ (.A(_13910_),
    .Y(_09788_));
 sky130_fd_sc_hd__o21bai_2 _24017_ (.A1(_09788_),
    .A2(_09782_),
    .B1_N(_13909_),
    .Y(_09789_));
 sky130_fd_sc_hd__a21oi_1 _24018_ (.A1(_13916_),
    .A2(_09789_),
    .B1(_13915_),
    .Y(_09790_));
 sky130_fd_sc_hd__xnor2_1 _24019_ (.A(_13923_),
    .B(_09790_),
    .Y(\hash.CA1.p5[15] ));
 sky130_fd_sc_hd__nor3_1 _24020_ (.A(_13909_),
    .B(_13915_),
    .C(_13922_),
    .Y(_09791_));
 sky130_fd_sc_hd__or2_0 _24021_ (.A(_13916_),
    .B(_13915_),
    .X(_09792_));
 sky130_fd_sc_hd__a21oi_1 _24022_ (.A1(_13923_),
    .A2(_09792_),
    .B1(_13922_),
    .Y(_09793_));
 sky130_fd_sc_hd__a21oi_1 _24023_ (.A1(_09786_),
    .A2(_09791_),
    .B1(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__xor2_1 _24024_ (.A(_13930_),
    .B(_09794_),
    .X(\hash.CA1.p5[16] ));
 sky130_fd_sc_hd__nand2_1 _24025_ (.A(_13923_),
    .B(_13930_),
    .Y(_09795_));
 sky130_fd_sc_hd__nand2_1 _24026_ (.A(_13916_),
    .B(_13937_),
    .Y(_09796_));
 sky130_fd_sc_hd__nor2_1 _24027_ (.A(_09795_),
    .B(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__inv_1 _24028_ (.A(_13937_),
    .Y(_09798_));
 sky130_fd_sc_hd__a21oi_1 _24029_ (.A1(_13930_),
    .A2(_13922_),
    .B1(_13929_),
    .Y(_09799_));
 sky130_fd_sc_hd__nand2_1 _24030_ (.A(_13937_),
    .B(_13915_),
    .Y(_09800_));
 sky130_fd_sc_hd__o22ai_1 _24031_ (.A1(_09798_),
    .A2(_09799_),
    .B1(_09795_),
    .B2(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__a21o_1 _24032_ (.A1(_09789_),
    .A2(_09797_),
    .B1(_09801_),
    .X(_09802_));
 sky130_fd_sc_hd__o21ai_0 _24033_ (.A1(_09790_),
    .A2(_09795_),
    .B1(_09799_),
    .Y(_09803_));
 sky130_fd_sc_hd__nor2_1 _24034_ (.A(_13937_),
    .B(_09803_),
    .Y(_09804_));
 sky130_fd_sc_hd__nor2_1 _24035_ (.A(_09802_),
    .B(_09804_),
    .Y(\hash.CA1.p5[17] ));
 sky130_fd_sc_hd__nand3_1 _24036_ (.A(_13930_),
    .B(_13937_),
    .C(_13943_),
    .Y(_09805_));
 sky130_fd_sc_hd__a211oi_2 _24037_ (.A1(_09786_),
    .A2(_09791_),
    .B1(_09793_),
    .C1(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_1 _24038_ (.A(_13943_),
    .B(_13936_),
    .Y(_09807_));
 sky130_fd_sc_hd__nand3_1 _24039_ (.A(_13937_),
    .B(_13943_),
    .C(_13929_),
    .Y(_09808_));
 sky130_fd_sc_hd__nand2_1 _24040_ (.A(_09807_),
    .B(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__a21o_1 _24041_ (.A1(_13930_),
    .A2(_09794_),
    .B1(_13929_),
    .X(_09810_));
 sky130_fd_sc_hd__a211oi_1 _24042_ (.A1(_13937_),
    .A2(_09810_),
    .B1(_13936_),
    .C1(_13943_),
    .Y(_09811_));
 sky130_fd_sc_hd__nor3_1 _24043_ (.A(_09806_),
    .B(_09809_),
    .C(_09811_),
    .Y(\hash.CA1.p5[18] ));
 sky130_fd_sc_hd__o21ai_0 _24044_ (.A1(_13936_),
    .A2(_09802_),
    .B1(_13943_),
    .Y(_09812_));
 sky130_fd_sc_hd__nand2b_1 _24045_ (.A_N(_13942_),
    .B(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__xor2_1 _24046_ (.A(_13948_),
    .B(_09813_),
    .X(\hash.CA1.p5[19] ));
 sky130_fd_sc_hd__o31ai_1 _24047_ (.A1(_13942_),
    .A2(_09806_),
    .A3(_09809_),
    .B1(_13948_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2b_1 _24048_ (.A_N(_13947_),
    .B(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__xor2_1 _24049_ (.A(_13953_),
    .B(_09815_),
    .X(\hash.CA1.p5[20] ));
 sky130_fd_sc_hd__nand2_1 _24050_ (.A(_13948_),
    .B(_13953_),
    .Y(_09816_));
 sky130_fd_sc_hd__a21oi_1 _24051_ (.A1(_13943_),
    .A2(_13936_),
    .B1(_13942_),
    .Y(_09817_));
 sky130_fd_sc_hd__nand2_1 _24052_ (.A(_13953_),
    .B(_13947_),
    .Y(_09818_));
 sky130_fd_sc_hd__o21ai_1 _24053_ (.A1(_09816_),
    .A2(_09817_),
    .B1(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__a41oi_4 _24054_ (.A1(_13943_),
    .A2(_13948_),
    .A3(_13953_),
    .A4(_09802_),
    .B1(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__nor2b_1 _24055_ (.A(_13952_),
    .B_N(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__xnor2_1 _24056_ (.A(_13958_),
    .B(_09821_),
    .Y(\hash.CA1.p5[21] ));
 sky130_fd_sc_hd__or3_1 _24057_ (.A(_13942_),
    .B(_13947_),
    .C(_13952_),
    .X(_09822_));
 sky130_fd_sc_hd__nor3_1 _24058_ (.A(_13948_),
    .B(_13947_),
    .C(_13952_),
    .Y(_09823_));
 sky130_fd_sc_hd__nor2_1 _24059_ (.A(_13953_),
    .B(_13952_),
    .Y(_09824_));
 sky130_fd_sc_hd__nor2_1 _24060_ (.A(_09823_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__o31a_1 _24061_ (.A1(_09806_),
    .A2(_09809_),
    .A3(_09822_),
    .B1(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__a21oi_1 _24062_ (.A1(_13958_),
    .A2(_09826_),
    .B1(_13957_),
    .Y(_09827_));
 sky130_fd_sc_hd__xnor2_1 _24063_ (.A(_13963_),
    .B(_09827_),
    .Y(\hash.CA1.p5[22] ));
 sky130_fd_sc_hd__nor3_1 _24064_ (.A(_13952_),
    .B(_13957_),
    .C(_13962_),
    .Y(_09828_));
 sky130_fd_sc_hd__or2_0 _24065_ (.A(_13958_),
    .B(_13957_),
    .X(_09829_));
 sky130_fd_sc_hd__a21oi_1 _24066_ (.A1(_13963_),
    .A2(_09829_),
    .B1(_13962_),
    .Y(_09830_));
 sky130_fd_sc_hd__a21oi_2 _24067_ (.A1(_09820_),
    .A2(_09828_),
    .B1(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__xor2_1 _24068_ (.A(_13969_),
    .B(_09831_),
    .X(\hash.CA1.p5[23] ));
 sky130_fd_sc_hd__and2_0 _24069_ (.A(_13963_),
    .B(_13957_),
    .X(_09832_));
 sky130_fd_sc_hd__a311o_1 _24070_ (.A1(_13958_),
    .A2(_13963_),
    .A3(_09826_),
    .B1(_09832_),
    .C1(_13962_),
    .X(_09833_));
 sky130_fd_sc_hd__a21oi_1 _24071_ (.A1(_13969_),
    .A2(_09833_),
    .B1(_13968_),
    .Y(_09834_));
 sky130_fd_sc_hd__xnor2_1 _24072_ (.A(_13976_),
    .B(_09834_),
    .Y(\hash.CA1.p5[24] ));
 sky130_fd_sc_hd__a21o_1 _24073_ (.A1(_13969_),
    .A2(_09831_),
    .B1(_13968_),
    .X(_09835_));
 sky130_fd_sc_hd__a21oi_1 _24074_ (.A1(_13976_),
    .A2(_09835_),
    .B1(_13975_),
    .Y(_09836_));
 sky130_fd_sc_hd__xnor2_1 _24075_ (.A(_13983_),
    .B(_09836_),
    .Y(\hash.CA1.p5[25] ));
 sky130_fd_sc_hd__a21o_1 _24076_ (.A1(_13976_),
    .A2(_13968_),
    .B1(_13975_),
    .X(_09837_));
 sky130_fd_sc_hd__a21oi_1 _24077_ (.A1(_13983_),
    .A2(_09837_),
    .B1(_13982_),
    .Y(_09838_));
 sky130_fd_sc_hd__inv_1 _24078_ (.A(_09838_),
    .Y(_09839_));
 sky130_fd_sc_hd__a41oi_4 _24079_ (.A1(_13969_),
    .A2(_13976_),
    .A3(_13983_),
    .A4(_09833_),
    .B1(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__xnor2_1 _24080_ (.A(_13990_),
    .B(_09840_),
    .Y(\hash.CA1.p5[26] ));
 sky130_fd_sc_hd__inv_1 _24081_ (.A(_13990_),
    .Y(_09841_));
 sky130_fd_sc_hd__a41oi_4 _24082_ (.A1(_13969_),
    .A2(_13976_),
    .A3(_13983_),
    .A4(_09831_),
    .B1(_09839_),
    .Y(_09842_));
 sky130_fd_sc_hd__o21bai_1 _24083_ (.A1(_09841_),
    .A2(_09842_),
    .B1_N(_13989_),
    .Y(_09843_));
 sky130_fd_sc_hd__xor2_1 _24084_ (.A(_13997_),
    .B(_09843_),
    .X(\hash.CA1.p5[27] ));
 sky130_fd_sc_hd__o21bai_1 _24085_ (.A1(_09841_),
    .A2(_09840_),
    .B1_N(_13989_),
    .Y(_09844_));
 sky130_fd_sc_hd__a21oi_1 _24086_ (.A1(_13997_),
    .A2(_09844_),
    .B1(_13996_),
    .Y(_09845_));
 sky130_fd_sc_hd__xnor2_1 _24087_ (.A(_14004_),
    .B(_09845_),
    .Y(\hash.CA1.p5[28] ));
 sky130_fd_sc_hd__nand3_1 _24088_ (.A(_13990_),
    .B(_13997_),
    .C(_14004_),
    .Y(_09846_));
 sky130_fd_sc_hd__nand2_1 _24089_ (.A(_13997_),
    .B(_13989_),
    .Y(_09847_));
 sky130_fd_sc_hd__nand2b_1 _24090_ (.A_N(_13996_),
    .B(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__a21oi_1 _24091_ (.A1(_14004_),
    .A2(_09848_),
    .B1(_14003_),
    .Y(_09849_));
 sky130_fd_sc_hd__o21ai_0 _24092_ (.A1(_09842_),
    .A2(_09846_),
    .B1(_09849_),
    .Y(_09850_));
 sky130_fd_sc_hd__xor2_1 _24093_ (.A(_14010_),
    .B(_09850_),
    .X(\hash.CA1.p5[29] ));
 sky130_fd_sc_hd__xnor2_1 _24094_ (.A(_13065_),
    .B(_13843_),
    .Y(\hash.CA1.p5[2] ));
 sky130_fd_sc_hd__o21ai_0 _24095_ (.A1(_09840_),
    .A2(_09846_),
    .B1(_09849_),
    .Y(_09851_));
 sky130_fd_sc_hd__a21oi_1 _24096_ (.A1(_14010_),
    .A2(_09851_),
    .B1(_14009_),
    .Y(_09852_));
 sky130_fd_sc_hd__xnor2_1 _24097_ (.A(_14015_),
    .B(_09852_),
    .Y(\hash.CA1.p5[30] ));
 sky130_fd_sc_hd__nand2_1 _24098_ (.A(_13990_),
    .B(_13997_),
    .Y(_09853_));
 sky130_fd_sc_hd__o21ai_0 _24099_ (.A1(_14004_),
    .A2(_14003_),
    .B1(_14010_),
    .Y(_09854_));
 sky130_fd_sc_hd__nand2b_1 _24100_ (.A_N(_14009_),
    .B(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__a21oi_1 _24101_ (.A1(_14015_),
    .A2(_09855_),
    .B1(_14014_),
    .Y(_09856_));
 sky130_fd_sc_hd__a2111oi_0 _24102_ (.A1(_14015_),
    .A2(_14009_),
    .B1(_14014_),
    .C1(_13996_),
    .D1(_14003_),
    .Y(_09857_));
 sky130_fd_sc_hd__a21o_1 _24103_ (.A1(_09847_),
    .A2(_09857_),
    .B1(_09856_),
    .X(_09858_));
 sky130_fd_sc_hd__o31ai_1 _24104_ (.A1(_09842_),
    .A2(_09853_),
    .A3(_09856_),
    .B1(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__nor2b_1 _24105_ (.A(net521),
    .B_N(\hash.CA2.a_dash[31] ),
    .Y(_09860_));
 sky130_fd_sc_hd__xnor2_1 _24106_ (.A(\hash.CA1.p4[31] ),
    .B(_09860_),
    .Y(_09861_));
 sky130_fd_sc_hd__xnor2_1 _24107_ (.A(_09859_),
    .B(_09861_),
    .Y(\hash.CA1.p5[31] ));
 sky130_fd_sc_hd__xnor2_1 _24108_ (.A(_13849_),
    .B(_09769_),
    .Y(\hash.CA1.p5[3] ));
 sky130_fd_sc_hd__o21a_1 _24109_ (.A1(_13848_),
    .A2(_09759_),
    .B1(_13855_),
    .X(_09862_));
 sky130_fd_sc_hd__nor3_1 _24110_ (.A(_13855_),
    .B(_13848_),
    .C(_09759_),
    .Y(_09863_));
 sky130_fd_sc_hd__nor2_1 _24111_ (.A(_09862_),
    .B(_09863_),
    .Y(\hash.CA1.p5[4] ));
 sky130_fd_sc_hd__a21oi_1 _24112_ (.A1(_13855_),
    .A2(_09770_),
    .B1(_13854_),
    .Y(_09864_));
 sky130_fd_sc_hd__xnor2_1 _24113_ (.A(_13861_),
    .B(_09864_),
    .Y(\hash.CA1.p5[5] ));
 sky130_fd_sc_hd__o21a_1 _24114_ (.A1(_13854_),
    .A2(_09862_),
    .B1(_13861_),
    .X(_09865_));
 sky130_fd_sc_hd__nor2_1 _24115_ (.A(_13860_),
    .B(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__xnor2_1 _24116_ (.A(_13867_),
    .B(_09866_),
    .Y(\hash.CA1.p5[6] ));
 sky130_fd_sc_hd__nor2_1 _24117_ (.A(_13866_),
    .B(_09762_),
    .Y(_09867_));
 sky130_fd_sc_hd__nor2_1 _24118_ (.A(_09867_),
    .B(_09771_),
    .Y(_09868_));
 sky130_fd_sc_hd__xor2_1 _24119_ (.A(_13873_),
    .B(_09868_),
    .X(\hash.CA1.p5[7] ));
 sky130_fd_sc_hd__nand2_1 _24120_ (.A(_09760_),
    .B(_09761_),
    .Y(_09869_));
 sky130_fd_sc_hd__a21o_1 _24121_ (.A1(_09869_),
    .A2(_09763_),
    .B1(_13872_),
    .X(_09870_));
 sky130_fd_sc_hd__xor2_1 _24122_ (.A(_13880_),
    .B(_09870_),
    .X(\hash.CA1.p5[8] ));
 sky130_fd_sc_hd__inv_1 _24123_ (.A(_09763_),
    .Y(_09871_));
 sky130_fd_sc_hd__o21bai_1 _24124_ (.A1(_09871_),
    .A2(_09771_),
    .B1_N(_13872_),
    .Y(_09872_));
 sky130_fd_sc_hd__a21oi_1 _24125_ (.A1(_13880_),
    .A2(_09872_),
    .B1(_13879_),
    .Y(_09873_));
 sky130_fd_sc_hd__xnor2_1 _24126_ (.A(_13886_),
    .B(_09873_),
    .Y(\hash.CA1.p5[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_633 ();
 sky130_fd_sc_hd__or2_0 _24138_ (.A(\hash.CA2.S1.X[2] ),
    .B(\hash.reset ),
    .X(\hash.CA1.f[2] ));
 sky130_fd_sc_hd__inv_1 _24139_ (.A(\hash.CA1.f[2] ),
    .Y(_00813_));
 sky130_fd_sc_hd__or2_2 _24140_ (.A(net520),
    .B(\hash.CA2.b_dash[1] ),
    .X(_12828_));
 sky130_fd_sc_hd__inv_1 _24141_ (.A(_12828_),
    .Y(_00751_));
 sky130_fd_sc_hd__or2_1 _24142_ (.A(net520),
    .B(\hash.CA2.a_dash[1] ),
    .X(_13067_));
 sky130_fd_sc_hd__inv_1 _24143_ (.A(_13067_),
    .Y(_00721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_632 ();
 sky130_fd_sc_hd__or2_0 _24145_ (.A(net520),
    .B(_13090_),
    .X(\hash.CA1.b[0] ));
 sky130_fd_sc_hd__inv_1 _24146_ (.A(\hash.CA1.b[0] ),
    .Y(_00690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_630 ();
 sky130_fd_sc_hd__or2_0 _24149_ (.A(\hash.reset ),
    .B(\hash.CA2.S1.X[3] ),
    .X(\hash.CA1.f[3] ));
 sky130_fd_sc_hd__inv_1 _24150_ (.A(\hash.CA1.f[3] ),
    .Y(_14019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_629 ();
 sky130_fd_sc_hd__nand4_4 _24152_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_13709_),
    .D(\count_2[5] ),
    .Y(_09889_));
 sky130_fd_sc_hd__or2_2 _24153_ (.A(\count_2[6] ),
    .B(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_628 ();
 sky130_fd_sc_hd__inv_1 _24155_ (.A(_09890_),
    .Y(_00128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_627 ();
 sky130_fd_sc_hd__clkinv_16 _24157_ (.A(net762),
    .Y(_09893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_623 ();
 sky130_fd_sc_hd__nor3_4 _24162_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .Y(_09897_));
 sky130_fd_sc_hd__nand2_1 _24163_ (.A(_13696_),
    .B(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__nand2_8 _24164_ (.A(_09893_),
    .B(_09898_),
    .Y(_00127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_621 ();
 sky130_fd_sc_hd__nor3b_4 _24167_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C_N(\count_1[3] ),
    .Y(_09901_));
 sky130_fd_sc_hd__nand2_2 _24168_ (.A(_13699_),
    .B(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__nand2_8 _24169_ (.A(_09893_),
    .B(_09902_),
    .Y(_00126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_620 ();
 sky130_fd_sc_hd__nand2_2 _24171_ (.A(_13697_),
    .B(_09901_),
    .Y(_09904_));
 sky130_fd_sc_hd__nand2_8 _24172_ (.A(_09893_),
    .B(_09904_),
    .Y(_00125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_619 ();
 sky130_fd_sc_hd__nand2_2 _24174_ (.A(_13701_),
    .B(_09901_),
    .Y(_09906_));
 sky130_fd_sc_hd__nand2_8 _24175_ (.A(_09893_),
    .B(_09906_),
    .Y(_00124_));
 sky130_fd_sc_hd__nor3b_4 _24176_ (.A(\count_1[5] ),
    .B(\count_1[3] ),
    .C_N(\count_1[4] ),
    .Y(_09907_));
 sky130_fd_sc_hd__nand2_2 _24177_ (.A(_13696_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__nand2_8 _24178_ (.A(_09893_),
    .B(_09908_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_2 _24179_ (.A(_13699_),
    .B(_09907_),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_8 _24180_ (.A(_09893_),
    .B(_09909_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_2 _24181_ (.A(_13697_),
    .B(_09907_),
    .Y(_09910_));
 sky130_fd_sc_hd__nand2_8 _24182_ (.A(_09893_),
    .B(_09910_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_1 _24183_ (.A(_13701_),
    .B(_09907_),
    .Y(_09911_));
 sky130_fd_sc_hd__nand2_8 _24184_ (.A(_09893_),
    .B(_09911_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_2 _24185_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .Y(_09912_));
 sky130_fd_sc_hd__nor2_8 _24186_ (.A(\count_1[5] ),
    .B(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__nand2_1 _24187_ (.A(_13696_),
    .B(_09913_),
    .Y(_09914_));
 sky130_fd_sc_hd__nand2_8 _24188_ (.A(_09893_),
    .B(_09914_),
    .Y(_00119_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_617 ();
 sky130_fd_sc_hd__nand2_2 _24191_ (.A(_13699_),
    .B(_09913_),
    .Y(_09917_));
 sky130_fd_sc_hd__nand2_8 _24192_ (.A(_09893_),
    .B(_09917_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_2 _24193_ (.A(_13697_),
    .B(_09913_),
    .Y(_09918_));
 sky130_fd_sc_hd__nand2_8 _24194_ (.A(_09893_),
    .B(_09918_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_2 _24195_ (.A(_13699_),
    .B(_09897_),
    .Y(_09919_));
 sky130_fd_sc_hd__nand2_8 _24196_ (.A(_09893_),
    .B(_09919_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_2 _24197_ (.A(_13701_),
    .B(_09913_),
    .Y(_09920_));
 sky130_fd_sc_hd__nand2_8 _24198_ (.A(_09893_),
    .B(_09920_),
    .Y(_00115_));
 sky130_fd_sc_hd__nor3b_4 _24199_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C_N(\count_1[5] ),
    .Y(_09921_));
 sky130_fd_sc_hd__nand2_2 _24200_ (.A(_13696_),
    .B(_09921_),
    .Y(_09922_));
 sky130_fd_sc_hd__nand2_8 _24201_ (.A(_09893_),
    .B(_09922_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_2 _24202_ (.A(_13699_),
    .B(_09921_),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_8 _24203_ (.A(_09893_),
    .B(_09923_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_2 _24204_ (.A(_13697_),
    .B(_09921_),
    .Y(_09924_));
 sky130_fd_sc_hd__nand2_8 _24205_ (.A(_09893_),
    .B(_09924_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_2 _24206_ (.A(_13701_),
    .B(_09921_),
    .Y(_09925_));
 sky130_fd_sc_hd__nand2_8 _24207_ (.A(_09893_),
    .B(_09925_),
    .Y(_00111_));
 sky130_fd_sc_hd__and3b_4 _24208_ (.A_N(\count_1[4] ),
    .B(\count_1[3] ),
    .C(\count_1[5] ),
    .X(_09926_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_616 ();
 sky130_fd_sc_hd__nand2_1 _24210_ (.A(_13696_),
    .B(_09926_),
    .Y(_09928_));
 sky130_fd_sc_hd__nand2_8 _24211_ (.A(_09893_),
    .B(_09928_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_2 _24212_ (.A(_13699_),
    .B(_09926_),
    .Y(_09929_));
 sky130_fd_sc_hd__nand2_8 _24213_ (.A(_09893_),
    .B(_09929_),
    .Y(_00109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_615 ();
 sky130_fd_sc_hd__nand2_2 _24215_ (.A(_13697_),
    .B(_09926_),
    .Y(_09931_));
 sky130_fd_sc_hd__nand2_8 _24216_ (.A(_09893_),
    .B(_09931_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_2 _24217_ (.A(_13701_),
    .B(_09926_),
    .Y(_09932_));
 sky130_fd_sc_hd__nand2_8 _24218_ (.A(_09893_),
    .B(_09932_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3b_4 _24219_ (.A_N(\count_1[3] ),
    .B(\count_1[4] ),
    .C(\count_1[5] ),
    .X(_09933_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_614 ();
 sky130_fd_sc_hd__nand2_2 _24221_ (.A(_13696_),
    .B(_09933_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_8 _24222_ (.A(_09893_),
    .B(_09935_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_2 _24223_ (.A(_13697_),
    .B(_09897_),
    .Y(_09936_));
 sky130_fd_sc_hd__nand2_8 _24224_ (.A(_09893_),
    .B(_09936_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_2 _24225_ (.A(_13699_),
    .B(_09933_),
    .Y(_09937_));
 sky130_fd_sc_hd__nand2_8 _24226_ (.A(_09893_),
    .B(_09937_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_2 _24227_ (.A(_13697_),
    .B(_09933_),
    .Y(_09938_));
 sky130_fd_sc_hd__nand2_8 _24228_ (.A(_09893_),
    .B(_09938_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_2 _24229_ (.A(_13701_),
    .B(_09933_),
    .Y(_09939_));
 sky130_fd_sc_hd__nand2_8 _24230_ (.A(_09893_),
    .B(_09939_),
    .Y(_00102_));
 sky130_fd_sc_hd__and3_4 _24231_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .X(_09940_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_613 ();
 sky130_fd_sc_hd__nand2_1 _24233_ (.A(_13696_),
    .B(_09940_),
    .Y(_09942_));
 sky130_fd_sc_hd__nand2_8 _24234_ (.A(_09893_),
    .B(_09942_),
    .Y(_00101_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_610 ();
 sky130_fd_sc_hd__nor3b_4 _24238_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .C_N(\count_2[3] ),
    .Y(_09946_));
 sky130_fd_sc_hd__nand2_2 _24239_ (.A(_13707_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__nand2_8 _24240_ (.A(_09893_),
    .B(_09947_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_2 _24241_ (.A(_13699_),
    .B(_09940_),
    .Y(_09948_));
 sky130_fd_sc_hd__nand2_8 _24242_ (.A(_09893_),
    .B(_09948_),
    .Y(_00100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_608 ();
 sky130_fd_sc_hd__nand2_2 _24245_ (.A(_13705_),
    .B(_09946_),
    .Y(_09951_));
 sky130_fd_sc_hd__nand2_8 _24246_ (.A(_09893_),
    .B(_09951_),
    .Y(_00094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_607 ();
 sky130_fd_sc_hd__nand2_1 _24248_ (.A(_13709_),
    .B(_09946_),
    .Y(_09953_));
 sky130_fd_sc_hd__nand2_8 _24249_ (.A(_09893_),
    .B(_09953_),
    .Y(_00093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_606 ();
 sky130_fd_sc_hd__nand2b_4 _24251_ (.A_N(\count_2[3] ),
    .B(\count_2[4] ),
    .Y(_09955_));
 sky130_fd_sc_hd__nor2_8 _24252_ (.A(\count_2[5] ),
    .B(_09955_),
    .Y(_09956_));
 sky130_fd_sc_hd__nand2_2 _24253_ (.A(_13704_),
    .B(_09956_),
    .Y(_09957_));
 sky130_fd_sc_hd__nand2_8 _24254_ (.A(_09893_),
    .B(_09957_),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_2 _24255_ (.A(_13707_),
    .B(_09956_),
    .Y(_09958_));
 sky130_fd_sc_hd__nand2_8 _24256_ (.A(_09893_),
    .B(_09958_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor3_4 _24257_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(\count_2[5] ),
    .Y(_09959_));
 sky130_fd_sc_hd__nand2_2 _24258_ (.A(_13704_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__nand2_8 _24259_ (.A(_09893_),
    .B(_09960_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_2 _24260_ (.A(_13705_),
    .B(_09956_),
    .Y(_09961_));
 sky130_fd_sc_hd__nand2_8 _24261_ (.A(_09893_),
    .B(_09961_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_2 _24262_ (.A(_13697_),
    .B(_09940_),
    .Y(_09962_));
 sky130_fd_sc_hd__nand2_8 _24263_ (.A(_09893_),
    .B(_09962_),
    .Y(_00099_));
 sky130_fd_sc_hd__clkinv_4 _24264_ (.A(\count_2[5] ),
    .Y(_09963_));
 sky130_fd_sc_hd__nand2_2 _24265_ (.A(_13709_),
    .B(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__o21ai_4 _24266_ (.A1(_09955_),
    .A2(_09964_),
    .B1(_09893_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_4 _24267_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .Y(_09965_));
 sky130_fd_sc_hd__nor2_8 _24268_ (.A(\count_2[5] ),
    .B(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__nand2_2 _24269_ (.A(_13704_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__nand2_8 _24270_ (.A(_09893_),
    .B(_09967_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand2_1 _24271_ (.A(_13707_),
    .B(_09966_),
    .Y(_09968_));
 sky130_fd_sc_hd__nand2_8 _24272_ (.A(_09893_),
    .B(_09968_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_1 _24273_ (.A(_13705_),
    .B(_09966_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand2_8 _24274_ (.A(_09893_),
    .B(_09969_),
    .Y(_00085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_605 ();
 sky130_fd_sc_hd__nand2_2 _24276_ (.A(_13709_),
    .B(_09966_),
    .Y(_09971_));
 sky130_fd_sc_hd__nand2_8 _24277_ (.A(_09893_),
    .B(_09971_),
    .Y(_00084_));
 sky130_fd_sc_hd__nor3_4 _24278_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_09963_),
    .Y(_09972_));
 sky130_fd_sc_hd__nand2_2 _24279_ (.A(_13704_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__nand2_8 _24280_ (.A(_09893_),
    .B(_09973_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_2 _24281_ (.A(_13701_),
    .B(_09940_),
    .Y(_09974_));
 sky130_fd_sc_hd__nand2_8 _24282_ (.A(_09893_),
    .B(_09974_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_2 _24283_ (.A(_13707_),
    .B(_09972_),
    .Y(_09975_));
 sky130_fd_sc_hd__nand2_8 _24284_ (.A(_09893_),
    .B(_09975_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand2_2 _24285_ (.A(_13705_),
    .B(_09972_),
    .Y(_09976_));
 sky130_fd_sc_hd__nand2_8 _24286_ (.A(_09893_),
    .B(_09976_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_2 _24287_ (.A(_13709_),
    .B(\count_2[5] ),
    .Y(_09977_));
 sky130_fd_sc_hd__o31ai_4 _24288_ (.A1(\count_2[4] ),
    .A2(\count_2[3] ),
    .A3(_09977_),
    .B1(_09893_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_2 _24289_ (.A(_13707_),
    .B(_09959_),
    .Y(_09978_));
 sky130_fd_sc_hd__nand2_8 _24290_ (.A(_09893_),
    .B(_09978_),
    .Y(_00079_));
 sky130_fd_sc_hd__nor3b_4 _24291_ (.A(_09963_),
    .B(\count_2[4] ),
    .C_N(\count_2[3] ),
    .Y(_09979_));
 sky130_fd_sc_hd__nand2_2 _24292_ (.A(_13704_),
    .B(_09979_),
    .Y(_09980_));
 sky130_fd_sc_hd__nand2_8 _24293_ (.A(_09893_),
    .B(_09980_),
    .Y(_00078_));
 sky130_fd_sc_hd__nand2_2 _24294_ (.A(_13707_),
    .B(_09979_),
    .Y(_09981_));
 sky130_fd_sc_hd__nand2_8 _24295_ (.A(_09893_),
    .B(_09981_),
    .Y(_00077_));
 sky130_fd_sc_hd__nand2_2 _24296_ (.A(_13701_),
    .B(_09897_),
    .Y(_09982_));
 sky130_fd_sc_hd__nand2_8 _24297_ (.A(_09893_),
    .B(_09982_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_2 _24298_ (.A(_13705_),
    .B(_09979_),
    .Y(_09983_));
 sky130_fd_sc_hd__nand2_8 _24299_ (.A(_09893_),
    .B(_09983_),
    .Y(_00076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_604 ();
 sky130_fd_sc_hd__nand2_2 _24301_ (.A(_13709_),
    .B(_09979_),
    .Y(_09985_));
 sky130_fd_sc_hd__nand2_8 _24302_ (.A(_09893_),
    .B(_09985_),
    .Y(_00075_));
 sky130_fd_sc_hd__nor2_8 _24303_ (.A(_09963_),
    .B(_09955_),
    .Y(_09986_));
 sky130_fd_sc_hd__nand2_2 _24304_ (.A(_13704_),
    .B(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_8 _24305_ (.A(_09893_),
    .B(_09987_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_2 _24306_ (.A(_13707_),
    .B(_09986_),
    .Y(_09988_));
 sky130_fd_sc_hd__nand2_8 _24307_ (.A(_09893_),
    .B(_09988_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_2 _24308_ (.A(_13705_),
    .B(_09986_),
    .Y(_09989_));
 sky130_fd_sc_hd__nand2_8 _24309_ (.A(_09893_),
    .B(_09989_),
    .Y(_00072_));
 sky130_fd_sc_hd__o21ai_4 _24310_ (.A1(_09977_),
    .A2(_09955_),
    .B1(_09893_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand2_2 _24311_ (.A(_13696_),
    .B(_09901_),
    .Y(_09990_));
 sky130_fd_sc_hd__nand2_8 _24312_ (.A(_09893_),
    .B(_09990_),
    .Y(_00096_));
 sky130_fd_sc_hd__nor2_8 _24313_ (.A(_09963_),
    .B(_09965_),
    .Y(_09991_));
 sky130_fd_sc_hd__nand2_2 _24314_ (.A(_13704_),
    .B(_09991_),
    .Y(_09992_));
 sky130_fd_sc_hd__nand2_8 _24315_ (.A(_09893_),
    .B(_09992_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_2 _24316_ (.A(_13707_),
    .B(_09991_),
    .Y(_09993_));
 sky130_fd_sc_hd__nand2_8 _24317_ (.A(_09893_),
    .B(_09993_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_2 _24318_ (.A(_13705_),
    .B(_09959_),
    .Y(_09994_));
 sky130_fd_sc_hd__nand2_8 _24319_ (.A(_09893_),
    .B(_09994_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_2 _24320_ (.A(_13705_),
    .B(_09991_),
    .Y(_09995_));
 sky130_fd_sc_hd__nand2_8 _24321_ (.A(_09893_),
    .B(_09995_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_8 _24322_ (.A(_09893_),
    .B(_09889_),
    .Y(_00066_));
 sky130_fd_sc_hd__o31ai_4 _24323_ (.A1(\count_2[4] ),
    .A2(\count_2[3] ),
    .A3(_09964_),
    .B1(_09893_),
    .Y(_00065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_603 ();
 sky130_fd_sc_hd__nand2_1 _24325_ (.A(_13704_),
    .B(_09946_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_8 _24326_ (.A(_09893_),
    .B(_09997_),
    .Y(_00064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_597 ();
 sky130_fd_sc_hd__mux4_1 _24333_ (.A0(\w[19][0] ),
    .A1(\w[17][0] ),
    .A2(\w[23][0] ),
    .A3(\w[21][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_595 ();
 sky130_fd_sc_hd__mux4_1 _24336_ (.A0(\w[27][0] ),
    .A1(\w[25][0] ),
    .A2(\w[31][0] ),
    .A3(\w[29][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10007_));
 sky130_fd_sc_hd__mux4_1 _24337_ (.A0(\w[3][0] ),
    .A1(\w[1][0] ),
    .A2(\w[7][0] ),
    .A3(\w[5][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_593 ();
 sky130_fd_sc_hd__mux4_1 _24340_ (.A0(\w[11][0] ),
    .A1(\w[9][0] ),
    .A2(\w[15][0] ),
    .A3(\w[13][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_592 ();
 sky130_fd_sc_hd__xor2_4 _24342_ (.A(\count_hash2[3] ),
    .B(_13076_),
    .X(_10013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_591 ();
 sky130_fd_sc_hd__nand3_4 _24344_ (.A(\count_hash2[3] ),
    .B(\count_hash2[2] ),
    .C(\count_hash2[1] ),
    .Y(_10015_));
 sky130_fd_sc_hd__xor2_4 _24345_ (.A(\count_hash2[4] ),
    .B(_10015_),
    .X(_10016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_590 ();
 sky130_fd_sc_hd__mux4_2 _24347_ (.A0(_10004_),
    .A1(_10007_),
    .A2(_10008_),
    .A3(_10011_),
    .S0(net515),
    .S1(net510),
    .X(_10018_));
 sky130_fd_sc_hd__mux4_1 _24348_ (.A0(\w[51][0] ),
    .A1(\w[49][0] ),
    .A2(\w[55][0] ),
    .A3(\w[53][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10019_));
 sky130_fd_sc_hd__mux4_1 _24349_ (.A0(\w[59][0] ),
    .A1(\w[57][0] ),
    .A2(\w[63][0] ),
    .A3(\w[61][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10020_));
 sky130_fd_sc_hd__mux4_1 _24350_ (.A0(\w[35][0] ),
    .A1(\w[33][0] ),
    .A2(\w[39][0] ),
    .A3(\w[37][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10021_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_588 ();
 sky130_fd_sc_hd__mux4_1 _24353_ (.A0(\w[43][0] ),
    .A1(\w[41][0] ),
    .A2(\w[47][0] ),
    .A3(\w[45][0] ),
    .S0(net540),
    .S1(net486),
    .X(_10024_));
 sky130_fd_sc_hd__mux4_1 _24354_ (.A0(_10019_),
    .A1(_10020_),
    .A2(_10021_),
    .A3(_10024_),
    .S0(net515),
    .S1(net510),
    .X(_10025_));
 sky130_fd_sc_hd__nand3_4 _24355_ (.A(\count_hash2[4] ),
    .B(\count_hash2[3] ),
    .C(_13076_),
    .Y(_10026_));
 sky130_fd_sc_hd__xnor2_4 _24356_ (.A(\count_hash2[5] ),
    .B(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_586 ();
 sky130_fd_sc_hd__mux2i_2 _24359_ (.A0(_10018_),
    .A1(_10025_),
    .S(_10027_),
    .Y(_10030_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_584 ();
 sky130_fd_sc_hd__nand4_2 _24362_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(_13088_),
    .D(\count_hash1[5] ),
    .Y(_10033_));
 sky130_fd_sc_hd__nor2_2 _24363_ (.A(_13082_),
    .B(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__or3_4 _24364_ (.A(\count_hash1[6] ),
    .B(net525),
    .C(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_580 ();
 sky130_fd_sc_hd__nand2_2 _24369_ (.A(reset_hash),
    .B(\w[1][0] ),
    .Y(_10040_));
 sky130_fd_sc_hd__o21ai_4 _24370_ (.A1(_10030_),
    .A2(net453),
    .B1(_10040_),
    .Y(_00032_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_576 ();
 sky130_fd_sc_hd__mux4_1 _24375_ (.A0(\w[19][1] ),
    .A1(\w[17][1] ),
    .A2(\w[23][1] ),
    .A3(\w[21][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_574 ();
 sky130_fd_sc_hd__mux4_1 _24378_ (.A0(\w[27][1] ),
    .A1(\w[25][1] ),
    .A2(\w[31][1] ),
    .A3(\w[29][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_572 ();
 sky130_fd_sc_hd__mux4_1 _24381_ (.A0(\w[3][1] ),
    .A1(\w[1][1] ),
    .A2(\w[7][1] ),
    .A3(\w[5][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_570 ();
 sky130_fd_sc_hd__mux4_1 _24384_ (.A0(\w[11][1] ),
    .A1(\w[9][1] ),
    .A2(\w[15][1] ),
    .A3(\w[13][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_567 ();
 sky130_fd_sc_hd__mux4_1 _24388_ (.A0(_10045_),
    .A1(_10048_),
    .A2(_10051_),
    .A3(_10054_),
    .S0(net515),
    .S1(net510),
    .X(_10058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_565 ();
 sky130_fd_sc_hd__mux4_1 _24391_ (.A0(\w[51][1] ),
    .A1(\w[49][1] ),
    .A2(\w[55][1] ),
    .A3(\w[53][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10061_));
 sky130_fd_sc_hd__mux4_1 _24392_ (.A0(\w[59][1] ),
    .A1(\w[57][1] ),
    .A2(\w[63][1] ),
    .A3(\w[61][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10062_));
 sky130_fd_sc_hd__mux4_1 _24393_ (.A0(\w[35][1] ),
    .A1(\w[33][1] ),
    .A2(\w[39][1] ),
    .A3(\w[37][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_563 ();
 sky130_fd_sc_hd__mux4_1 _24396_ (.A0(\w[43][1] ),
    .A1(\w[41][1] ),
    .A2(\w[47][1] ),
    .A3(\w[45][1] ),
    .S0(net540),
    .S1(net486),
    .X(_10066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_561 ();
 sky130_fd_sc_hd__mux4_1 _24399_ (.A0(_10061_),
    .A1(_10062_),
    .A2(_10063_),
    .A3(_10066_),
    .S0(net515),
    .S1(net510),
    .X(_10069_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_560 ();
 sky130_fd_sc_hd__mux2i_2 _24401_ (.A0(_10058_),
    .A1(_10069_),
    .S(net464),
    .Y(_10071_));
 sky130_fd_sc_hd__nand2_1 _24402_ (.A(reset_hash),
    .B(\w[1][1] ),
    .Y(_10072_));
 sky130_fd_sc_hd__o21ai_4 _24403_ (.A1(net453),
    .A2(_10071_),
    .B1(_10072_),
    .Y(_00043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_559 ();
 sky130_fd_sc_hd__mux4_1 _24405_ (.A0(\w[19][2] ),
    .A1(\w[17][2] ),
    .A2(\w[23][2] ),
    .A3(\w[21][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10074_));
 sky130_fd_sc_hd__mux4_1 _24406_ (.A0(\w[27][2] ),
    .A1(\w[25][2] ),
    .A2(\w[31][2] ),
    .A3(\w[29][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10075_));
 sky130_fd_sc_hd__mux4_1 _24407_ (.A0(\w[3][2] ),
    .A1(\w[1][2] ),
    .A2(\w[7][2] ),
    .A3(\w[5][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10076_));
 sky130_fd_sc_hd__mux4_1 _24408_ (.A0(\w[11][2] ),
    .A1(\w[9][2] ),
    .A2(\w[15][2] ),
    .A3(\w[13][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10077_));
 sky130_fd_sc_hd__mux4_1 _24409_ (.A0(_10074_),
    .A1(_10075_),
    .A2(_10076_),
    .A3(_10077_),
    .S0(net514),
    .S1(net509),
    .X(_10078_));
 sky130_fd_sc_hd__mux4_1 _24410_ (.A0(\w[51][2] ),
    .A1(\w[49][2] ),
    .A2(\w[55][2] ),
    .A3(\w[53][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10079_));
 sky130_fd_sc_hd__mux4_1 _24411_ (.A0(\w[59][2] ),
    .A1(\w[57][2] ),
    .A2(\w[63][2] ),
    .A3(\w[61][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10080_));
 sky130_fd_sc_hd__mux4_1 _24412_ (.A0(\w[35][2] ),
    .A1(\w[33][2] ),
    .A2(\w[39][2] ),
    .A3(\w[37][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10081_));
 sky130_fd_sc_hd__mux4_1 _24413_ (.A0(\w[43][2] ),
    .A1(\w[41][2] ),
    .A2(\w[47][2] ),
    .A3(\w[45][2] ),
    .S0(net542),
    .S1(net487),
    .X(_10082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_557 ();
 sky130_fd_sc_hd__mux4_4 _24416_ (.A0(_10079_),
    .A1(_10080_),
    .A2(_10081_),
    .A3(_10082_),
    .S0(net514),
    .S1(net509),
    .X(_10085_));
 sky130_fd_sc_hd__mux2i_2 _24417_ (.A0(_10078_),
    .A1(_10085_),
    .S(net465),
    .Y(_10086_));
 sky130_fd_sc_hd__nand2_1 _24418_ (.A(reset_hash),
    .B(\w[1][2] ),
    .Y(_10087_));
 sky130_fd_sc_hd__o21ai_4 _24419_ (.A1(net454),
    .A2(_10086_),
    .B1(_10087_),
    .Y(_00054_));
 sky130_fd_sc_hd__mux4_1 _24420_ (.A0(\w[19][3] ),
    .A1(\w[17][3] ),
    .A2(\w[23][3] ),
    .A3(\w[21][3] ),
    .S0(net543),
    .S1(net486),
    .X(_10088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_555 ();
 sky130_fd_sc_hd__mux4_1 _24423_ (.A0(\w[27][3] ),
    .A1(\w[25][3] ),
    .A2(\w[31][3] ),
    .A3(\w[29][3] ),
    .S0(net543),
    .S1(net486),
    .X(_10091_));
 sky130_fd_sc_hd__mux4_1 _24424_ (.A0(\w[3][3] ),
    .A1(\w[1][3] ),
    .A2(\w[7][3] ),
    .A3(\w[5][3] ),
    .S0(net543),
    .S1(net486),
    .X(_10092_));
 sky130_fd_sc_hd__mux4_1 _24425_ (.A0(\w[11][3] ),
    .A1(\w[9][3] ),
    .A2(\w[15][3] ),
    .A3(\w[13][3] ),
    .S0(net543),
    .S1(net486),
    .X(_10093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_553 ();
 sky130_fd_sc_hd__mux4_1 _24428_ (.A0(_10088_),
    .A1(_10091_),
    .A2(_10092_),
    .A3(_10093_),
    .S0(net515),
    .S1(net510),
    .X(_10096_));
 sky130_fd_sc_hd__mux4_1 _24429_ (.A0(\w[51][3] ),
    .A1(\w[49][3] ),
    .A2(\w[55][3] ),
    .A3(\w[53][3] ),
    .S0(net540),
    .S1(net486),
    .X(_10097_));
 sky130_fd_sc_hd__mux4_1 _24430_ (.A0(\w[59][3] ),
    .A1(\w[57][3] ),
    .A2(\w[63][3] ),
    .A3(\w[61][3] ),
    .S0(net540),
    .S1(net486),
    .X(_10098_));
 sky130_fd_sc_hd__mux4_1 _24431_ (.A0(\w[35][3] ),
    .A1(\w[33][3] ),
    .A2(\w[39][3] ),
    .A3(\w[37][3] ),
    .S0(net540),
    .S1(net486),
    .X(_10099_));
 sky130_fd_sc_hd__mux4_1 _24432_ (.A0(\w[43][3] ),
    .A1(\w[41][3] ),
    .A2(\w[47][3] ),
    .A3(\w[45][3] ),
    .S0(net540),
    .S1(net486),
    .X(_10100_));
 sky130_fd_sc_hd__mux4_2 _24433_ (.A0(_10097_),
    .A1(_10098_),
    .A2(_10099_),
    .A3(_10100_),
    .S0(net513),
    .S1(net508),
    .X(_10101_));
 sky130_fd_sc_hd__mux2i_2 _24434_ (.A0(_10096_),
    .A1(_10101_),
    .S(net464),
    .Y(_10102_));
 sky130_fd_sc_hd__nand2_1 _24435_ (.A(reset_hash),
    .B(\w[1][3] ),
    .Y(_10103_));
 sky130_fd_sc_hd__o21ai_4 _24436_ (.A1(net453),
    .A2(_10102_),
    .B1(_10103_),
    .Y(_00057_));
 sky130_fd_sc_hd__mux4_1 _24437_ (.A0(\w[19][4] ),
    .A1(\w[17][4] ),
    .A2(\w[23][4] ),
    .A3(\w[21][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10104_));
 sky130_fd_sc_hd__mux4_1 _24438_ (.A0(\w[27][4] ),
    .A1(\w[25][4] ),
    .A2(\w[31][4] ),
    .A3(\w[29][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10105_));
 sky130_fd_sc_hd__mux4_1 _24439_ (.A0(\w[3][4] ),
    .A1(\w[1][4] ),
    .A2(\w[7][4] ),
    .A3(\w[5][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10106_));
 sky130_fd_sc_hd__mux4_1 _24440_ (.A0(\w[11][4] ),
    .A1(\w[9][4] ),
    .A2(\w[15][4] ),
    .A3(\w[13][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10107_));
 sky130_fd_sc_hd__mux4_1 _24441_ (.A0(_10104_),
    .A1(_10105_),
    .A2(_10106_),
    .A3(_10107_),
    .S0(net515),
    .S1(net510),
    .X(_10108_));
 sky130_fd_sc_hd__mux4_1 _24442_ (.A0(\w[51][4] ),
    .A1(\w[49][4] ),
    .A2(\w[55][4] ),
    .A3(\w[53][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10109_));
 sky130_fd_sc_hd__mux4_1 _24443_ (.A0(\w[59][4] ),
    .A1(\w[57][4] ),
    .A2(\w[63][4] ),
    .A3(\w[61][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10110_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_551 ();
 sky130_fd_sc_hd__mux4_1 _24446_ (.A0(\w[35][4] ),
    .A1(\w[33][4] ),
    .A2(\w[39][4] ),
    .A3(\w[37][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10113_));
 sky130_fd_sc_hd__mux4_1 _24447_ (.A0(\w[43][4] ),
    .A1(\w[41][4] ),
    .A2(\w[47][4] ),
    .A3(\w[45][4] ),
    .S0(net540),
    .S1(net486),
    .X(_10114_));
 sky130_fd_sc_hd__mux4_2 _24448_ (.A0(_10109_),
    .A1(_10110_),
    .A2(_10113_),
    .A3(_10114_),
    .S0(net515),
    .S1(net510),
    .X(_10115_));
 sky130_fd_sc_hd__mux2i_2 _24449_ (.A0(_10108_),
    .A1(_10115_),
    .S(_10027_),
    .Y(_10116_));
 sky130_fd_sc_hd__nand2_1 _24450_ (.A(reset_hash),
    .B(\w[1][4] ),
    .Y(_10117_));
 sky130_fd_sc_hd__o21ai_4 _24451_ (.A1(net453),
    .A2(_10116_),
    .B1(_10117_),
    .Y(_00058_));
 sky130_fd_sc_hd__mux4_1 _24452_ (.A0(\w[19][5] ),
    .A1(\w[17][5] ),
    .A2(\w[23][5] ),
    .A3(\w[21][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10118_));
 sky130_fd_sc_hd__mux4_1 _24453_ (.A0(\w[27][5] ),
    .A1(\w[25][5] ),
    .A2(\w[31][5] ),
    .A3(\w[29][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10119_));
 sky130_fd_sc_hd__mux4_1 _24454_ (.A0(\w[3][5] ),
    .A1(\w[1][5] ),
    .A2(\w[7][5] ),
    .A3(\w[5][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10120_));
 sky130_fd_sc_hd__mux4_1 _24455_ (.A0(\w[11][5] ),
    .A1(\w[9][5] ),
    .A2(\w[15][5] ),
    .A3(\w[13][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10121_));
 sky130_fd_sc_hd__mux4_1 _24456_ (.A0(_10118_),
    .A1(_10119_),
    .A2(_10120_),
    .A3(_10121_),
    .S0(net515),
    .S1(net510),
    .X(_10122_));
 sky130_fd_sc_hd__mux4_1 _24457_ (.A0(\w[51][5] ),
    .A1(\w[49][5] ),
    .A2(\w[55][5] ),
    .A3(\w[53][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10123_));
 sky130_fd_sc_hd__mux4_1 _24458_ (.A0(\w[59][5] ),
    .A1(\w[57][5] ),
    .A2(\w[63][5] ),
    .A3(\w[61][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10124_));
 sky130_fd_sc_hd__mux4_1 _24459_ (.A0(\w[35][5] ),
    .A1(\w[33][5] ),
    .A2(\w[39][5] ),
    .A3(\w[37][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10125_));
 sky130_fd_sc_hd__mux4_1 _24460_ (.A0(\w[43][5] ),
    .A1(\w[41][5] ),
    .A2(\w[47][5] ),
    .A3(\w[45][5] ),
    .S0(net543),
    .S1(net486),
    .X(_10126_));
 sky130_fd_sc_hd__mux4_1 _24461_ (.A0(_10123_),
    .A1(_10124_),
    .A2(_10125_),
    .A3(_10126_),
    .S0(net513),
    .S1(net508),
    .X(_10127_));
 sky130_fd_sc_hd__mux2i_2 _24462_ (.A0(_10122_),
    .A1(_10127_),
    .S(net464),
    .Y(_10128_));
 sky130_fd_sc_hd__nand2_1 _24463_ (.A(reset_hash),
    .B(\w[1][5] ),
    .Y(_10129_));
 sky130_fd_sc_hd__o21ai_4 _24464_ (.A1(net453),
    .A2(_10128_),
    .B1(_10129_),
    .Y(_00059_));
 sky130_fd_sc_hd__mux4_1 _24465_ (.A0(\w[19][6] ),
    .A1(\w[17][6] ),
    .A2(\w[23][6] ),
    .A3(\w[21][6] ),
    .S0(net539),
    .S1(net484),
    .X(_10130_));
 sky130_fd_sc_hd__mux4_1 _24466_ (.A0(\w[27][6] ),
    .A1(\w[25][6] ),
    .A2(\w[31][6] ),
    .A3(\w[29][6] ),
    .S0(net539),
    .S1(net484),
    .X(_10131_));
 sky130_fd_sc_hd__mux4_1 _24467_ (.A0(\w[3][6] ),
    .A1(\w[1][6] ),
    .A2(\w[7][6] ),
    .A3(\w[5][6] ),
    .S0(net539),
    .S1(net484),
    .X(_10132_));
 sky130_fd_sc_hd__mux4_1 _24468_ (.A0(\w[11][6] ),
    .A1(\w[9][6] ),
    .A2(\w[15][6] ),
    .A3(\w[13][6] ),
    .S0(net539),
    .S1(net484),
    .X(_10133_));
 sky130_fd_sc_hd__mux4_1 _24469_ (.A0(_10130_),
    .A1(_10131_),
    .A2(_10132_),
    .A3(_10133_),
    .S0(net516),
    .S1(net511),
    .X(_10134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_549 ();
 sky130_fd_sc_hd__mux4_1 _24472_ (.A0(\w[51][6] ),
    .A1(\w[49][6] ),
    .A2(\w[55][6] ),
    .A3(\w[53][6] ),
    .S0(net543),
    .S1(net487),
    .X(_10137_));
 sky130_fd_sc_hd__mux4_1 _24473_ (.A0(\w[59][6] ),
    .A1(\w[57][6] ),
    .A2(\w[63][6] ),
    .A3(\w[61][6] ),
    .S0(net543),
    .S1(net487),
    .X(_10138_));
 sky130_fd_sc_hd__mux4_1 _24474_ (.A0(\w[35][6] ),
    .A1(\w[33][6] ),
    .A2(\w[39][6] ),
    .A3(\w[37][6] ),
    .S0(net543),
    .S1(net487),
    .X(_10139_));
 sky130_fd_sc_hd__mux4_1 _24475_ (.A0(\w[43][6] ),
    .A1(\w[41][6] ),
    .A2(\w[47][6] ),
    .A3(\w[45][6] ),
    .S0(net543),
    .S1(net487),
    .X(_10140_));
 sky130_fd_sc_hd__mux4_4 _24476_ (.A0(_10137_),
    .A1(_10138_),
    .A2(_10139_),
    .A3(_10140_),
    .S0(net514),
    .S1(net509),
    .X(_10141_));
 sky130_fd_sc_hd__mux2i_2 _24477_ (.A0(_10134_),
    .A1(_10141_),
    .S(net465),
    .Y(_10142_));
 sky130_fd_sc_hd__nand2_1 _24478_ (.A(reset_hash),
    .B(\w[1][6] ),
    .Y(_10143_));
 sky130_fd_sc_hd__o21ai_4 _24479_ (.A1(net454),
    .A2(_10142_),
    .B1(_10143_),
    .Y(_00060_));
 sky130_fd_sc_hd__mux4_1 _24480_ (.A0(\w[19][7] ),
    .A1(\w[17][7] ),
    .A2(\w[23][7] ),
    .A3(\w[21][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10144_));
 sky130_fd_sc_hd__mux4_1 _24481_ (.A0(\w[27][7] ),
    .A1(\w[25][7] ),
    .A2(\w[31][7] ),
    .A3(\w[29][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_547 ();
 sky130_fd_sc_hd__mux4_1 _24484_ (.A0(\w[3][7] ),
    .A1(\w[1][7] ),
    .A2(\w[7][7] ),
    .A3(\w[5][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10148_));
 sky130_fd_sc_hd__mux4_1 _24485_ (.A0(\w[11][7] ),
    .A1(\w[9][7] ),
    .A2(\w[15][7] ),
    .A3(\w[13][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10149_));
 sky130_fd_sc_hd__mux4_1 _24486_ (.A0(_10144_),
    .A1(_10145_),
    .A2(_10148_),
    .A3(_10149_),
    .S0(net513),
    .S1(net508),
    .X(_10150_));
 sky130_fd_sc_hd__mux4_1 _24487_ (.A0(\w[51][7] ),
    .A1(\w[49][7] ),
    .A2(\w[55][7] ),
    .A3(\w[53][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10151_));
 sky130_fd_sc_hd__mux4_1 _24488_ (.A0(\w[59][7] ),
    .A1(\w[57][7] ),
    .A2(\w[63][7] ),
    .A3(\w[61][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10152_));
 sky130_fd_sc_hd__mux4_1 _24489_ (.A0(\w[35][7] ),
    .A1(\w[33][7] ),
    .A2(\w[39][7] ),
    .A3(\w[37][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10153_));
 sky130_fd_sc_hd__mux4_1 _24490_ (.A0(\w[43][7] ),
    .A1(\w[41][7] ),
    .A2(\w[47][7] ),
    .A3(\w[45][7] ),
    .S0(net541),
    .S1(net485),
    .X(_10154_));
 sky130_fd_sc_hd__mux4_2 _24491_ (.A0(_10151_),
    .A1(_10152_),
    .A2(_10153_),
    .A3(_10154_),
    .S0(net513),
    .S1(net508),
    .X(_10155_));
 sky130_fd_sc_hd__mux2i_2 _24492_ (.A0(_10150_),
    .A1(_10155_),
    .S(net464),
    .Y(_10156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_546 ();
 sky130_fd_sc_hd__nand2_1 _24494_ (.A(reset_hash),
    .B(\w[1][7] ),
    .Y(_10158_));
 sky130_fd_sc_hd__o21ai_4 _24495_ (.A1(net453),
    .A2(_10156_),
    .B1(_10158_),
    .Y(_00061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_544 ();
 sky130_fd_sc_hd__mux4_1 _24498_ (.A0(\w[19][8] ),
    .A1(\w[17][8] ),
    .A2(\w[23][8] ),
    .A3(\w[21][8] ),
    .S0(net539),
    .S1(net484),
    .X(_10161_));
 sky130_fd_sc_hd__mux4_1 _24499_ (.A0(\w[27][8] ),
    .A1(\w[25][8] ),
    .A2(\w[31][8] ),
    .A3(\w[29][8] ),
    .S0(net539),
    .S1(net484),
    .X(_10162_));
 sky130_fd_sc_hd__mux4_1 _24500_ (.A0(\w[3][8] ),
    .A1(\w[1][8] ),
    .A2(\w[7][8] ),
    .A3(\w[5][8] ),
    .S0(net539),
    .S1(net484),
    .X(_10163_));
 sky130_fd_sc_hd__mux4_1 _24501_ (.A0(\w[11][8] ),
    .A1(\w[9][8] ),
    .A2(\w[15][8] ),
    .A3(\w[13][8] ),
    .S0(net539),
    .S1(net484),
    .X(_10164_));
 sky130_fd_sc_hd__mux4_1 _24502_ (.A0(_10161_),
    .A1(_10162_),
    .A2(_10163_),
    .A3(_10164_),
    .S0(net516),
    .S1(net511),
    .X(_10165_));
 sky130_fd_sc_hd__mux4_1 _24503_ (.A0(\w[51][8] ),
    .A1(\w[49][8] ),
    .A2(\w[55][8] ),
    .A3(\w[53][8] ),
    .S0(net542),
    .S1(net487),
    .X(_10166_));
 sky130_fd_sc_hd__mux4_1 _24504_ (.A0(\w[59][8] ),
    .A1(\w[57][8] ),
    .A2(\w[63][8] ),
    .A3(\w[61][8] ),
    .S0(net543),
    .S1(net487),
    .X(_10167_));
 sky130_fd_sc_hd__mux4_1 _24505_ (.A0(\w[35][8] ),
    .A1(\w[33][8] ),
    .A2(\w[39][8] ),
    .A3(\w[37][8] ),
    .S0(net542),
    .S1(net487),
    .X(_10168_));
 sky130_fd_sc_hd__mux4_1 _24506_ (.A0(\w[43][8] ),
    .A1(\w[41][8] ),
    .A2(\w[47][8] ),
    .A3(\w[45][8] ),
    .S0(net542),
    .S1(net487),
    .X(_10169_));
 sky130_fd_sc_hd__mux4_4 _24507_ (.A0(_10166_),
    .A1(_10167_),
    .A2(_10168_),
    .A3(_10169_),
    .S0(net514),
    .S1(net508),
    .X(_10170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_543 ();
 sky130_fd_sc_hd__mux2i_2 _24509_ (.A0(_10165_),
    .A1(_10170_),
    .S(net465),
    .Y(_10172_));
 sky130_fd_sc_hd__nand2_1 _24510_ (.A(reset_hash),
    .B(\w[1][8] ),
    .Y(_10173_));
 sky130_fd_sc_hd__o21ai_4 _24511_ (.A1(net454),
    .A2(_10172_),
    .B1(_10173_),
    .Y(_00062_));
 sky130_fd_sc_hd__mux4_1 _24512_ (.A0(\w[19][9] ),
    .A1(\w[17][9] ),
    .A2(\w[23][9] ),
    .A3(\w[21][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10174_));
 sky130_fd_sc_hd__mux4_1 _24513_ (.A0(\w[27][9] ),
    .A1(\w[25][9] ),
    .A2(\w[31][9] ),
    .A3(\w[29][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10175_));
 sky130_fd_sc_hd__mux4_1 _24514_ (.A0(\w[3][9] ),
    .A1(\w[1][9] ),
    .A2(\w[7][9] ),
    .A3(\w[5][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10176_));
 sky130_fd_sc_hd__mux4_1 _24515_ (.A0(\w[11][9] ),
    .A1(\w[9][9] ),
    .A2(\w[15][9] ),
    .A3(\w[13][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10177_));
 sky130_fd_sc_hd__mux4_1 _24516_ (.A0(_10174_),
    .A1(_10175_),
    .A2(_10176_),
    .A3(_10177_),
    .S0(net517),
    .S1(net512),
    .X(_10178_));
 sky130_fd_sc_hd__mux4_1 _24517_ (.A0(\w[51][9] ),
    .A1(\w[49][9] ),
    .A2(\w[55][9] ),
    .A3(\w[53][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10179_));
 sky130_fd_sc_hd__mux4_1 _24518_ (.A0(\w[59][9] ),
    .A1(\w[57][9] ),
    .A2(\w[63][9] ),
    .A3(\w[61][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10180_));
 sky130_fd_sc_hd__mux4_1 _24519_ (.A0(\w[35][9] ),
    .A1(\w[33][9] ),
    .A2(\w[39][9] ),
    .A3(\w[37][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_541 ();
 sky130_fd_sc_hd__mux4_1 _24522_ (.A0(\w[43][9] ),
    .A1(\w[41][9] ),
    .A2(\w[47][9] ),
    .A3(\w[45][9] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10184_));
 sky130_fd_sc_hd__mux4_1 _24523_ (.A0(_10179_),
    .A1(_10180_),
    .A2(_10181_),
    .A3(_10184_),
    .S0(_10013_),
    .S1(net510),
    .X(_10185_));
 sky130_fd_sc_hd__mux2i_1 _24524_ (.A0(_10178_),
    .A1(_10185_),
    .S(net466),
    .Y(_10186_));
 sky130_fd_sc_hd__nand2_1 _24525_ (.A(net525),
    .B(\w[1][9] ),
    .Y(_10187_));
 sky130_fd_sc_hd__o21ai_1 _24526_ (.A1(net454),
    .A2(_10186_),
    .B1(_10187_),
    .Y(_00063_));
 sky130_fd_sc_hd__mux4_1 _24527_ (.A0(\w[19][10] ),
    .A1(\w[17][10] ),
    .A2(\w[23][10] ),
    .A3(\w[21][10] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10188_));
 sky130_fd_sc_hd__mux4_1 _24528_ (.A0(\w[27][10] ),
    .A1(\w[25][10] ),
    .A2(\w[31][10] ),
    .A3(\w[29][10] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10189_));
 sky130_fd_sc_hd__mux4_1 _24529_ (.A0(\w[3][10] ),
    .A1(\w[1][10] ),
    .A2(\w[7][10] ),
    .A3(\w[5][10] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_539 ();
 sky130_fd_sc_hd__mux4_1 _24532_ (.A0(\w[11][10] ),
    .A1(\w[9][10] ),
    .A2(\w[15][10] ),
    .A3(\w[13][10] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10193_));
 sky130_fd_sc_hd__mux4_1 _24533_ (.A0(_10188_),
    .A1(_10189_),
    .A2(_10190_),
    .A3(_10193_),
    .S0(net517),
    .S1(net512),
    .X(_10194_));
 sky130_fd_sc_hd__mux4_1 _24534_ (.A0(\w[51][10] ),
    .A1(\w[49][10] ),
    .A2(\w[55][10] ),
    .A3(\w[53][10] ),
    .S0(net539),
    .S1(net484),
    .X(_10195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_537 ();
 sky130_fd_sc_hd__mux4_1 _24537_ (.A0(\w[59][10] ),
    .A1(\w[57][10] ),
    .A2(\w[63][10] ),
    .A3(\w[61][10] ),
    .S0(net539),
    .S1(net484),
    .X(_10198_));
 sky130_fd_sc_hd__mux4_1 _24538_ (.A0(\w[35][10] ),
    .A1(\w[33][10] ),
    .A2(\w[39][10] ),
    .A3(\w[37][10] ),
    .S0(net544),
    .S1(net488),
    .X(_10199_));
 sky130_fd_sc_hd__mux4_1 _24539_ (.A0(\w[43][10] ),
    .A1(\w[41][10] ),
    .A2(\w[47][10] ),
    .A3(\w[45][10] ),
    .S0(net544),
    .S1(net488),
    .X(_10200_));
 sky130_fd_sc_hd__mux4_1 _24540_ (.A0(_10195_),
    .A1(_10198_),
    .A2(_10199_),
    .A3(_10200_),
    .S0(net516),
    .S1(net511),
    .X(_10201_));
 sky130_fd_sc_hd__mux2i_1 _24541_ (.A0(_10194_),
    .A1(_10201_),
    .S(net466),
    .Y(_10202_));
 sky130_fd_sc_hd__nand2_1 _24542_ (.A(net525),
    .B(\w[1][10] ),
    .Y(_10203_));
 sky130_fd_sc_hd__o21ai_1 _24543_ (.A1(net454),
    .A2(_10202_),
    .B1(_10203_),
    .Y(_00033_));
 sky130_fd_sc_hd__mux4_1 _24544_ (.A0(\w[19][11] ),
    .A1(\w[17][11] ),
    .A2(\w[23][11] ),
    .A3(\w[21][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10204_));
 sky130_fd_sc_hd__mux4_1 _24545_ (.A0(\w[27][11] ),
    .A1(\w[25][11] ),
    .A2(\w[31][11] ),
    .A3(\w[29][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10205_));
 sky130_fd_sc_hd__mux4_1 _24546_ (.A0(\w[3][11] ),
    .A1(\w[1][11] ),
    .A2(\w[7][11] ),
    .A3(\w[5][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10206_));
 sky130_fd_sc_hd__mux4_1 _24547_ (.A0(\w[11][11] ),
    .A1(\w[9][11] ),
    .A2(\w[15][11] ),
    .A3(\w[13][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10207_));
 sky130_fd_sc_hd__mux4_1 _24548_ (.A0(_10204_),
    .A1(_10205_),
    .A2(_10206_),
    .A3(_10207_),
    .S0(net517),
    .S1(net511),
    .X(_10208_));
 sky130_fd_sc_hd__mux4_1 _24549_ (.A0(\w[51][11] ),
    .A1(\w[49][11] ),
    .A2(\w[55][11] ),
    .A3(\w[53][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10209_));
 sky130_fd_sc_hd__mux4_1 _24550_ (.A0(\w[59][11] ),
    .A1(\w[57][11] ),
    .A2(\w[63][11] ),
    .A3(\w[61][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10210_));
 sky130_fd_sc_hd__mux4_1 _24551_ (.A0(\w[35][11] ),
    .A1(\w[33][11] ),
    .A2(\w[39][11] ),
    .A3(\w[37][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10211_));
 sky130_fd_sc_hd__mux4_1 _24552_ (.A0(\w[43][11] ),
    .A1(\w[41][11] ),
    .A2(\w[47][11] ),
    .A3(\w[45][11] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10212_));
 sky130_fd_sc_hd__mux4_2 _24553_ (.A0(_10209_),
    .A1(_10210_),
    .A2(_10211_),
    .A3(_10212_),
    .S0(net515),
    .S1(net510),
    .X(_10213_));
 sky130_fd_sc_hd__mux2i_1 _24554_ (.A0(_10208_),
    .A1(_10213_),
    .S(net466),
    .Y(_10214_));
 sky130_fd_sc_hd__nand2_1 _24555_ (.A(net525),
    .B(\w[1][11] ),
    .Y(_10215_));
 sky130_fd_sc_hd__o21ai_1 _24556_ (.A1(_10035_),
    .A2(_10214_),
    .B1(_10215_),
    .Y(_00034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_536 ();
 sky130_fd_sc_hd__mux4_1 _24558_ (.A0(\w[19][12] ),
    .A1(\w[17][12] ),
    .A2(\w[23][12] ),
    .A3(\w[21][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10217_));
 sky130_fd_sc_hd__mux4_1 _24559_ (.A0(\w[27][12] ),
    .A1(\w[25][12] ),
    .A2(\w[31][12] ),
    .A3(\w[29][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10218_));
 sky130_fd_sc_hd__mux4_1 _24560_ (.A0(\w[3][12] ),
    .A1(\w[1][12] ),
    .A2(\w[7][12] ),
    .A3(\w[5][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10219_));
 sky130_fd_sc_hd__mux4_1 _24561_ (.A0(\w[11][12] ),
    .A1(\w[9][12] ),
    .A2(\w[15][12] ),
    .A3(\w[13][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10220_));
 sky130_fd_sc_hd__mux4_1 _24562_ (.A0(_10217_),
    .A1(_10218_),
    .A2(_10219_),
    .A3(_10220_),
    .S0(net515),
    .S1(net510),
    .X(_10221_));
 sky130_fd_sc_hd__mux4_1 _24563_ (.A0(\w[51][12] ),
    .A1(\w[49][12] ),
    .A2(\w[55][12] ),
    .A3(\w[53][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10222_));
 sky130_fd_sc_hd__mux4_1 _24564_ (.A0(\w[59][12] ),
    .A1(\w[57][12] ),
    .A2(\w[63][12] ),
    .A3(\w[61][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10223_));
 sky130_fd_sc_hd__mux4_1 _24565_ (.A0(\w[35][12] ),
    .A1(\w[33][12] ),
    .A2(\w[39][12] ),
    .A3(\w[37][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10224_));
 sky130_fd_sc_hd__mux4_1 _24566_ (.A0(\w[43][12] ),
    .A1(\w[41][12] ),
    .A2(\w[47][12] ),
    .A3(\w[45][12] ),
    .S0(net543),
    .S1(net486),
    .X(_10225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_534 ();
 sky130_fd_sc_hd__mux4_4 _24569_ (.A0(_10222_),
    .A1(_10223_),
    .A2(_10224_),
    .A3(_10225_),
    .S0(net513),
    .S1(net508),
    .X(_10228_));
 sky130_fd_sc_hd__mux2i_2 _24570_ (.A0(_10221_),
    .A1(_10228_),
    .S(net464),
    .Y(_10229_));
 sky130_fd_sc_hd__nand2_1 _24571_ (.A(reset_hash),
    .B(\w[1][12] ),
    .Y(_10230_));
 sky130_fd_sc_hd__o21ai_4 _24572_ (.A1(net453),
    .A2(_10229_),
    .B1(_10230_),
    .Y(_00035_));
 sky130_fd_sc_hd__mux4_1 _24573_ (.A0(\w[19][13] ),
    .A1(\w[17][13] ),
    .A2(\w[23][13] ),
    .A3(\w[21][13] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10231_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_532 ();
 sky130_fd_sc_hd__mux4_1 _24576_ (.A0(\w[27][13] ),
    .A1(\w[25][13] ),
    .A2(\w[31][13] ),
    .A3(\w[29][13] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10234_));
 sky130_fd_sc_hd__mux4_1 _24577_ (.A0(\w[3][13] ),
    .A1(\w[1][13] ),
    .A2(\w[7][13] ),
    .A3(\w[5][13] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10235_));
 sky130_fd_sc_hd__mux4_1 _24578_ (.A0(\w[11][13] ),
    .A1(\w[9][13] ),
    .A2(\w[15][13] ),
    .A3(\w[13][13] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10236_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_530 ();
 sky130_fd_sc_hd__mux4_1 _24581_ (.A0(_10231_),
    .A1(_10234_),
    .A2(_10235_),
    .A3(_10236_),
    .S0(net517),
    .S1(net512),
    .X(_10239_));
 sky130_fd_sc_hd__mux4_1 _24582_ (.A0(\w[51][13] ),
    .A1(\w[49][13] ),
    .A2(\w[55][13] ),
    .A3(\w[53][13] ),
    .S0(net544),
    .S1(net488),
    .X(_10240_));
 sky130_fd_sc_hd__mux4_1 _24583_ (.A0(\w[59][13] ),
    .A1(\w[57][13] ),
    .A2(\w[63][13] ),
    .A3(\w[61][13] ),
    .S0(net544),
    .S1(net488),
    .X(_10241_));
 sky130_fd_sc_hd__mux4_1 _24584_ (.A0(\w[35][13] ),
    .A1(\w[33][13] ),
    .A2(\w[39][13] ),
    .A3(\w[37][13] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10242_));
 sky130_fd_sc_hd__mux4_1 _24585_ (.A0(\w[43][13] ),
    .A1(\w[41][13] ),
    .A2(\w[47][13] ),
    .A3(\w[45][13] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10243_));
 sky130_fd_sc_hd__mux4_2 _24586_ (.A0(_10240_),
    .A1(_10241_),
    .A2(_10242_),
    .A3(_10243_),
    .S0(_10013_),
    .S1(net509),
    .X(_10244_));
 sky130_fd_sc_hd__mux2i_1 _24587_ (.A0(_10239_),
    .A1(_10244_),
    .S(net466),
    .Y(_10245_));
 sky130_fd_sc_hd__nand2_1 _24588_ (.A(net525),
    .B(\w[1][13] ),
    .Y(_10246_));
 sky130_fd_sc_hd__o21ai_0 _24589_ (.A1(net454),
    .A2(_10245_),
    .B1(_10246_),
    .Y(_00036_));
 sky130_fd_sc_hd__mux4_1 _24590_ (.A0(\w[19][14] ),
    .A1(\w[17][14] ),
    .A2(\w[23][14] ),
    .A3(\w[21][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10247_));
 sky130_fd_sc_hd__mux4_1 _24591_ (.A0(\w[27][14] ),
    .A1(\w[25][14] ),
    .A2(\w[31][14] ),
    .A3(\w[29][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10248_));
 sky130_fd_sc_hd__mux4_1 _24592_ (.A0(\w[3][14] ),
    .A1(\w[1][14] ),
    .A2(\w[7][14] ),
    .A3(\w[5][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10249_));
 sky130_fd_sc_hd__mux4_1 _24593_ (.A0(\w[11][14] ),
    .A1(\w[9][14] ),
    .A2(\w[15][14] ),
    .A3(\w[13][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10250_));
 sky130_fd_sc_hd__mux4_1 _24594_ (.A0(_10247_),
    .A1(_10248_),
    .A2(_10249_),
    .A3(_10250_),
    .S0(net513),
    .S1(net508),
    .X(_10251_));
 sky130_fd_sc_hd__mux4_1 _24595_ (.A0(\w[51][14] ),
    .A1(\w[49][14] ),
    .A2(\w[55][14] ),
    .A3(\w[53][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10252_));
 sky130_fd_sc_hd__mux4_1 _24596_ (.A0(\w[59][14] ),
    .A1(\w[57][14] ),
    .A2(\w[63][14] ),
    .A3(\w[61][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10253_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_528 ();
 sky130_fd_sc_hd__mux4_1 _24599_ (.A0(\w[35][14] ),
    .A1(\w[33][14] ),
    .A2(\w[39][14] ),
    .A3(\w[37][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10256_));
 sky130_fd_sc_hd__mux4_1 _24600_ (.A0(\w[43][14] ),
    .A1(\w[41][14] ),
    .A2(\w[47][14] ),
    .A3(\w[45][14] ),
    .S0(net541),
    .S1(net485),
    .X(_10257_));
 sky130_fd_sc_hd__mux4_1 _24601_ (.A0(_10252_),
    .A1(_10253_),
    .A2(_10256_),
    .A3(_10257_),
    .S0(net513),
    .S1(net508),
    .X(_10258_));
 sky130_fd_sc_hd__mux2i_2 _24602_ (.A0(_10251_),
    .A1(_10258_),
    .S(net464),
    .Y(_10259_));
 sky130_fd_sc_hd__nand2_1 _24603_ (.A(reset_hash),
    .B(\w[1][14] ),
    .Y(_10260_));
 sky130_fd_sc_hd__o21ai_4 _24604_ (.A1(net453),
    .A2(_10259_),
    .B1(_10260_),
    .Y(_00037_));
 sky130_fd_sc_hd__mux4_1 _24605_ (.A0(\w[19][15] ),
    .A1(\w[17][15] ),
    .A2(\w[23][15] ),
    .A3(\w[21][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10261_));
 sky130_fd_sc_hd__mux4_1 _24606_ (.A0(\w[27][15] ),
    .A1(\w[25][15] ),
    .A2(\w[31][15] ),
    .A3(\w[29][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10262_));
 sky130_fd_sc_hd__mux4_1 _24607_ (.A0(\w[3][15] ),
    .A1(\w[1][15] ),
    .A2(\w[7][15] ),
    .A3(\w[5][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10263_));
 sky130_fd_sc_hd__mux4_1 _24608_ (.A0(\w[11][15] ),
    .A1(\w[9][15] ),
    .A2(\w[15][15] ),
    .A3(\w[13][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10264_));
 sky130_fd_sc_hd__mux4_1 _24609_ (.A0(_10261_),
    .A1(_10262_),
    .A2(_10263_),
    .A3(_10264_),
    .S0(net513),
    .S1(net508),
    .X(_10265_));
 sky130_fd_sc_hd__mux4_1 _24610_ (.A0(\w[51][15] ),
    .A1(\w[49][15] ),
    .A2(\w[55][15] ),
    .A3(\w[53][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10266_));
 sky130_fd_sc_hd__mux4_1 _24611_ (.A0(\w[59][15] ),
    .A1(\w[57][15] ),
    .A2(\w[63][15] ),
    .A3(\w[61][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10267_));
 sky130_fd_sc_hd__mux4_1 _24612_ (.A0(\w[35][15] ),
    .A1(\w[33][15] ),
    .A2(\w[39][15] ),
    .A3(\w[37][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10268_));
 sky130_fd_sc_hd__mux4_1 _24613_ (.A0(\w[43][15] ),
    .A1(\w[41][15] ),
    .A2(\w[47][15] ),
    .A3(\w[45][15] ),
    .S0(net541),
    .S1(net485),
    .X(_10269_));
 sky130_fd_sc_hd__mux4_1 _24614_ (.A0(_10266_),
    .A1(_10267_),
    .A2(_10268_),
    .A3(_10269_),
    .S0(net513),
    .S1(net508),
    .X(_10270_));
 sky130_fd_sc_hd__mux2i_2 _24615_ (.A0(_10265_),
    .A1(_10270_),
    .S(net464),
    .Y(_10271_));
 sky130_fd_sc_hd__nand2_1 _24616_ (.A(reset_hash),
    .B(\w[1][15] ),
    .Y(_10272_));
 sky130_fd_sc_hd__o21ai_4 _24617_ (.A1(net453),
    .A2(_10271_),
    .B1(_10272_),
    .Y(_00038_));
 sky130_fd_sc_hd__mux4_1 _24618_ (.A0(\w[19][16] ),
    .A1(\w[17][16] ),
    .A2(\w[23][16] ),
    .A3(\w[21][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10273_));
 sky130_fd_sc_hd__mux4_1 _24619_ (.A0(\w[27][16] ),
    .A1(\w[25][16] ),
    .A2(\w[31][16] ),
    .A3(\w[29][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10274_));
 sky130_fd_sc_hd__mux4_1 _24620_ (.A0(\w[3][16] ),
    .A1(\w[1][16] ),
    .A2(\w[7][16] ),
    .A3(\w[5][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10275_));
 sky130_fd_sc_hd__mux4_1 _24621_ (.A0(\w[11][16] ),
    .A1(\w[9][16] ),
    .A2(\w[15][16] ),
    .A3(\w[13][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10276_));
 sky130_fd_sc_hd__mux4_1 _24622_ (.A0(_10273_),
    .A1(_10274_),
    .A2(_10275_),
    .A3(_10276_),
    .S0(net513),
    .S1(net508),
    .X(_10277_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_526 ();
 sky130_fd_sc_hd__mux4_1 _24625_ (.A0(\w[51][16] ),
    .A1(\w[49][16] ),
    .A2(\w[55][16] ),
    .A3(\w[53][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10280_));
 sky130_fd_sc_hd__mux4_1 _24626_ (.A0(\w[59][16] ),
    .A1(\w[57][16] ),
    .A2(\w[63][16] ),
    .A3(\w[61][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10281_));
 sky130_fd_sc_hd__mux4_1 _24627_ (.A0(\w[35][16] ),
    .A1(\w[33][16] ),
    .A2(\w[39][16] ),
    .A3(\w[37][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10282_));
 sky130_fd_sc_hd__mux4_1 _24628_ (.A0(\w[43][16] ),
    .A1(\w[41][16] ),
    .A2(\w[47][16] ),
    .A3(\w[45][16] ),
    .S0(net541),
    .S1(net485),
    .X(_10283_));
 sky130_fd_sc_hd__mux4_1 _24629_ (.A0(_10280_),
    .A1(_10281_),
    .A2(_10282_),
    .A3(_10283_),
    .S0(net513),
    .S1(net508),
    .X(_10284_));
 sky130_fd_sc_hd__mux2i_2 _24630_ (.A0(_10277_),
    .A1(_10284_),
    .S(net464),
    .Y(_10285_));
 sky130_fd_sc_hd__nand2_1 _24631_ (.A(reset_hash),
    .B(\w[1][16] ),
    .Y(_10286_));
 sky130_fd_sc_hd__o21ai_4 _24632_ (.A1(net453),
    .A2(_10285_),
    .B1(_10286_),
    .Y(_00039_));
 sky130_fd_sc_hd__mux4_1 _24633_ (.A0(\w[19][17] ),
    .A1(\w[17][17] ),
    .A2(\w[23][17] ),
    .A3(\w[21][17] ),
    .S0(net541),
    .S1(net485),
    .X(_10287_));
 sky130_fd_sc_hd__mux4_1 _24634_ (.A0(\w[27][17] ),
    .A1(\w[25][17] ),
    .A2(\w[31][17] ),
    .A3(\w[29][17] ),
    .S0(net541),
    .S1(net485),
    .X(_10288_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_524 ();
 sky130_fd_sc_hd__mux4_1 _24637_ (.A0(\w[3][17] ),
    .A1(\w[1][17] ),
    .A2(\w[7][17] ),
    .A3(\w[5][17] ),
    .S0(net541),
    .S1(net485),
    .X(_10291_));
 sky130_fd_sc_hd__mux4_1 _24638_ (.A0(\w[11][17] ),
    .A1(\w[9][17] ),
    .A2(\w[15][17] ),
    .A3(\w[13][17] ),
    .S0(net541),
    .S1(net485),
    .X(_10292_));
 sky130_fd_sc_hd__mux4_2 _24639_ (.A0(_10287_),
    .A1(_10288_),
    .A2(_10291_),
    .A3(_10292_),
    .S0(net513),
    .S1(net508),
    .X(_10293_));
 sky130_fd_sc_hd__mux4_1 _24640_ (.A0(\w[51][17] ),
    .A1(\w[49][17] ),
    .A2(\w[55][17] ),
    .A3(\w[53][17] ),
    .S0(net542),
    .S1(net487),
    .X(_10294_));
 sky130_fd_sc_hd__mux4_1 _24641_ (.A0(\w[59][17] ),
    .A1(\w[57][17] ),
    .A2(\w[63][17] ),
    .A3(\w[61][17] ),
    .S0(net542),
    .S1(net487),
    .X(_10295_));
 sky130_fd_sc_hd__mux4_1 _24642_ (.A0(\w[35][17] ),
    .A1(\w[33][17] ),
    .A2(\w[39][17] ),
    .A3(\w[37][17] ),
    .S0(net542),
    .S1(net487),
    .X(_10296_));
 sky130_fd_sc_hd__mux4_1 _24643_ (.A0(\w[43][17] ),
    .A1(\w[41][17] ),
    .A2(\w[47][17] ),
    .A3(\w[45][17] ),
    .S0(net542),
    .S1(net487),
    .X(_10297_));
 sky130_fd_sc_hd__mux4_1 _24644_ (.A0(_10294_),
    .A1(_10295_),
    .A2(_10296_),
    .A3(_10297_),
    .S0(net513),
    .S1(net508),
    .X(_10298_));
 sky130_fd_sc_hd__mux2i_2 _24645_ (.A0(_10293_),
    .A1(_10298_),
    .S(net464),
    .Y(_10299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_523 ();
 sky130_fd_sc_hd__nand2_1 _24647_ (.A(reset_hash),
    .B(\w[1][17] ),
    .Y(_10301_));
 sky130_fd_sc_hd__o21ai_4 _24648_ (.A1(net454),
    .A2(_10299_),
    .B1(_10301_),
    .Y(_00040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_521 ();
 sky130_fd_sc_hd__mux4_1 _24651_ (.A0(\w[19][18] ),
    .A1(\w[17][18] ),
    .A2(\w[23][18] ),
    .A3(\w[21][18] ),
    .S0(net544),
    .S1(net488),
    .X(_10304_));
 sky130_fd_sc_hd__mux4_1 _24652_ (.A0(\w[27][18] ),
    .A1(\w[25][18] ),
    .A2(\w[31][18] ),
    .A3(\w[29][18] ),
    .S0(net544),
    .S1(net488),
    .X(_10305_));
 sky130_fd_sc_hd__mux4_1 _24653_ (.A0(\w[3][18] ),
    .A1(\w[1][18] ),
    .A2(\w[7][18] ),
    .A3(\w[5][18] ),
    .S0(net544),
    .S1(net488),
    .X(_10306_));
 sky130_fd_sc_hd__mux4_1 _24654_ (.A0(\w[11][18] ),
    .A1(\w[9][18] ),
    .A2(\w[15][18] ),
    .A3(\w[13][18] ),
    .S0(net544),
    .S1(net488),
    .X(_10307_));
 sky130_fd_sc_hd__mux4_1 _24655_ (.A0(_10304_),
    .A1(_10305_),
    .A2(_10306_),
    .A3(_10307_),
    .S0(net517),
    .S1(net512),
    .X(_10308_));
 sky130_fd_sc_hd__mux4_1 _24656_ (.A0(\w[51][18] ),
    .A1(\w[49][18] ),
    .A2(\w[55][18] ),
    .A3(\w[53][18] ),
    .S0(net539),
    .S1(net484),
    .X(_10309_));
 sky130_fd_sc_hd__mux4_1 _24657_ (.A0(\w[59][18] ),
    .A1(\w[57][18] ),
    .A2(\w[63][18] ),
    .A3(\w[61][18] ),
    .S0(net539),
    .S1(net484),
    .X(_10310_));
 sky130_fd_sc_hd__mux4_1 _24658_ (.A0(\w[35][18] ),
    .A1(\w[33][18] ),
    .A2(\w[39][18] ),
    .A3(\w[37][18] ),
    .S0(net539),
    .S1(net484),
    .X(_10311_));
 sky130_fd_sc_hd__mux4_1 _24659_ (.A0(\w[43][18] ),
    .A1(\w[41][18] ),
    .A2(\w[47][18] ),
    .A3(\w[45][18] ),
    .S0(net539),
    .S1(net484),
    .X(_10312_));
 sky130_fd_sc_hd__mux4_4 _24660_ (.A0(_10309_),
    .A1(_10310_),
    .A2(_10311_),
    .A3(_10312_),
    .S0(net516),
    .S1(net511),
    .X(_10313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_520 ();
 sky130_fd_sc_hd__mux2i_2 _24662_ (.A0(_10308_),
    .A1(_10313_),
    .S(net465),
    .Y(_10315_));
 sky130_fd_sc_hd__nand2_1 _24663_ (.A(reset_hash),
    .B(\w[1][18] ),
    .Y(_10316_));
 sky130_fd_sc_hd__o21ai_4 _24664_ (.A1(net454),
    .A2(_10315_),
    .B1(_10316_),
    .Y(_00041_));
 sky130_fd_sc_hd__mux4_1 _24665_ (.A0(\w[19][19] ),
    .A1(\w[17][19] ),
    .A2(\w[23][19] ),
    .A3(\w[21][19] ),
    .S0(net544),
    .S1(net488),
    .X(_10317_));
 sky130_fd_sc_hd__mux4_1 _24666_ (.A0(\w[27][19] ),
    .A1(\w[25][19] ),
    .A2(\w[31][19] ),
    .A3(\w[29][19] ),
    .S0(net544),
    .S1(net488),
    .X(_10318_));
 sky130_fd_sc_hd__mux4_1 _24667_ (.A0(\w[3][19] ),
    .A1(\w[1][19] ),
    .A2(\w[7][19] ),
    .A3(\w[5][19] ),
    .S0(net544),
    .S1(net488),
    .X(_10319_));
 sky130_fd_sc_hd__mux4_1 _24668_ (.A0(\w[11][19] ),
    .A1(\w[9][19] ),
    .A2(\w[15][19] ),
    .A3(\w[13][19] ),
    .S0(net544),
    .S1(net488),
    .X(_10320_));
 sky130_fd_sc_hd__mux4_1 _24669_ (.A0(_10317_),
    .A1(_10318_),
    .A2(_10319_),
    .A3(_10320_),
    .S0(net517),
    .S1(net512),
    .X(_10321_));
 sky130_fd_sc_hd__mux4_1 _24670_ (.A0(\w[51][19] ),
    .A1(\w[49][19] ),
    .A2(\w[55][19] ),
    .A3(\w[53][19] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10322_));
 sky130_fd_sc_hd__mux4_1 _24671_ (.A0(\w[59][19] ),
    .A1(\w[57][19] ),
    .A2(\w[63][19] ),
    .A3(\w[61][19] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10323_));
 sky130_fd_sc_hd__mux4_1 _24672_ (.A0(\w[35][19] ),
    .A1(\w[33][19] ),
    .A2(\w[39][19] ),
    .A3(\w[37][19] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10324_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_518 ();
 sky130_fd_sc_hd__mux4_1 _24675_ (.A0(\w[43][19] ),
    .A1(\w[41][19] ),
    .A2(\w[47][19] ),
    .A3(\w[45][19] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10327_));
 sky130_fd_sc_hd__mux4_4 _24676_ (.A0(_10322_),
    .A1(_10323_),
    .A2(_10324_),
    .A3(_10327_),
    .S0(net515),
    .S1(net510),
    .X(_10328_));
 sky130_fd_sc_hd__mux2i_1 _24677_ (.A0(_10321_),
    .A1(_10328_),
    .S(net465),
    .Y(_10329_));
 sky130_fd_sc_hd__nand2_1 _24678_ (.A(reset_hash),
    .B(\w[1][19] ),
    .Y(_10330_));
 sky130_fd_sc_hd__o21ai_2 _24679_ (.A1(net454),
    .A2(_10329_),
    .B1(_10330_),
    .Y(_00042_));
 sky130_fd_sc_hd__mux4_1 _24680_ (.A0(\w[19][20] ),
    .A1(\w[17][20] ),
    .A2(\w[23][20] ),
    .A3(\w[21][20] ),
    .S0(\count_hash2[1] ),
    .S1(_00657_),
    .X(_10331_));
 sky130_fd_sc_hd__mux4_1 _24681_ (.A0(\w[27][20] ),
    .A1(\w[25][20] ),
    .A2(\w[31][20] ),
    .A3(\w[29][20] ),
    .S0(\count_hash2[1] ),
    .S1(_00657_),
    .X(_10332_));
 sky130_fd_sc_hd__mux4_1 _24682_ (.A0(\w[3][20] ),
    .A1(\w[1][20] ),
    .A2(\w[7][20] ),
    .A3(\w[5][20] ),
    .S0(\count_hash2[1] ),
    .S1(_00657_),
    .X(_10333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_516 ();
 sky130_fd_sc_hd__mux4_1 _24685_ (.A0(\w[11][20] ),
    .A1(\w[9][20] ),
    .A2(\w[15][20] ),
    .A3(\w[13][20] ),
    .S0(\count_hash2[1] ),
    .S1(_00657_),
    .X(_10336_));
 sky130_fd_sc_hd__mux4_1 _24686_ (.A0(_10331_),
    .A1(_10332_),
    .A2(_10333_),
    .A3(_10336_),
    .S0(_10013_),
    .S1(_10016_),
    .X(_10337_));
 sky130_fd_sc_hd__mux4_1 _24687_ (.A0(\w[51][20] ),
    .A1(\w[49][20] ),
    .A2(\w[55][20] ),
    .A3(\w[53][20] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_514 ();
 sky130_fd_sc_hd__mux4_1 _24690_ (.A0(\w[59][20] ),
    .A1(\w[57][20] ),
    .A2(\w[63][20] ),
    .A3(\w[61][20] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10341_));
 sky130_fd_sc_hd__mux4_1 _24691_ (.A0(\w[35][20] ),
    .A1(\w[33][20] ),
    .A2(\w[39][20] ),
    .A3(\w[37][20] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10342_));
 sky130_fd_sc_hd__mux4_1 _24692_ (.A0(\w[43][20] ),
    .A1(\w[41][20] ),
    .A2(\w[47][20] ),
    .A3(\w[45][20] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10343_));
 sky130_fd_sc_hd__mux4_2 _24693_ (.A0(_10338_),
    .A1(_10341_),
    .A2(_10342_),
    .A3(_10343_),
    .S0(net515),
    .S1(net510),
    .X(_10344_));
 sky130_fd_sc_hd__mux2i_2 _24694_ (.A0(_10337_),
    .A1(_10344_),
    .S(_10027_),
    .Y(_10345_));
 sky130_fd_sc_hd__nand2_1 _24695_ (.A(net525),
    .B(\w[1][20] ),
    .Y(_10346_));
 sky130_fd_sc_hd__o21ai_4 _24696_ (.A1(_10035_),
    .A2(_10345_),
    .B1(_10346_),
    .Y(_00044_));
 sky130_fd_sc_hd__mux4_1 _24697_ (.A0(\w[19][21] ),
    .A1(\w[17][21] ),
    .A2(\w[23][21] ),
    .A3(\w[21][21] ),
    .S0(net544),
    .S1(net488),
    .X(_10347_));
 sky130_fd_sc_hd__mux4_1 _24698_ (.A0(\w[27][21] ),
    .A1(\w[25][21] ),
    .A2(\w[31][21] ),
    .A3(\w[29][21] ),
    .S0(net544),
    .S1(net488),
    .X(_10348_));
 sky130_fd_sc_hd__mux4_1 _24699_ (.A0(\w[3][21] ),
    .A1(\w[1][21] ),
    .A2(\w[7][21] ),
    .A3(\w[5][21] ),
    .S0(net544),
    .S1(net488),
    .X(_10349_));
 sky130_fd_sc_hd__mux4_1 _24700_ (.A0(\w[11][21] ),
    .A1(\w[9][21] ),
    .A2(\w[15][21] ),
    .A3(\w[13][21] ),
    .S0(net544),
    .S1(net488),
    .X(_10350_));
 sky130_fd_sc_hd__mux4_1 _24701_ (.A0(_10347_),
    .A1(_10348_),
    .A2(_10349_),
    .A3(_10350_),
    .S0(net517),
    .S1(net512),
    .X(_10351_));
 sky130_fd_sc_hd__mux4_1 _24702_ (.A0(\w[51][21] ),
    .A1(\w[49][21] ),
    .A2(\w[55][21] ),
    .A3(\w[53][21] ),
    .S0(net543),
    .S1(net487),
    .X(_10352_));
 sky130_fd_sc_hd__mux4_1 _24703_ (.A0(\w[59][21] ),
    .A1(\w[57][21] ),
    .A2(\w[63][21] ),
    .A3(\w[61][21] ),
    .S0(net543),
    .S1(net487),
    .X(_10353_));
 sky130_fd_sc_hd__mux4_1 _24704_ (.A0(\w[35][21] ),
    .A1(\w[33][21] ),
    .A2(\w[39][21] ),
    .A3(\w[37][21] ),
    .S0(net543),
    .S1(net487),
    .X(_10354_));
 sky130_fd_sc_hd__mux4_1 _24705_ (.A0(\w[43][21] ),
    .A1(\w[41][21] ),
    .A2(\w[47][21] ),
    .A3(\w[45][21] ),
    .S0(net543),
    .S1(net487),
    .X(_10355_));
 sky130_fd_sc_hd__mux4_4 _24706_ (.A0(_10352_),
    .A1(_10353_),
    .A2(_10354_),
    .A3(_10355_),
    .S0(net514),
    .S1(net509),
    .X(_10356_));
 sky130_fd_sc_hd__mux2i_1 _24707_ (.A0(_10351_),
    .A1(_10356_),
    .S(net466),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_1 _24708_ (.A(reset_hash),
    .B(\w[1][21] ),
    .Y(_10358_));
 sky130_fd_sc_hd__o21ai_1 _24709_ (.A1(net454),
    .A2(_10357_),
    .B1(_10358_),
    .Y(_00045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_513 ();
 sky130_fd_sc_hd__mux4_1 _24711_ (.A0(\w[19][22] ),
    .A1(\w[17][22] ),
    .A2(\w[23][22] ),
    .A3(\w[21][22] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10360_));
 sky130_fd_sc_hd__mux4_1 _24712_ (.A0(\w[27][22] ),
    .A1(\w[25][22] ),
    .A2(\w[31][22] ),
    .A3(\w[29][22] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10361_));
 sky130_fd_sc_hd__mux4_1 _24713_ (.A0(\w[3][22] ),
    .A1(\w[1][22] ),
    .A2(\w[7][22] ),
    .A3(\w[5][22] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10362_));
 sky130_fd_sc_hd__mux4_1 _24714_ (.A0(\w[11][22] ),
    .A1(\w[9][22] ),
    .A2(\w[15][22] ),
    .A3(\w[13][22] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10363_));
 sky130_fd_sc_hd__mux4_1 _24715_ (.A0(_10360_),
    .A1(_10361_),
    .A2(_10362_),
    .A3(_10363_),
    .S0(net517),
    .S1(net512),
    .X(_10364_));
 sky130_fd_sc_hd__mux4_1 _24716_ (.A0(\w[51][22] ),
    .A1(\w[49][22] ),
    .A2(\w[55][22] ),
    .A3(\w[53][22] ),
    .S0(net544),
    .S1(net488),
    .X(_10365_));
 sky130_fd_sc_hd__mux4_1 _24717_ (.A0(\w[59][22] ),
    .A1(\w[57][22] ),
    .A2(\w[63][22] ),
    .A3(\w[61][22] ),
    .S0(net544),
    .S1(net488),
    .X(_10366_));
 sky130_fd_sc_hd__mux4_1 _24718_ (.A0(\w[35][22] ),
    .A1(\w[33][22] ),
    .A2(\w[39][22] ),
    .A3(\w[37][22] ),
    .S0(net544),
    .S1(net488),
    .X(_10367_));
 sky130_fd_sc_hd__mux4_1 _24719_ (.A0(\w[43][22] ),
    .A1(\w[41][22] ),
    .A2(\w[47][22] ),
    .A3(\w[45][22] ),
    .S0(net544),
    .S1(net488),
    .X(_10368_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_511 ();
 sky130_fd_sc_hd__mux4_2 _24722_ (.A0(_10365_),
    .A1(_10366_),
    .A2(_10367_),
    .A3(_10368_),
    .S0(net516),
    .S1(net511),
    .X(_10371_));
 sky130_fd_sc_hd__mux2i_1 _24723_ (.A0(_10364_),
    .A1(_10371_),
    .S(net466),
    .Y(_10372_));
 sky130_fd_sc_hd__nand2_1 _24724_ (.A(reset_hash),
    .B(\w[1][22] ),
    .Y(_10373_));
 sky130_fd_sc_hd__o21ai_0 _24725_ (.A1(net454),
    .A2(_10372_),
    .B1(_10373_),
    .Y(_00046_));
 sky130_fd_sc_hd__mux4_1 _24726_ (.A0(\w[19][23] ),
    .A1(\w[17][23] ),
    .A2(\w[23][23] ),
    .A3(\w[21][23] ),
    .S0(net539),
    .S1(net484),
    .X(_10374_));
 sky130_fd_sc_hd__mux4_1 _24727_ (.A0(\w[27][23] ),
    .A1(\w[25][23] ),
    .A2(\w[31][23] ),
    .A3(\w[29][23] ),
    .S0(net539),
    .S1(net484),
    .X(_10375_));
 sky130_fd_sc_hd__mux4_1 _24728_ (.A0(\w[3][23] ),
    .A1(\w[1][23] ),
    .A2(\w[7][23] ),
    .A3(\w[5][23] ),
    .S0(net539),
    .S1(net484),
    .X(_10376_));
 sky130_fd_sc_hd__mux4_1 _24729_ (.A0(\w[11][23] ),
    .A1(\w[9][23] ),
    .A2(\w[15][23] ),
    .A3(\w[13][23] ),
    .S0(net539),
    .S1(net484),
    .X(_10377_));
 sky130_fd_sc_hd__mux4_1 _24730_ (.A0(_10374_),
    .A1(_10375_),
    .A2(_10376_),
    .A3(_10377_),
    .S0(net516),
    .S1(net511),
    .X(_10378_));
 sky130_fd_sc_hd__mux4_1 _24731_ (.A0(\w[51][23] ),
    .A1(\w[49][23] ),
    .A2(\w[55][23] ),
    .A3(\w[53][23] ),
    .S0(net543),
    .S1(net487),
    .X(_10379_));
 sky130_fd_sc_hd__mux4_1 _24732_ (.A0(\w[59][23] ),
    .A1(\w[57][23] ),
    .A2(\w[63][23] ),
    .A3(\w[61][23] ),
    .S0(net543),
    .S1(net487),
    .X(_10380_));
 sky130_fd_sc_hd__mux4_1 _24733_ (.A0(\w[35][23] ),
    .A1(\w[33][23] ),
    .A2(\w[39][23] ),
    .A3(\w[37][23] ),
    .S0(net543),
    .S1(net487),
    .X(_10381_));
 sky130_fd_sc_hd__mux4_1 _24734_ (.A0(\w[43][23] ),
    .A1(\w[41][23] ),
    .A2(\w[47][23] ),
    .A3(\w[45][23] ),
    .S0(net543),
    .S1(net487),
    .X(_10382_));
 sky130_fd_sc_hd__mux4_2 _24735_ (.A0(_10379_),
    .A1(_10380_),
    .A2(_10381_),
    .A3(_10382_),
    .S0(net514),
    .S1(net509),
    .X(_10383_));
 sky130_fd_sc_hd__mux2i_2 _24736_ (.A0(_10378_),
    .A1(_10383_),
    .S(net465),
    .Y(_10384_));
 sky130_fd_sc_hd__nand2_1 _24737_ (.A(reset_hash),
    .B(\w[1][23] ),
    .Y(_10385_));
 sky130_fd_sc_hd__o21ai_4 _24738_ (.A1(net454),
    .A2(_10384_),
    .B1(_10385_),
    .Y(_00047_));
 sky130_fd_sc_hd__mux4_1 _24739_ (.A0(\w[19][24] ),
    .A1(\w[17][24] ),
    .A2(\w[23][24] ),
    .A3(\w[21][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10386_));
 sky130_fd_sc_hd__mux4_1 _24740_ (.A0(\w[27][24] ),
    .A1(\w[25][24] ),
    .A2(\w[31][24] ),
    .A3(\w[29][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10387_));
 sky130_fd_sc_hd__mux4_1 _24741_ (.A0(\w[3][24] ),
    .A1(\w[1][24] ),
    .A2(\w[7][24] ),
    .A3(\w[5][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10388_));
 sky130_fd_sc_hd__mux4_1 _24742_ (.A0(\w[11][24] ),
    .A1(\w[9][24] ),
    .A2(\w[15][24] ),
    .A3(\w[13][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10389_));
 sky130_fd_sc_hd__mux4_1 _24743_ (.A0(_10386_),
    .A1(_10387_),
    .A2(_10388_),
    .A3(_10389_),
    .S0(net514),
    .S1(net509),
    .X(_10390_));
 sky130_fd_sc_hd__mux4_1 _24744_ (.A0(\w[51][24] ),
    .A1(\w[49][24] ),
    .A2(\w[55][24] ),
    .A3(\w[53][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10391_));
 sky130_fd_sc_hd__mux4_1 _24745_ (.A0(\w[59][24] ),
    .A1(\w[57][24] ),
    .A2(\w[63][24] ),
    .A3(\w[61][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10392_));
 sky130_fd_sc_hd__mux4_1 _24746_ (.A0(\w[35][24] ),
    .A1(\w[33][24] ),
    .A2(\w[39][24] ),
    .A3(\w[37][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10393_));
 sky130_fd_sc_hd__mux4_1 _24747_ (.A0(\w[43][24] ),
    .A1(\w[41][24] ),
    .A2(\w[47][24] ),
    .A3(\w[45][24] ),
    .S0(net542),
    .S1(net487),
    .X(_10394_));
 sky130_fd_sc_hd__mux4_1 _24748_ (.A0(_10391_),
    .A1(_10392_),
    .A2(_10393_),
    .A3(_10394_),
    .S0(net514),
    .S1(net509),
    .X(_10395_));
 sky130_fd_sc_hd__mux2i_2 _24749_ (.A0(_10390_),
    .A1(_10395_),
    .S(net464),
    .Y(_10396_));
 sky130_fd_sc_hd__nand2_1 _24750_ (.A(reset_hash),
    .B(\w[1][24] ),
    .Y(_10397_));
 sky130_fd_sc_hd__o21ai_4 _24751_ (.A1(net454),
    .A2(_10396_),
    .B1(_10397_),
    .Y(_00048_));
 sky130_fd_sc_hd__mux4_1 _24752_ (.A0(\w[19][25] ),
    .A1(\w[17][25] ),
    .A2(\w[23][25] ),
    .A3(\w[21][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10398_));
 sky130_fd_sc_hd__mux4_1 _24753_ (.A0(\w[27][25] ),
    .A1(\w[25][25] ),
    .A2(\w[31][25] ),
    .A3(\w[29][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10399_));
 sky130_fd_sc_hd__mux4_1 _24754_ (.A0(\w[3][25] ),
    .A1(\w[1][25] ),
    .A2(\w[7][25] ),
    .A3(\w[5][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10400_));
 sky130_fd_sc_hd__mux4_1 _24755_ (.A0(\w[11][25] ),
    .A1(\w[9][25] ),
    .A2(\w[15][25] ),
    .A3(\w[13][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10401_));
 sky130_fd_sc_hd__mux4_1 _24756_ (.A0(_10398_),
    .A1(_10399_),
    .A2(_10400_),
    .A3(_10401_),
    .S0(net514),
    .S1(net509),
    .X(_10402_));
 sky130_fd_sc_hd__mux4_1 _24757_ (.A0(\w[51][25] ),
    .A1(\w[49][25] ),
    .A2(\w[55][25] ),
    .A3(\w[53][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10403_));
 sky130_fd_sc_hd__mux4_1 _24758_ (.A0(\w[59][25] ),
    .A1(\w[57][25] ),
    .A2(\w[63][25] ),
    .A3(\w[61][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10404_));
 sky130_fd_sc_hd__mux4_1 _24759_ (.A0(\w[35][25] ),
    .A1(\w[33][25] ),
    .A2(\w[39][25] ),
    .A3(\w[37][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10405_));
 sky130_fd_sc_hd__mux4_1 _24760_ (.A0(\w[43][25] ),
    .A1(\w[41][25] ),
    .A2(\w[47][25] ),
    .A3(\w[45][25] ),
    .S0(net542),
    .S1(net487),
    .X(_10406_));
 sky130_fd_sc_hd__mux4_2 _24761_ (.A0(_10403_),
    .A1(_10404_),
    .A2(_10405_),
    .A3(_10406_),
    .S0(net514),
    .S1(net509),
    .X(_10407_));
 sky130_fd_sc_hd__mux2i_2 _24762_ (.A0(_10402_),
    .A1(_10407_),
    .S(net464),
    .Y(_10408_));
 sky130_fd_sc_hd__nand2_1 _24763_ (.A(reset_hash),
    .B(\w[1][25] ),
    .Y(_10409_));
 sky130_fd_sc_hd__o21ai_4 _24764_ (.A1(net454),
    .A2(_10408_),
    .B1(_10409_),
    .Y(_00049_));
 sky130_fd_sc_hd__mux4_1 _24765_ (.A0(\w[19][26] ),
    .A1(\w[17][26] ),
    .A2(\w[23][26] ),
    .A3(\w[21][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10410_));
 sky130_fd_sc_hd__mux4_1 _24766_ (.A0(\w[27][26] ),
    .A1(\w[25][26] ),
    .A2(\w[31][26] ),
    .A3(\w[29][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10411_));
 sky130_fd_sc_hd__mux4_1 _24767_ (.A0(\w[3][26] ),
    .A1(\w[1][26] ),
    .A2(\w[7][26] ),
    .A3(\w[5][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10412_));
 sky130_fd_sc_hd__mux4_1 _24768_ (.A0(\w[11][26] ),
    .A1(\w[9][26] ),
    .A2(\w[15][26] ),
    .A3(\w[13][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10413_));
 sky130_fd_sc_hd__mux4_1 _24769_ (.A0(_10410_),
    .A1(_10411_),
    .A2(_10412_),
    .A3(_10413_),
    .S0(net516),
    .S1(net511),
    .X(_10414_));
 sky130_fd_sc_hd__mux4_1 _24770_ (.A0(\w[51][26] ),
    .A1(\w[49][26] ),
    .A2(\w[55][26] ),
    .A3(\w[53][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10415_));
 sky130_fd_sc_hd__mux4_1 _24771_ (.A0(\w[59][26] ),
    .A1(\w[57][26] ),
    .A2(\w[63][26] ),
    .A3(\w[61][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10416_));
 sky130_fd_sc_hd__mux4_1 _24772_ (.A0(\w[35][26] ),
    .A1(\w[33][26] ),
    .A2(\w[39][26] ),
    .A3(\w[37][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10417_));
 sky130_fd_sc_hd__mux4_1 _24773_ (.A0(\w[43][26] ),
    .A1(\w[41][26] ),
    .A2(\w[47][26] ),
    .A3(\w[45][26] ),
    .S0(net539),
    .S1(net484),
    .X(_10418_));
 sky130_fd_sc_hd__mux4_2 _24774_ (.A0(_10415_),
    .A1(_10416_),
    .A2(_10417_),
    .A3(_10418_),
    .S0(net516),
    .S1(net511),
    .X(_10419_));
 sky130_fd_sc_hd__mux2i_2 _24775_ (.A0(_10414_),
    .A1(_10419_),
    .S(net465),
    .Y(_10420_));
 sky130_fd_sc_hd__nand2_1 _24776_ (.A(reset_hash),
    .B(\w[1][26] ),
    .Y(_10421_));
 sky130_fd_sc_hd__o21ai_4 _24777_ (.A1(net454),
    .A2(_10420_),
    .B1(_10421_),
    .Y(_00050_));
 sky130_fd_sc_hd__mux4_1 _24778_ (.A0(\w[19][27] ),
    .A1(\w[17][27] ),
    .A2(\w[23][27] ),
    .A3(\w[21][27] ),
    .S0(net539),
    .S1(net484),
    .X(_10422_));
 sky130_fd_sc_hd__mux4_1 _24779_ (.A0(\w[27][27] ),
    .A1(\w[25][27] ),
    .A2(\w[31][27] ),
    .A3(\w[29][27] ),
    .S0(net539),
    .S1(net484),
    .X(_10423_));
 sky130_fd_sc_hd__mux4_1 _24780_ (.A0(\w[3][27] ),
    .A1(\w[1][27] ),
    .A2(\w[7][27] ),
    .A3(\w[5][27] ),
    .S0(net539),
    .S1(net484),
    .X(_10424_));
 sky130_fd_sc_hd__mux4_1 _24781_ (.A0(\w[11][27] ),
    .A1(\w[9][27] ),
    .A2(\w[15][27] ),
    .A3(\w[13][27] ),
    .S0(net539),
    .S1(net484),
    .X(_10425_));
 sky130_fd_sc_hd__mux4_1 _24782_ (.A0(_10422_),
    .A1(_10423_),
    .A2(_10424_),
    .A3(_10425_),
    .S0(net516),
    .S1(net511),
    .X(_10426_));
 sky130_fd_sc_hd__mux4_1 _24783_ (.A0(\w[51][27] ),
    .A1(\w[49][27] ),
    .A2(\w[55][27] ),
    .A3(\w[53][27] ),
    .S0(net543),
    .S1(net487),
    .X(_10427_));
 sky130_fd_sc_hd__mux4_1 _24784_ (.A0(\w[59][27] ),
    .A1(\w[57][27] ),
    .A2(\w[63][27] ),
    .A3(\w[61][27] ),
    .S0(net543),
    .S1(net487),
    .X(_10428_));
 sky130_fd_sc_hd__mux4_1 _24785_ (.A0(\w[35][27] ),
    .A1(\w[33][27] ),
    .A2(\w[39][27] ),
    .A3(\w[37][27] ),
    .S0(net543),
    .S1(net487),
    .X(_10429_));
 sky130_fd_sc_hd__mux4_1 _24786_ (.A0(\w[43][27] ),
    .A1(\w[41][27] ),
    .A2(\w[47][27] ),
    .A3(\w[45][27] ),
    .S0(net543),
    .S1(net487),
    .X(_10430_));
 sky130_fd_sc_hd__mux4_4 _24787_ (.A0(_10427_),
    .A1(_10428_),
    .A2(_10429_),
    .A3(_10430_),
    .S0(net514),
    .S1(net509),
    .X(_10431_));
 sky130_fd_sc_hd__mux2i_2 _24788_ (.A0(_10426_),
    .A1(_10431_),
    .S(net464),
    .Y(_10432_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_510 ();
 sky130_fd_sc_hd__nand2_1 _24790_ (.A(reset_hash),
    .B(\w[1][27] ),
    .Y(_10434_));
 sky130_fd_sc_hd__o21ai_4 _24791_ (.A1(net454),
    .A2(_10432_),
    .B1(_10434_),
    .Y(_00051_));
 sky130_fd_sc_hd__mux4_1 _24792_ (.A0(\w[19][28] ),
    .A1(\w[17][28] ),
    .A2(\w[23][28] ),
    .A3(\w[21][28] ),
    .S0(net544),
    .S1(net488),
    .X(_10435_));
 sky130_fd_sc_hd__mux4_1 _24793_ (.A0(\w[27][28] ),
    .A1(\w[25][28] ),
    .A2(\w[31][28] ),
    .A3(\w[29][28] ),
    .S0(net544),
    .S1(net488),
    .X(_10436_));
 sky130_fd_sc_hd__mux4_1 _24794_ (.A0(\w[3][28] ),
    .A1(\w[1][28] ),
    .A2(\w[7][28] ),
    .A3(\w[5][28] ),
    .S0(net544),
    .S1(net488),
    .X(_10437_));
 sky130_fd_sc_hd__mux4_1 _24795_ (.A0(\w[11][28] ),
    .A1(\w[9][28] ),
    .A2(\w[15][28] ),
    .A3(\w[13][28] ),
    .S0(net544),
    .S1(net488),
    .X(_10438_));
 sky130_fd_sc_hd__mux4_1 _24796_ (.A0(_10435_),
    .A1(_10436_),
    .A2(_10437_),
    .A3(_10438_),
    .S0(net517),
    .S1(net512),
    .X(_10439_));
 sky130_fd_sc_hd__mux4_1 _24797_ (.A0(\w[51][28] ),
    .A1(\w[49][28] ),
    .A2(\w[55][28] ),
    .A3(\w[53][28] ),
    .S0(net539),
    .S1(net484),
    .X(_10440_));
 sky130_fd_sc_hd__mux4_1 _24798_ (.A0(\w[59][28] ),
    .A1(\w[57][28] ),
    .A2(\w[63][28] ),
    .A3(\w[61][28] ),
    .S0(net539),
    .S1(net484),
    .X(_10441_));
 sky130_fd_sc_hd__mux4_1 _24799_ (.A0(\w[35][28] ),
    .A1(\w[33][28] ),
    .A2(\w[39][28] ),
    .A3(\w[37][28] ),
    .S0(net539),
    .S1(net484),
    .X(_10442_));
 sky130_fd_sc_hd__mux4_1 _24800_ (.A0(\w[43][28] ),
    .A1(\w[41][28] ),
    .A2(\w[47][28] ),
    .A3(\w[45][28] ),
    .S0(net539),
    .S1(net484),
    .X(_10443_));
 sky130_fd_sc_hd__mux4_4 _24801_ (.A0(_10440_),
    .A1(_10441_),
    .A2(_10442_),
    .A3(_10443_),
    .S0(net516),
    .S1(net511),
    .X(_10444_));
 sky130_fd_sc_hd__mux2i_1 _24802_ (.A0(_10439_),
    .A1(_10444_),
    .S(net465),
    .Y(_10445_));
 sky130_fd_sc_hd__nand2_1 _24803_ (.A(reset_hash),
    .B(\w[1][28] ),
    .Y(_10446_));
 sky130_fd_sc_hd__o21ai_2 _24804_ (.A1(net454),
    .A2(_10445_),
    .B1(_10446_),
    .Y(_00052_));
 sky130_fd_sc_hd__mux4_1 _24805_ (.A0(\w[19][29] ),
    .A1(\w[17][29] ),
    .A2(\w[23][29] ),
    .A3(\w[21][29] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10447_));
 sky130_fd_sc_hd__mux4_1 _24806_ (.A0(\w[27][29] ),
    .A1(\w[25][29] ),
    .A2(\w[31][29] ),
    .A3(\w[29][29] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10448_));
 sky130_fd_sc_hd__mux4_1 _24807_ (.A0(\w[3][29] ),
    .A1(\w[1][29] ),
    .A2(\w[7][29] ),
    .A3(\w[5][29] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10449_));
 sky130_fd_sc_hd__mux4_1 _24808_ (.A0(\w[11][29] ),
    .A1(\w[9][29] ),
    .A2(\w[15][29] ),
    .A3(\w[13][29] ),
    .S0(net545),
    .S1(_00657_),
    .X(_10450_));
 sky130_fd_sc_hd__mux4_1 _24809_ (.A0(_10447_),
    .A1(_10448_),
    .A2(_10449_),
    .A3(_10450_),
    .S0(net517),
    .S1(net512),
    .X(_10451_));
 sky130_fd_sc_hd__mux4_1 _24810_ (.A0(\w[51][29] ),
    .A1(\w[49][29] ),
    .A2(\w[55][29] ),
    .A3(\w[53][29] ),
    .S0(net544),
    .S1(net488),
    .X(_10452_));
 sky130_fd_sc_hd__mux4_1 _24811_ (.A0(\w[59][29] ),
    .A1(\w[57][29] ),
    .A2(\w[63][29] ),
    .A3(\w[61][29] ),
    .S0(net544),
    .S1(net488),
    .X(_10453_));
 sky130_fd_sc_hd__mux4_1 _24812_ (.A0(\w[35][29] ),
    .A1(\w[33][29] ),
    .A2(\w[39][29] ),
    .A3(\w[37][29] ),
    .S0(net544),
    .S1(net488),
    .X(_10454_));
 sky130_fd_sc_hd__mux4_1 _24813_ (.A0(\w[43][29] ),
    .A1(\w[41][29] ),
    .A2(\w[47][29] ),
    .A3(\w[45][29] ),
    .S0(net544),
    .S1(net488),
    .X(_10455_));
 sky130_fd_sc_hd__mux4_2 _24814_ (.A0(_10452_),
    .A1(_10453_),
    .A2(_10454_),
    .A3(_10455_),
    .S0(net516),
    .S1(net511),
    .X(_10456_));
 sky130_fd_sc_hd__mux2i_1 _24815_ (.A0(_10451_),
    .A1(_10456_),
    .S(net466),
    .Y(_10457_));
 sky130_fd_sc_hd__nand2_1 _24816_ (.A(reset_hash),
    .B(\w[1][29] ),
    .Y(_10458_));
 sky130_fd_sc_hd__o21ai_0 _24817_ (.A1(net454),
    .A2(_10457_),
    .B1(_10458_),
    .Y(_00053_));
 sky130_fd_sc_hd__mux4_1 _24818_ (.A0(\w[19][30] ),
    .A1(\w[17][30] ),
    .A2(\w[23][30] ),
    .A3(\w[21][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10459_));
 sky130_fd_sc_hd__mux4_1 _24819_ (.A0(\w[27][30] ),
    .A1(\w[25][30] ),
    .A2(\w[31][30] ),
    .A3(\w[29][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10460_));
 sky130_fd_sc_hd__mux4_1 _24820_ (.A0(\w[3][30] ),
    .A1(\w[1][30] ),
    .A2(\w[7][30] ),
    .A3(\w[5][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10461_));
 sky130_fd_sc_hd__mux4_1 _24821_ (.A0(\w[11][30] ),
    .A1(\w[9][30] ),
    .A2(\w[15][30] ),
    .A3(\w[13][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10462_));
 sky130_fd_sc_hd__mux4_1 _24822_ (.A0(_10459_),
    .A1(_10460_),
    .A2(_10461_),
    .A3(_10462_),
    .S0(net517),
    .S1(net512),
    .X(_10463_));
 sky130_fd_sc_hd__mux4_1 _24823_ (.A0(\w[51][30] ),
    .A1(\w[49][30] ),
    .A2(\w[55][30] ),
    .A3(\w[53][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10464_));
 sky130_fd_sc_hd__mux4_1 _24824_ (.A0(\w[59][30] ),
    .A1(\w[57][30] ),
    .A2(\w[63][30] ),
    .A3(\w[61][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10465_));
 sky130_fd_sc_hd__mux4_1 _24825_ (.A0(\w[35][30] ),
    .A1(\w[33][30] ),
    .A2(\w[39][30] ),
    .A3(\w[37][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10466_));
 sky130_fd_sc_hd__mux4_1 _24826_ (.A0(\w[43][30] ),
    .A1(\w[41][30] ),
    .A2(\w[47][30] ),
    .A3(\w[45][30] ),
    .S0(net544),
    .S1(net488),
    .X(_10467_));
 sky130_fd_sc_hd__mux4_1 _24827_ (.A0(_10464_),
    .A1(_10465_),
    .A2(_10466_),
    .A3(_10467_),
    .S0(net517),
    .S1(net512),
    .X(_10468_));
 sky130_fd_sc_hd__mux2i_1 _24828_ (.A0(_10463_),
    .A1(_10468_),
    .S(net465),
    .Y(_10469_));
 sky130_fd_sc_hd__nand2_1 _24829_ (.A(reset_hash),
    .B(\w[1][30] ),
    .Y(_10470_));
 sky130_fd_sc_hd__o21ai_2 _24830_ (.A1(net454),
    .A2(_10469_),
    .B1(_10470_),
    .Y(_00055_));
 sky130_fd_sc_hd__mux4_1 _24831_ (.A0(\w[19][31] ),
    .A1(\w[17][31] ),
    .A2(\w[23][31] ),
    .A3(\w[21][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10471_));
 sky130_fd_sc_hd__mux4_1 _24832_ (.A0(\w[27][31] ),
    .A1(\w[25][31] ),
    .A2(\w[31][31] ),
    .A3(\w[29][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10472_));
 sky130_fd_sc_hd__mux4_1 _24833_ (.A0(\w[3][31] ),
    .A1(\w[1][31] ),
    .A2(\w[7][31] ),
    .A3(\w[5][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10473_));
 sky130_fd_sc_hd__mux4_1 _24834_ (.A0(\w[11][31] ),
    .A1(\w[9][31] ),
    .A2(\w[15][31] ),
    .A3(\w[13][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10474_));
 sky130_fd_sc_hd__mux4_1 _24835_ (.A0(_10471_),
    .A1(_10472_),
    .A2(_10473_),
    .A3(_10474_),
    .S0(net516),
    .S1(net511),
    .X(_10475_));
 sky130_fd_sc_hd__mux4_1 _24836_ (.A0(\w[51][31] ),
    .A1(\w[49][31] ),
    .A2(\w[55][31] ),
    .A3(\w[53][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10476_));
 sky130_fd_sc_hd__mux4_1 _24837_ (.A0(\w[59][31] ),
    .A1(\w[57][31] ),
    .A2(\w[63][31] ),
    .A3(\w[61][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10477_));
 sky130_fd_sc_hd__mux4_1 _24838_ (.A0(\w[35][31] ),
    .A1(\w[33][31] ),
    .A2(\w[39][31] ),
    .A3(\w[37][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10478_));
 sky130_fd_sc_hd__mux4_1 _24839_ (.A0(\w[43][31] ),
    .A1(\w[41][31] ),
    .A2(\w[47][31] ),
    .A3(\w[45][31] ),
    .S0(net539),
    .S1(net484),
    .X(_10479_));
 sky130_fd_sc_hd__mux4_2 _24840_ (.A0(_10476_),
    .A1(_10477_),
    .A2(_10478_),
    .A3(_10479_),
    .S0(net516),
    .S1(net511),
    .X(_10480_));
 sky130_fd_sc_hd__mux2i_2 _24841_ (.A0(_10475_),
    .A1(_10480_),
    .S(net465),
    .Y(_10481_));
 sky130_fd_sc_hd__nand2_1 _24842_ (.A(reset_hash),
    .B(\w[1][31] ),
    .Y(_10482_));
 sky130_fd_sc_hd__o21ai_4 _24843_ (.A1(net454),
    .A2(_10481_),
    .B1(_10482_),
    .Y(_00056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_503 ();
 sky130_fd_sc_hd__mux4_1 _24851_ (.A0(\w[18][0] ),
    .A1(\w[16][0] ),
    .A2(\w[22][0] ),
    .A3(\w[20][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_501 ();
 sky130_fd_sc_hd__mux4_1 _24854_ (.A0(\w[26][0] ),
    .A1(\w[24][0] ),
    .A2(\w[30][0] ),
    .A3(\w[28][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10493_));
 sky130_fd_sc_hd__mux4_1 _24855_ (.A0(\w[2][0] ),
    .A1(\w[0][0] ),
    .A2(\w[6][0] ),
    .A3(\w[4][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_498 ();
 sky130_fd_sc_hd__mux4_1 _24859_ (.A0(\w[10][0] ),
    .A1(\w[8][0] ),
    .A2(\w[14][0] ),
    .A3(\w[12][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10498_));
 sky130_fd_sc_hd__xor2_4 _24860_ (.A(\count_hash1[3] ),
    .B(_13088_),
    .X(_10499_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_496 ();
 sky130_fd_sc_hd__nand3_4 _24863_ (.A(\count_hash1[3] ),
    .B(\count_hash1[2] ),
    .C(\count_hash1[1] ),
    .Y(_10502_));
 sky130_fd_sc_hd__xor2_4 _24864_ (.A(\count_hash1[4] ),
    .B(_10502_),
    .X(_10503_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_494 ();
 sky130_fd_sc_hd__mux4_1 _24867_ (.A0(_10490_),
    .A1(_10493_),
    .A2(_10494_),
    .A3(_10498_),
    .S0(net505),
    .S1(net497),
    .X(_10506_));
 sky130_fd_sc_hd__nand3_4 _24868_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(_13088_),
    .Y(_10507_));
 sky130_fd_sc_hd__xor2_4 _24869_ (.A(\count_hash1[5] ),
    .B(_10507_),
    .X(_10508_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_491 ();
 sky130_fd_sc_hd__xnor2_4 _24873_ (.A(\count_hash1[4] ),
    .B(_10502_),
    .Y(_10512_));
 sky130_fd_sc_hd__nor2_8 _24874_ (.A(_10512_),
    .B(net507),
    .Y(_10513_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_484 ();
 sky130_fd_sc_hd__mux4_1 _24882_ (.A0(\w[34][0] ),
    .A1(\w[32][0] ),
    .A2(\w[38][0] ),
    .A3(\w[36][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10521_));
 sky130_fd_sc_hd__nand2_1 _24883_ (.A(net460),
    .B(_10521_),
    .Y(_10522_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_476 ();
 sky130_fd_sc_hd__mux4_1 _24892_ (.A0(\w[42][0] ),
    .A1(\w[40][0] ),
    .A2(\w[46][0] ),
    .A3(\w[44][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10531_));
 sky130_fd_sc_hd__xnor2_4 _24893_ (.A(\count_hash1[3] ),
    .B(_13088_),
    .Y(_10532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_474 ();
 sky130_fd_sc_hd__mux4_1 _24896_ (.A0(\w[50][0] ),
    .A1(\w[48][0] ),
    .A2(\w[54][0] ),
    .A3(\w[52][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10535_));
 sky130_fd_sc_hd__nand2_1 _24897_ (.A(net491),
    .B(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_471 ();
 sky130_fd_sc_hd__mux4_1 _24901_ (.A0(\w[58][0] ),
    .A1(\w[56][0] ),
    .A2(\w[62][0] ),
    .A3(\w[60][0] ),
    .S0(net547),
    .S1(net481),
    .X(_10540_));
 sky130_fd_sc_hd__nand2_1 _24902_ (.A(net505),
    .B(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_470 ();
 sky130_fd_sc_hd__a21oi_1 _24904_ (.A1(_10536_),
    .A2(_10541_),
    .B1(net498),
    .Y(_10543_));
 sky130_fd_sc_hd__a31oi_1 _24905_ (.A1(net498),
    .A2(net505),
    .A3(_10531_),
    .B1(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__a21oi_1 _24906_ (.A1(_10522_),
    .A2(_10544_),
    .B1(net462),
    .Y(_10545_));
 sky130_fd_sc_hd__a21oi_1 _24907_ (.A1(_10506_),
    .A2(net462),
    .B1(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__nand2_1 _24908_ (.A(net526),
    .B(\w[0][0] ),
    .Y(_10547_));
 sky130_fd_sc_hd__o21ai_4 _24909_ (.A1(net455),
    .A2(_10546_),
    .B1(_10547_),
    .Y(_00000_));
 sky130_fd_sc_hd__mux4_1 _24910_ (.A0(\w[18][1] ),
    .A1(\w[16][1] ),
    .A2(\w[22][1] ),
    .A3(\w[20][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10548_));
 sky130_fd_sc_hd__mux4_1 _24911_ (.A0(\w[26][1] ),
    .A1(\w[24][1] ),
    .A2(\w[30][1] ),
    .A3(\w[28][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10549_));
 sky130_fd_sc_hd__mux4_1 _24912_ (.A0(\w[2][1] ),
    .A1(\w[0][1] ),
    .A2(\w[6][1] ),
    .A3(\w[4][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10550_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_469 ();
 sky130_fd_sc_hd__mux4_1 _24914_ (.A0(\w[10][1] ),
    .A1(\w[8][1] ),
    .A2(\w[14][1] ),
    .A3(\w[12][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10552_));
 sky130_fd_sc_hd__mux4_2 _24915_ (.A0(_10548_),
    .A1(_10549_),
    .A2(_10550_),
    .A3(_10552_),
    .S0(net502),
    .S1(net497),
    .X(_10553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_467 ();
 sky130_fd_sc_hd__mux4_1 _24918_ (.A0(\w[50][1] ),
    .A1(\w[48][1] ),
    .A2(\w[54][1] ),
    .A3(\w[52][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_466 ();
 sky130_fd_sc_hd__mux4_1 _24920_ (.A0(\w[58][1] ),
    .A1(\w[56][1] ),
    .A2(\w[62][1] ),
    .A3(\w[60][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10558_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_465 ();
 sky130_fd_sc_hd__mux4_1 _24922_ (.A0(\w[34][1] ),
    .A1(\w[32][1] ),
    .A2(\w[38][1] ),
    .A3(\w[36][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10560_));
 sky130_fd_sc_hd__mux4_1 _24923_ (.A0(\w[42][1] ),
    .A1(\w[40][1] ),
    .A2(\w[46][1] ),
    .A3(\w[44][1] ),
    .S0(net551),
    .S1(net479),
    .X(_10561_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_464 ();
 sky130_fd_sc_hd__mux4_2 _24925_ (.A0(_10556_),
    .A1(_10558_),
    .A2(_10560_),
    .A3(_10561_),
    .S0(net502),
    .S1(net498),
    .X(_10563_));
 sky130_fd_sc_hd__xnor2_4 _24926_ (.A(\count_hash1[5] ),
    .B(_10507_),
    .Y(_10564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_461 ();
 sky130_fd_sc_hd__mux2i_2 _24930_ (.A0(_10553_),
    .A1(_10563_),
    .S(net457),
    .Y(_10568_));
 sky130_fd_sc_hd__nand2_1 _24931_ (.A(net526),
    .B(\w[0][1] ),
    .Y(_10569_));
 sky130_fd_sc_hd__o21ai_4 _24932_ (.A1(net455),
    .A2(_10568_),
    .B1(_10569_),
    .Y(_00011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_460 ();
 sky130_fd_sc_hd__or2_4 _24934_ (.A(\count_hash1[6] ),
    .B(_10034_),
    .X(_10571_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_459 ();
 sky130_fd_sc_hd__nor2_8 _24936_ (.A(net525),
    .B(_10571_),
    .Y(_10573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_458 ();
 sky130_fd_sc_hd__nand2_8 _24938_ (.A(net493),
    .B(net490),
    .Y(_10575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_454 ();
 sky130_fd_sc_hd__mux4_1 _24943_ (.A0(\w[2][2] ),
    .A1(\w[0][2] ),
    .A2(\w[6][2] ),
    .A3(\w[4][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10580_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_452 ();
 sky130_fd_sc_hd__mux4_1 _24946_ (.A0(\w[34][2] ),
    .A1(\w[32][2] ),
    .A2(\w[38][2] ),
    .A3(\w[36][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10583_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_451 ();
 sky130_fd_sc_hd__mux2i_1 _24948_ (.A0(_10580_),
    .A1(_10583_),
    .S(net457),
    .Y(_10585_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_447 ();
 sky130_fd_sc_hd__mux4_1 _24953_ (.A0(\w[10][2] ),
    .A1(\w[8][2] ),
    .A2(\w[14][2] ),
    .A3(\w[12][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_444 ();
 sky130_fd_sc_hd__mux4_1 _24957_ (.A0(\w[18][2] ),
    .A1(\w[16][2] ),
    .A2(\w[22][2] ),
    .A3(\w[20][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10594_));
 sky130_fd_sc_hd__nand2_1 _24958_ (.A(net489),
    .B(_10594_),
    .Y(_10595_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_441 ();
 sky130_fd_sc_hd__mux4_1 _24962_ (.A0(\w[26][2] ),
    .A1(\w[24][2] ),
    .A2(\w[30][2] ),
    .A3(\w[28][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10599_));
 sky130_fd_sc_hd__nand2_1 _24963_ (.A(net500),
    .B(_10599_),
    .Y(_10600_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_440 ();
 sky130_fd_sc_hd__a21oi_1 _24965_ (.A1(_10595_),
    .A2(_10600_),
    .B1(net495),
    .Y(_10602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_439 ();
 sky130_fd_sc_hd__a311oi_1 _24967_ (.A1(net495),
    .A2(net500),
    .A3(_10590_),
    .B1(_10602_),
    .C1(net457),
    .Y(_10604_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_435 ();
 sky130_fd_sc_hd__mux4_1 _24972_ (.A0(\w[42][2] ),
    .A1(\w[40][2] ),
    .A2(\w[46][2] ),
    .A3(\w[44][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_432 ();
 sky130_fd_sc_hd__mux4_1 _24976_ (.A0(\w[50][2] ),
    .A1(\w[48][2] ),
    .A2(\w[54][2] ),
    .A3(\w[52][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10613_));
 sky130_fd_sc_hd__nand2_1 _24977_ (.A(net489),
    .B(_10613_),
    .Y(_10614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_431 ();
 sky130_fd_sc_hd__mux4_1 _24979_ (.A0(\w[58][2] ),
    .A1(\w[56][2] ),
    .A2(\w[62][2] ),
    .A3(\w[60][2] ),
    .S0(net552),
    .S1(net483),
    .X(_10616_));
 sky130_fd_sc_hd__nand2_1 _24980_ (.A(net500),
    .B(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_430 ();
 sky130_fd_sc_hd__a21oi_1 _24982_ (.A1(_10614_),
    .A2(_10617_),
    .B1(net495),
    .Y(_10619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_429 ();
 sky130_fd_sc_hd__a311oi_2 _24984_ (.A1(net495),
    .A2(net500),
    .A3(_10609_),
    .B1(_10619_),
    .C1(net462),
    .Y(_10621_));
 sky130_fd_sc_hd__o22ai_1 _24985_ (.A1(_10575_),
    .A2(_10585_),
    .B1(_10604_),
    .B2(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__a22o_2 _24986_ (.A1(net526),
    .A2(\w[0][2] ),
    .B1(_10573_),
    .B2(_10622_),
    .X(_00022_));
 sky130_fd_sc_hd__mux4_1 _24987_ (.A0(\w[2][3] ),
    .A1(\w[0][3] ),
    .A2(\w[6][3] ),
    .A3(\w[4][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_428 ();
 sky130_fd_sc_hd__mux4_1 _24989_ (.A0(\w[34][3] ),
    .A1(\w[32][3] ),
    .A2(\w[38][3] ),
    .A3(\w[36][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10625_));
 sky130_fd_sc_hd__mux2i_1 _24990_ (.A0(_10623_),
    .A1(_10625_),
    .S(net456),
    .Y(_10626_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_427 ();
 sky130_fd_sc_hd__mux4_1 _24992_ (.A0(\w[10][3] ),
    .A1(\w[8][3] ),
    .A2(\w[14][3] ),
    .A3(\w[12][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10628_));
 sky130_fd_sc_hd__mux4_1 _24993_ (.A0(\w[18][3] ),
    .A1(\w[16][3] ),
    .A2(\w[22][3] ),
    .A3(\w[20][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10629_));
 sky130_fd_sc_hd__nand2_1 _24994_ (.A(net491),
    .B(_10629_),
    .Y(_10630_));
 sky130_fd_sc_hd__mux4_1 _24995_ (.A0(\w[26][3] ),
    .A1(\w[24][3] ),
    .A2(\w[30][3] ),
    .A3(\w[28][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10631_));
 sky130_fd_sc_hd__nand2_1 _24996_ (.A(net506),
    .B(_10631_),
    .Y(_10632_));
 sky130_fd_sc_hd__a21oi_1 _24997_ (.A1(_10630_),
    .A2(_10632_),
    .B1(net497),
    .Y(_10633_));
 sky130_fd_sc_hd__a311oi_1 _24998_ (.A1(net497),
    .A2(net506),
    .A3(_10628_),
    .B1(_10633_),
    .C1(net456),
    .Y(_10634_));
 sky130_fd_sc_hd__mux4_1 _24999_ (.A0(\w[42][3] ),
    .A1(\w[40][3] ),
    .A2(\w[46][3] ),
    .A3(\w[44][3] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10635_));
 sky130_fd_sc_hd__mux4_1 _25000_ (.A0(\w[50][3] ),
    .A1(\w[48][3] ),
    .A2(\w[54][3] ),
    .A3(\w[52][3] ),
    .S0(net547),
    .S1(net481),
    .X(_10636_));
 sky130_fd_sc_hd__nand2_1 _25001_ (.A(net491),
    .B(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_426 ();
 sky130_fd_sc_hd__mux4_1 _25003_ (.A0(\w[58][3] ),
    .A1(\w[56][3] ),
    .A2(\w[62][3] ),
    .A3(\w[60][3] ),
    .S0(net547),
    .S1(net481),
    .X(_10639_));
 sky130_fd_sc_hd__nand2_1 _25004_ (.A(net506),
    .B(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__a21oi_2 _25005_ (.A1(_10637_),
    .A2(_10640_),
    .B1(net498),
    .Y(_10641_));
 sky130_fd_sc_hd__a311oi_2 _25006_ (.A1(net497),
    .A2(net506),
    .A3(_10635_),
    .B1(_10641_),
    .C1(net462),
    .Y(_10642_));
 sky130_fd_sc_hd__o22ai_1 _25007_ (.A1(_10575_),
    .A2(_10626_),
    .B1(_10634_),
    .B2(_10642_),
    .Y(_10643_));
 sky130_fd_sc_hd__a22o_2 _25008_ (.A1(net526),
    .A2(\w[0][3] ),
    .B1(_10573_),
    .B2(_10643_),
    .X(_00025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_425 ();
 sky130_fd_sc_hd__mux4_1 _25010_ (.A0(\w[18][4] ),
    .A1(\w[16][4] ),
    .A2(\w[22][4] ),
    .A3(\w[20][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10645_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_424 ();
 sky130_fd_sc_hd__mux4_1 _25012_ (.A0(\w[26][4] ),
    .A1(\w[24][4] ),
    .A2(\w[30][4] ),
    .A3(\w[28][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10647_));
 sky130_fd_sc_hd__mux4_1 _25013_ (.A0(\w[2][4] ),
    .A1(\w[0][4] ),
    .A2(\w[6][4] ),
    .A3(\w[4][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10648_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_422 ();
 sky130_fd_sc_hd__mux4_1 _25016_ (.A0(\w[10][4] ),
    .A1(\w[8][4] ),
    .A2(\w[14][4] ),
    .A3(\w[12][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10651_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_421 ();
 sky130_fd_sc_hd__mux4_1 _25018_ (.A0(_10645_),
    .A1(_10647_),
    .A2(_10648_),
    .A3(_10651_),
    .S0(net505),
    .S1(net498),
    .X(_10653_));
 sky130_fd_sc_hd__mux4_1 _25019_ (.A0(\w[34][4] ),
    .A1(\w[32][4] ),
    .A2(\w[38][4] ),
    .A3(\w[36][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10654_));
 sky130_fd_sc_hd__nand2_1 _25020_ (.A(net460),
    .B(_10654_),
    .Y(_10655_));
 sky130_fd_sc_hd__mux4_1 _25021_ (.A0(\w[42][4] ),
    .A1(\w[40][4] ),
    .A2(\w[46][4] ),
    .A3(\w[44][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10656_));
 sky130_fd_sc_hd__mux4_1 _25022_ (.A0(\w[50][4] ),
    .A1(\w[48][4] ),
    .A2(\w[54][4] ),
    .A3(\w[52][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10657_));
 sky130_fd_sc_hd__nand2_1 _25023_ (.A(net492),
    .B(_10657_),
    .Y(_10658_));
 sky130_fd_sc_hd__mux4_1 _25024_ (.A0(\w[58][4] ),
    .A1(\w[56][4] ),
    .A2(\w[62][4] ),
    .A3(\w[60][4] ),
    .S0(net547),
    .S1(net481),
    .X(_10659_));
 sky130_fd_sc_hd__nand2_1 _25025_ (.A(net506),
    .B(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__a21oi_1 _25026_ (.A1(_10658_),
    .A2(_10660_),
    .B1(net498),
    .Y(_10661_));
 sky130_fd_sc_hd__a31oi_2 _25027_ (.A1(net498),
    .A2(net506),
    .A3(_10656_),
    .B1(_10661_),
    .Y(_10662_));
 sky130_fd_sc_hd__a21oi_1 _25028_ (.A1(_10655_),
    .A2(_10662_),
    .B1(net462),
    .Y(_10663_));
 sky130_fd_sc_hd__a21oi_1 _25029_ (.A1(net462),
    .A2(_10653_),
    .B1(_10663_),
    .Y(_10664_));
 sky130_fd_sc_hd__nand2_1 _25030_ (.A(net526),
    .B(\w[0][4] ),
    .Y(_10665_));
 sky130_fd_sc_hd__o21ai_4 _25031_ (.A1(net455),
    .A2(_10664_),
    .B1(_10665_),
    .Y(_00026_));
 sky130_fd_sc_hd__mux4_1 _25032_ (.A0(\w[18][5] ),
    .A1(\w[16][5] ),
    .A2(\w[22][5] ),
    .A3(\w[20][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10666_));
 sky130_fd_sc_hd__mux4_1 _25033_ (.A0(\w[26][5] ),
    .A1(\w[24][5] ),
    .A2(\w[30][5] ),
    .A3(\w[28][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10667_));
 sky130_fd_sc_hd__mux4_1 _25034_ (.A0(\w[2][5] ),
    .A1(\w[0][5] ),
    .A2(\w[6][5] ),
    .A3(\w[4][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10668_));
 sky130_fd_sc_hd__mux4_1 _25035_ (.A0(\w[10][5] ),
    .A1(\w[8][5] ),
    .A2(\w[14][5] ),
    .A3(\w[12][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10669_));
 sky130_fd_sc_hd__mux4_2 _25036_ (.A0(_10666_),
    .A1(_10667_),
    .A2(_10668_),
    .A3(_10669_),
    .S0(net505),
    .S1(net496),
    .X(_10670_));
 sky130_fd_sc_hd__mux4_1 _25037_ (.A0(\w[50][5] ),
    .A1(\w[48][5] ),
    .A2(\w[54][5] ),
    .A3(\w[52][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10671_));
 sky130_fd_sc_hd__mux4_1 _25038_ (.A0(\w[58][5] ),
    .A1(\w[56][5] ),
    .A2(\w[62][5] ),
    .A3(\w[60][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10672_));
 sky130_fd_sc_hd__mux4_1 _25039_ (.A0(\w[34][5] ),
    .A1(\w[32][5] ),
    .A2(\w[38][5] ),
    .A3(\w[36][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10673_));
 sky130_fd_sc_hd__mux4_1 _25040_ (.A0(\w[42][5] ),
    .A1(\w[40][5] ),
    .A2(\w[46][5] ),
    .A3(\w[44][5] ),
    .S0(net546),
    .S1(net480),
    .X(_10674_));
 sky130_fd_sc_hd__mux4_1 _25041_ (.A0(_10671_),
    .A1(_10672_),
    .A2(_10673_),
    .A3(_10674_),
    .S0(net506),
    .S1(net499),
    .X(_10675_));
 sky130_fd_sc_hd__mux2i_2 _25042_ (.A0(_10670_),
    .A1(_10675_),
    .S(net456),
    .Y(_10676_));
 sky130_fd_sc_hd__nand2_1 _25043_ (.A(net526),
    .B(\w[0][5] ),
    .Y(_10677_));
 sky130_fd_sc_hd__o21ai_4 _25044_ (.A1(net455),
    .A2(_10676_),
    .B1(_10677_),
    .Y(_00027_));
 sky130_fd_sc_hd__mux4_1 _25045_ (.A0(\w[18][6] ),
    .A1(\w[16][6] ),
    .A2(\w[22][6] ),
    .A3(\w[20][6] ),
    .S0(net547),
    .S1(net481),
    .X(_10678_));
 sky130_fd_sc_hd__mux4_1 _25046_ (.A0(\w[26][6] ),
    .A1(\w[24][6] ),
    .A2(\w[30][6] ),
    .A3(\w[28][6] ),
    .S0(net547),
    .S1(net481),
    .X(_10679_));
 sky130_fd_sc_hd__mux4_1 _25047_ (.A0(\w[2][6] ),
    .A1(\w[0][6] ),
    .A2(\w[6][6] ),
    .A3(\w[4][6] ),
    .S0(net547),
    .S1(net481),
    .X(_10680_));
 sky130_fd_sc_hd__mux4_1 _25048_ (.A0(\w[10][6] ),
    .A1(\w[8][6] ),
    .A2(\w[14][6] ),
    .A3(\w[12][6] ),
    .S0(net547),
    .S1(net481),
    .X(_10681_));
 sky130_fd_sc_hd__mux4_2 _25049_ (.A0(_10678_),
    .A1(_10679_),
    .A2(_10680_),
    .A3(_10681_),
    .S0(net505),
    .S1(net498),
    .X(_10682_));
 sky130_fd_sc_hd__mux4_1 _25050_ (.A0(\w[34][6] ),
    .A1(\w[32][6] ),
    .A2(\w[38][6] ),
    .A3(\w[36][6] ),
    .S0(net546),
    .S1(net480),
    .X(_10683_));
 sky130_fd_sc_hd__nand2_1 _25051_ (.A(net460),
    .B(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_420 ();
 sky130_fd_sc_hd__mux4_1 _25053_ (.A0(\w[42][6] ),
    .A1(\w[40][6] ),
    .A2(\w[46][6] ),
    .A3(\w[44][6] ),
    .S0(net546),
    .S1(net480),
    .X(_10686_));
 sky130_fd_sc_hd__mux4_1 _25054_ (.A0(\w[50][6] ),
    .A1(\w[48][6] ),
    .A2(\w[54][6] ),
    .A3(\w[52][6] ),
    .S0(net546),
    .S1(net480),
    .X(_10687_));
 sky130_fd_sc_hd__nand2_1 _25055_ (.A(net492),
    .B(_10687_),
    .Y(_10688_));
 sky130_fd_sc_hd__mux4_1 _25056_ (.A0(\w[58][6] ),
    .A1(\w[56][6] ),
    .A2(\w[62][6] ),
    .A3(\w[60][6] ),
    .S0(net546),
    .S1(net480),
    .X(_10689_));
 sky130_fd_sc_hd__nand2_1 _25057_ (.A(net506),
    .B(_10689_),
    .Y(_10690_));
 sky130_fd_sc_hd__a21oi_1 _25058_ (.A1(_10688_),
    .A2(_10690_),
    .B1(net499),
    .Y(_10691_));
 sky130_fd_sc_hd__a31oi_1 _25059_ (.A1(net499),
    .A2(net506),
    .A3(_10686_),
    .B1(_10691_),
    .Y(_10692_));
 sky130_fd_sc_hd__a21oi_1 _25060_ (.A1(_10684_),
    .A2(_10692_),
    .B1(_10508_),
    .Y(_10693_));
 sky130_fd_sc_hd__a21oi_1 _25061_ (.A1(_10508_),
    .A2(_10682_),
    .B1(_10693_),
    .Y(_10694_));
 sky130_fd_sc_hd__nand2_1 _25062_ (.A(net526),
    .B(\w[0][6] ),
    .Y(_10695_));
 sky130_fd_sc_hd__o21ai_4 _25063_ (.A1(net455),
    .A2(_10694_),
    .B1(_10695_),
    .Y(_00028_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_419 ();
 sky130_fd_sc_hd__mux4_1 _25065_ (.A0(\w[2][7] ),
    .A1(\w[0][7] ),
    .A2(\w[6][7] ),
    .A3(\w[4][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10697_));
 sky130_fd_sc_hd__mux4_1 _25066_ (.A0(\w[34][7] ),
    .A1(\w[32][7] ),
    .A2(\w[38][7] ),
    .A3(\w[36][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10698_));
 sky130_fd_sc_hd__mux2i_1 _25067_ (.A0(_10697_),
    .A1(_10698_),
    .S(net457),
    .Y(_10699_));
 sky130_fd_sc_hd__mux4_1 _25068_ (.A0(\w[10][7] ),
    .A1(\w[8][7] ),
    .A2(\w[14][7] ),
    .A3(\w[12][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10700_));
 sky130_fd_sc_hd__mux4_1 _25069_ (.A0(\w[18][7] ),
    .A1(\w[16][7] ),
    .A2(\w[22][7] ),
    .A3(\w[20][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10701_));
 sky130_fd_sc_hd__nand2_1 _25070_ (.A(net489),
    .B(_10701_),
    .Y(_10702_));
 sky130_fd_sc_hd__mux4_1 _25071_ (.A0(\w[26][7] ),
    .A1(\w[24][7] ),
    .A2(\w[30][7] ),
    .A3(\w[28][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10703_));
 sky130_fd_sc_hd__nand2_1 _25072_ (.A(net500),
    .B(_10703_),
    .Y(_10704_));
 sky130_fd_sc_hd__a21oi_1 _25073_ (.A1(_10702_),
    .A2(_10704_),
    .B1(net495),
    .Y(_10705_));
 sky130_fd_sc_hd__a311oi_1 _25074_ (.A1(net495),
    .A2(net500),
    .A3(_10700_),
    .B1(_10705_),
    .C1(net457),
    .Y(_10706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_418 ();
 sky130_fd_sc_hd__mux4_1 _25076_ (.A0(\w[42][7] ),
    .A1(\w[40][7] ),
    .A2(\w[46][7] ),
    .A3(\w[44][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10708_));
 sky130_fd_sc_hd__mux4_1 _25077_ (.A0(\w[50][7] ),
    .A1(\w[48][7] ),
    .A2(\w[54][7] ),
    .A3(\w[52][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10709_));
 sky130_fd_sc_hd__nand2_1 _25078_ (.A(net489),
    .B(_10709_),
    .Y(_10710_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_417 ();
 sky130_fd_sc_hd__mux4_1 _25080_ (.A0(\w[58][7] ),
    .A1(\w[56][7] ),
    .A2(\w[62][7] ),
    .A3(\w[60][7] ),
    .S0(net552),
    .S1(net483),
    .X(_10712_));
 sky130_fd_sc_hd__nand2_1 _25081_ (.A(net500),
    .B(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_416 ();
 sky130_fd_sc_hd__a21oi_1 _25083_ (.A1(_10710_),
    .A2(_10713_),
    .B1(net495),
    .Y(_10715_));
 sky130_fd_sc_hd__a311oi_1 _25084_ (.A1(net495),
    .A2(net500),
    .A3(_10708_),
    .B1(_10715_),
    .C1(net461),
    .Y(_10716_));
 sky130_fd_sc_hd__o22ai_1 _25085_ (.A1(_10575_),
    .A2(_10699_),
    .B1(_10706_),
    .B2(_10716_),
    .Y(_10717_));
 sky130_fd_sc_hd__a22o_2 _25086_ (.A1(net526),
    .A2(\w[0][7] ),
    .B1(_10573_),
    .B2(_10717_),
    .X(_00029_));
 sky130_fd_sc_hd__mux4_1 _25087_ (.A0(\w[2][8] ),
    .A1(\w[0][8] ),
    .A2(\w[6][8] ),
    .A3(\w[4][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10718_));
 sky130_fd_sc_hd__mux4_1 _25088_ (.A0(\w[34][8] ),
    .A1(\w[32][8] ),
    .A2(\w[38][8] ),
    .A3(\w[36][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10719_));
 sky130_fd_sc_hd__mux2i_1 _25089_ (.A0(_10718_),
    .A1(_10719_),
    .S(net458),
    .Y(_10720_));
 sky130_fd_sc_hd__mux4_2 _25090_ (.A0(\w[10][8] ),
    .A1(\w[8][8] ),
    .A2(\w[14][8] ),
    .A3(\w[12][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10721_));
 sky130_fd_sc_hd__mux4_1 _25091_ (.A0(\w[18][8] ),
    .A1(\w[16][8] ),
    .A2(\w[22][8] ),
    .A3(\w[20][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10722_));
 sky130_fd_sc_hd__nand2_1 _25092_ (.A(net489),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__mux4_1 _25093_ (.A0(\w[26][8] ),
    .A1(\w[24][8] ),
    .A2(\w[30][8] ),
    .A3(\w[28][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10724_));
 sky130_fd_sc_hd__nand2_1 _25094_ (.A(net501),
    .B(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__a21oi_1 _25095_ (.A1(_10723_),
    .A2(_10725_),
    .B1(net494),
    .Y(_10726_));
 sky130_fd_sc_hd__a311oi_1 _25096_ (.A1(net494),
    .A2(net501),
    .A3(_10721_),
    .B1(_10726_),
    .C1(net457),
    .Y(_10727_));
 sky130_fd_sc_hd__mux4_1 _25097_ (.A0(\w[42][8] ),
    .A1(\w[40][8] ),
    .A2(\w[46][8] ),
    .A3(\w[44][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10728_));
 sky130_fd_sc_hd__mux4_1 _25098_ (.A0(\w[50][8] ),
    .A1(\w[48][8] ),
    .A2(\w[54][8] ),
    .A3(\w[52][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10729_));
 sky130_fd_sc_hd__nand2_1 _25099_ (.A(net489),
    .B(_10729_),
    .Y(_10730_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_415 ();
 sky130_fd_sc_hd__mux4_1 _25101_ (.A0(\w[58][8] ),
    .A1(\w[56][8] ),
    .A2(\w[62][8] ),
    .A3(\w[60][8] ),
    .S0(net549),
    .S1(net477),
    .X(_10732_));
 sky130_fd_sc_hd__nand2_1 _25102_ (.A(net503),
    .B(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__a21oi_1 _25103_ (.A1(_10730_),
    .A2(_10733_),
    .B1(net494),
    .Y(_10734_));
 sky130_fd_sc_hd__a311oi_1 _25104_ (.A1(net494),
    .A2(net503),
    .A3(_10728_),
    .B1(_10734_),
    .C1(net461),
    .Y(_10735_));
 sky130_fd_sc_hd__o22ai_1 _25105_ (.A1(_10575_),
    .A2(_10720_),
    .B1(_10727_),
    .B2(_10735_),
    .Y(_10736_));
 sky130_fd_sc_hd__a22o_2 _25106_ (.A1(net525),
    .A2(\w[0][8] ),
    .B1(_10573_),
    .B2(_10736_),
    .X(_00030_));
 sky130_fd_sc_hd__mux4_1 _25107_ (.A0(\w[18][9] ),
    .A1(\w[16][9] ),
    .A2(\w[22][9] ),
    .A3(\w[20][9] ),
    .S0(net546),
    .S1(net480),
    .X(_10737_));
 sky130_fd_sc_hd__mux4_1 _25108_ (.A0(\w[26][9] ),
    .A1(\w[24][9] ),
    .A2(\w[30][9] ),
    .A3(\w[28][9] ),
    .S0(net546),
    .S1(net480),
    .X(_10738_));
 sky130_fd_sc_hd__mux4_1 _25109_ (.A0(\w[2][9] ),
    .A1(\w[0][9] ),
    .A2(\w[6][9] ),
    .A3(\w[4][9] ),
    .S0(net546),
    .S1(net480),
    .X(_10739_));
 sky130_fd_sc_hd__mux4_1 _25110_ (.A0(\w[10][9] ),
    .A1(\w[8][9] ),
    .A2(\w[14][9] ),
    .A3(\w[12][9] ),
    .S0(net546),
    .S1(net480),
    .X(_10740_));
 sky130_fd_sc_hd__mux4_1 _25111_ (.A0(_10737_),
    .A1(_10738_),
    .A2(_10739_),
    .A3(_10740_),
    .S0(net504),
    .S1(net496),
    .X(_10741_));
 sky130_fd_sc_hd__mux4_1 _25112_ (.A0(\w[34][9] ),
    .A1(\w[32][9] ),
    .A2(\w[38][9] ),
    .A3(\w[36][9] ),
    .S0(net548),
    .S1(net482),
    .X(_10742_));
 sky130_fd_sc_hd__nand2_1 _25113_ (.A(net460),
    .B(_10742_),
    .Y(_10743_));
 sky130_fd_sc_hd__mux4_1 _25114_ (.A0(\w[42][9] ),
    .A1(\w[40][9] ),
    .A2(\w[46][9] ),
    .A3(\w[44][9] ),
    .S0(net548),
    .S1(net482),
    .X(_10744_));
 sky130_fd_sc_hd__mux4_1 _25115_ (.A0(\w[50][9] ),
    .A1(\w[48][9] ),
    .A2(\w[54][9] ),
    .A3(\w[52][9] ),
    .S0(net548),
    .S1(net482),
    .X(_10745_));
 sky130_fd_sc_hd__nand2_1 _25116_ (.A(net492),
    .B(_10745_),
    .Y(_10746_));
 sky130_fd_sc_hd__mux4_1 _25117_ (.A0(\w[58][9] ),
    .A1(\w[56][9] ),
    .A2(\w[62][9] ),
    .A3(\w[60][9] ),
    .S0(net548),
    .S1(net482),
    .X(_10747_));
 sky130_fd_sc_hd__nand2_1 _25118_ (.A(net504),
    .B(_10747_),
    .Y(_10748_));
 sky130_fd_sc_hd__a21oi_1 _25119_ (.A1(_10746_),
    .A2(_10748_),
    .B1(net499),
    .Y(_10749_));
 sky130_fd_sc_hd__a31oi_1 _25120_ (.A1(net499),
    .A2(net504),
    .A3(_10744_),
    .B1(_10749_),
    .Y(_10750_));
 sky130_fd_sc_hd__a21oi_1 _25121_ (.A1(_10743_),
    .A2(_10750_),
    .B1(_10508_),
    .Y(_10751_));
 sky130_fd_sc_hd__a21oi_1 _25122_ (.A1(_10508_),
    .A2(_10741_),
    .B1(_10751_),
    .Y(_10752_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_414 ();
 sky130_fd_sc_hd__nand2_1 _25124_ (.A(net526),
    .B(\w[0][9] ),
    .Y(_10754_));
 sky130_fd_sc_hd__o21ai_4 _25125_ (.A1(net453),
    .A2(_10752_),
    .B1(_10754_),
    .Y(_00031_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__mux4_1 _25128_ (.A0(\w[50][10] ),
    .A1(\w[48][10] ),
    .A2(\w[54][10] ),
    .A3(\w[52][10] ),
    .S0(net552),
    .S1(net483),
    .X(_10757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__mux4_1 _25130_ (.A0(\w[58][10] ),
    .A1(\w[56][10] ),
    .A2(\w[62][10] ),
    .A3(\w[60][10] ),
    .S0(net551),
    .S1(net479),
    .X(_10759_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__mux4_1 _25132_ (.A0(\w[34][10] ),
    .A1(\w[32][10] ),
    .A2(\w[38][10] ),
    .A3(\w[36][10] ),
    .S0(net552),
    .S1(net483),
    .X(_10761_));
 sky130_fd_sc_hd__mux4_1 _25133_ (.A0(\w[42][10] ),
    .A1(\w[40][10] ),
    .A2(\w[46][10] ),
    .A3(\w[44][10] ),
    .S0(net552),
    .S1(net483),
    .X(_10762_));
 sky130_fd_sc_hd__mux4_1 _25134_ (.A0(_10757_),
    .A1(_10759_),
    .A2(_10761_),
    .A3(_10762_),
    .S0(net502),
    .S1(net495),
    .X(_10763_));
 sky130_fd_sc_hd__mux4_1 _25135_ (.A0(\w[2][10] ),
    .A1(\w[0][10] ),
    .A2(\w[6][10] ),
    .A3(\w[4][10] ),
    .S0(net550),
    .S1(net478),
    .X(_10764_));
 sky130_fd_sc_hd__nand2_1 _25136_ (.A(_10513_),
    .B(_10764_),
    .Y(_10765_));
 sky130_fd_sc_hd__mux4_1 _25137_ (.A0(\w[10][10] ),
    .A1(\w[8][10] ),
    .A2(\w[14][10] ),
    .A3(\w[12][10] ),
    .S0(net550),
    .S1(net478),
    .X(_10766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__mux4_1 _25139_ (.A0(\w[18][10] ),
    .A1(\w[16][10] ),
    .A2(\w[22][10] ),
    .A3(\w[20][10] ),
    .S0(net550),
    .S1(net478),
    .X(_10768_));
 sky130_fd_sc_hd__nand2_1 _25140_ (.A(net490),
    .B(_10768_),
    .Y(_10769_));
 sky130_fd_sc_hd__mux4_1 _25141_ (.A0(\w[26][10] ),
    .A1(\w[24][10] ),
    .A2(\w[30][10] ),
    .A3(\w[28][10] ),
    .S0(net550),
    .S1(net478),
    .X(_10770_));
 sky130_fd_sc_hd__nand2_1 _25142_ (.A(net501),
    .B(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__a21oi_1 _25143_ (.A1(_10769_),
    .A2(_10771_),
    .B1(net493),
    .Y(_10772_));
 sky130_fd_sc_hd__a31oi_1 _25144_ (.A1(net493),
    .A2(net501),
    .A3(_10766_),
    .B1(_10772_),
    .Y(_10773_));
 sky130_fd_sc_hd__a21oi_2 _25145_ (.A1(_10765_),
    .A2(_10773_),
    .B1(net458),
    .Y(_10774_));
 sky130_fd_sc_hd__a21oi_1 _25146_ (.A1(net458),
    .A2(_10763_),
    .B1(_10774_),
    .Y(_10775_));
 sky130_fd_sc_hd__nand2_1 _25147_ (.A(net525),
    .B(\w[0][10] ),
    .Y(_10776_));
 sky130_fd_sc_hd__o21ai_1 _25148_ (.A1(net455),
    .A2(_10775_),
    .B1(_10776_),
    .Y(_00001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__mux4_1 _25150_ (.A0(\w[2][11] ),
    .A1(\w[0][11] ),
    .A2(\w[6][11] ),
    .A3(\w[4][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10778_));
 sky130_fd_sc_hd__mux4_1 _25151_ (.A0(\w[34][11] ),
    .A1(\w[32][11] ),
    .A2(\w[38][11] ),
    .A3(\w[36][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10779_));
 sky130_fd_sc_hd__mux2i_1 _25152_ (.A0(_10778_),
    .A1(_10779_),
    .S(net457),
    .Y(_10780_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__mux4_1 _25154_ (.A0(\w[10][11] ),
    .A1(\w[8][11] ),
    .A2(\w[14][11] ),
    .A3(\w[12][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10782_));
 sky130_fd_sc_hd__mux4_1 _25155_ (.A0(\w[18][11] ),
    .A1(\w[16][11] ),
    .A2(\w[22][11] ),
    .A3(\w[20][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10783_));
 sky130_fd_sc_hd__nand2_1 _25156_ (.A(net489),
    .B(_10783_),
    .Y(_10784_));
 sky130_fd_sc_hd__mux4_1 _25157_ (.A0(\w[26][11] ),
    .A1(\w[24][11] ),
    .A2(\w[30][11] ),
    .A3(\w[28][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10785_));
 sky130_fd_sc_hd__nand2_1 _25158_ (.A(net502),
    .B(_10785_),
    .Y(_10786_));
 sky130_fd_sc_hd__a21oi_1 _25159_ (.A1(_10784_),
    .A2(_10786_),
    .B1(net495),
    .Y(_10787_));
 sky130_fd_sc_hd__a311oi_1 _25160_ (.A1(net495),
    .A2(net502),
    .A3(_10782_),
    .B1(_10787_),
    .C1(net457),
    .Y(_10788_));
 sky130_fd_sc_hd__mux4_1 _25161_ (.A0(\w[42][11] ),
    .A1(\w[40][11] ),
    .A2(\w[46][11] ),
    .A3(\w[44][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10789_));
 sky130_fd_sc_hd__mux4_1 _25162_ (.A0(\w[50][11] ),
    .A1(\w[48][11] ),
    .A2(\w[54][11] ),
    .A3(\w[52][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10790_));
 sky130_fd_sc_hd__nand2_1 _25163_ (.A(net491),
    .B(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__mux4_1 _25164_ (.A0(\w[58][11] ),
    .A1(\w[56][11] ),
    .A2(\w[62][11] ),
    .A3(\w[60][11] ),
    .S0(net551),
    .S1(net479),
    .X(_10792_));
 sky130_fd_sc_hd__nand2_1 _25165_ (.A(net500),
    .B(_10792_),
    .Y(_10793_));
 sky130_fd_sc_hd__a21oi_1 _25166_ (.A1(_10791_),
    .A2(_10793_),
    .B1(net495),
    .Y(_10794_));
 sky130_fd_sc_hd__a311oi_2 _25167_ (.A1(net495),
    .A2(net500),
    .A3(_10789_),
    .B1(_10794_),
    .C1(net462),
    .Y(_10795_));
 sky130_fd_sc_hd__o22ai_1 _25168_ (.A1(_10575_),
    .A2(_10780_),
    .B1(_10788_),
    .B2(_10795_),
    .Y(_10796_));
 sky130_fd_sc_hd__a22o_2 _25169_ (.A1(net526),
    .A2(\w[0][11] ),
    .B1(_10573_),
    .B2(_10796_),
    .X(_00002_));
 sky130_fd_sc_hd__mux4_1 _25170_ (.A0(\w[50][12] ),
    .A1(\w[48][12] ),
    .A2(\w[54][12] ),
    .A3(\w[52][12] ),
    .S0(net547),
    .S1(net481),
    .X(_10797_));
 sky130_fd_sc_hd__mux4_1 _25171_ (.A0(\w[58][12] ),
    .A1(\w[56][12] ),
    .A2(\w[62][12] ),
    .A3(\w[60][12] ),
    .S0(net548),
    .S1(net482),
    .X(_10798_));
 sky130_fd_sc_hd__mux4_1 _25172_ (.A0(\w[34][12] ),
    .A1(\w[32][12] ),
    .A2(\w[38][12] ),
    .A3(\w[36][12] ),
    .S0(net547),
    .S1(net481),
    .X(_10799_));
 sky130_fd_sc_hd__mux4_1 _25173_ (.A0(\w[42][12] ),
    .A1(\w[40][12] ),
    .A2(\w[46][12] ),
    .A3(\w[44][12] ),
    .S0(net547),
    .S1(net481),
    .X(_10800_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__mux4_2 _25175_ (.A0(_10797_),
    .A1(_10798_),
    .A2(_10799_),
    .A3(_10800_),
    .S0(net506),
    .S1(net499),
    .X(_10802_));
 sky130_fd_sc_hd__mux4_1 _25176_ (.A0(\w[2][12] ),
    .A1(\w[0][12] ),
    .A2(\w[6][12] ),
    .A3(\w[4][12] ),
    .S0(net547),
    .S1(net481),
    .X(_10803_));
 sky130_fd_sc_hd__nand2_1 _25177_ (.A(net460),
    .B(_10803_),
    .Y(_10804_));
 sky130_fd_sc_hd__mux4_1 _25178_ (.A0(\w[10][12] ),
    .A1(\w[8][12] ),
    .A2(\w[14][12] ),
    .A3(\w[12][12] ),
    .S0(net547),
    .S1(net481),
    .X(_10805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__mux4_1 _25180_ (.A0(\w[18][12] ),
    .A1(\w[16][12] ),
    .A2(\w[22][12] ),
    .A3(\w[20][12] ),
    .S0(net547),
    .S1(net481),
    .X(_10807_));
 sky130_fd_sc_hd__nand2_1 _25181_ (.A(net491),
    .B(_10807_),
    .Y(_10808_));
 sky130_fd_sc_hd__mux4_1 _25182_ (.A0(\w[26][12] ),
    .A1(\w[24][12] ),
    .A2(\w[30][12] ),
    .A3(\w[28][12] ),
    .S0(net547),
    .S1(net481),
    .X(_10809_));
 sky130_fd_sc_hd__nand2_1 _25183_ (.A(net505),
    .B(_10809_),
    .Y(_10810_));
 sky130_fd_sc_hd__a21oi_1 _25184_ (.A1(_10808_),
    .A2(_10810_),
    .B1(net498),
    .Y(_10811_));
 sky130_fd_sc_hd__a31oi_1 _25185_ (.A1(net498),
    .A2(net505),
    .A3(_10805_),
    .B1(_10811_),
    .Y(_10812_));
 sky130_fd_sc_hd__a21oi_1 _25186_ (.A1(_10804_),
    .A2(_10812_),
    .B1(net456),
    .Y(_10813_));
 sky130_fd_sc_hd__a21oi_1 _25187_ (.A1(net456),
    .A2(_10802_),
    .B1(_10813_),
    .Y(_10814_));
 sky130_fd_sc_hd__nand2_1 _25188_ (.A(net526),
    .B(\w[0][12] ),
    .Y(_10815_));
 sky130_fd_sc_hd__o21ai_4 _25189_ (.A1(net455),
    .A2(_10814_),
    .B1(_10815_),
    .Y(_00003_));
 sky130_fd_sc_hd__mux4_1 _25190_ (.A0(\w[2][13] ),
    .A1(\w[0][13] ),
    .A2(\w[6][13] ),
    .A3(\w[4][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10816_));
 sky130_fd_sc_hd__mux4_1 _25191_ (.A0(\w[34][13] ),
    .A1(\w[32][13] ),
    .A2(\w[38][13] ),
    .A3(\w[36][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10817_));
 sky130_fd_sc_hd__mux2i_1 _25192_ (.A0(_10816_),
    .A1(_10817_),
    .S(net457),
    .Y(_10818_));
 sky130_fd_sc_hd__mux4_1 _25193_ (.A0(\w[10][13] ),
    .A1(\w[8][13] ),
    .A2(\w[14][13] ),
    .A3(\w[12][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10819_));
 sky130_fd_sc_hd__mux4_1 _25194_ (.A0(\w[18][13] ),
    .A1(\w[16][13] ),
    .A2(\w[22][13] ),
    .A3(\w[20][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10820_));
 sky130_fd_sc_hd__nand2_1 _25195_ (.A(net489),
    .B(_10820_),
    .Y(_10821_));
 sky130_fd_sc_hd__mux4_1 _25196_ (.A0(\w[26][13] ),
    .A1(\w[24][13] ),
    .A2(\w[30][13] ),
    .A3(\w[28][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10822_));
 sky130_fd_sc_hd__nand2_1 _25197_ (.A(net500),
    .B(_10822_),
    .Y(_10823_));
 sky130_fd_sc_hd__a21oi_1 _25198_ (.A1(_10821_),
    .A2(_10823_),
    .B1(net494),
    .Y(_10824_));
 sky130_fd_sc_hd__a311oi_1 _25199_ (.A1(net494),
    .A2(net500),
    .A3(_10819_),
    .B1(_10824_),
    .C1(net457),
    .Y(_10825_));
 sky130_fd_sc_hd__mux4_1 _25200_ (.A0(\w[42][13] ),
    .A1(\w[40][13] ),
    .A2(\w[46][13] ),
    .A3(\w[44][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10826_));
 sky130_fd_sc_hd__mux4_1 _25201_ (.A0(\w[50][13] ),
    .A1(\w[48][13] ),
    .A2(\w[54][13] ),
    .A3(\w[52][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10827_));
 sky130_fd_sc_hd__nand2_1 _25202_ (.A(net489),
    .B(_10827_),
    .Y(_10828_));
 sky130_fd_sc_hd__mux4_1 _25203_ (.A0(\w[58][13] ),
    .A1(\w[56][13] ),
    .A2(\w[62][13] ),
    .A3(\w[60][13] ),
    .S0(net549),
    .S1(net477),
    .X(_10829_));
 sky130_fd_sc_hd__nand2_1 _25204_ (.A(net503),
    .B(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__a21oi_1 _25205_ (.A1(_10828_),
    .A2(_10830_),
    .B1(net494),
    .Y(_10831_));
 sky130_fd_sc_hd__a311oi_2 _25206_ (.A1(net494),
    .A2(net503),
    .A3(_10826_),
    .B1(_10831_),
    .C1(net461),
    .Y(_10832_));
 sky130_fd_sc_hd__o22ai_1 _25207_ (.A1(_10575_),
    .A2(_10818_),
    .B1(_10825_),
    .B2(_10832_),
    .Y(_10833_));
 sky130_fd_sc_hd__a22o_2 _25208_ (.A1(net526),
    .A2(\w[0][13] ),
    .B1(_10573_),
    .B2(_10833_),
    .X(_00004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_404 ();
 sky130_fd_sc_hd__mux4_1 _25210_ (.A0(\w[50][14] ),
    .A1(\w[48][14] ),
    .A2(\w[54][14] ),
    .A3(\w[52][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10835_));
 sky130_fd_sc_hd__mux4_1 _25211_ (.A0(\w[58][14] ),
    .A1(\w[56][14] ),
    .A2(\w[62][14] ),
    .A3(\w[60][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10836_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_403 ();
 sky130_fd_sc_hd__mux4_1 _25213_ (.A0(\w[34][14] ),
    .A1(\w[32][14] ),
    .A2(\w[38][14] ),
    .A3(\w[36][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10838_));
 sky130_fd_sc_hd__mux4_1 _25214_ (.A0(\w[42][14] ),
    .A1(\w[40][14] ),
    .A2(\w[46][14] ),
    .A3(\w[44][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10839_));
 sky130_fd_sc_hd__mux4_1 _25215_ (.A0(_10835_),
    .A1(_10836_),
    .A2(_10838_),
    .A3(_10839_),
    .S0(net504),
    .S1(net496),
    .X(_10840_));
 sky130_fd_sc_hd__mux4_1 _25216_ (.A0(\w[2][14] ),
    .A1(\w[0][14] ),
    .A2(\w[6][14] ),
    .A3(\w[4][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10841_));
 sky130_fd_sc_hd__nand2_1 _25217_ (.A(net460),
    .B(_10841_),
    .Y(_10842_));
 sky130_fd_sc_hd__mux4_1 _25218_ (.A0(\w[10][14] ),
    .A1(\w[8][14] ),
    .A2(\w[14][14] ),
    .A3(\w[12][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_402 ();
 sky130_fd_sc_hd__mux4_1 _25220_ (.A0(\w[18][14] ),
    .A1(\w[16][14] ),
    .A2(\w[22][14] ),
    .A3(\w[20][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10845_));
 sky130_fd_sc_hd__nand2_1 _25221_ (.A(net492),
    .B(_10845_),
    .Y(_10846_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__mux4_1 _25223_ (.A0(\w[26][14] ),
    .A1(\w[24][14] ),
    .A2(\w[30][14] ),
    .A3(\w[28][14] ),
    .S0(net548),
    .S1(net482),
    .X(_10848_));
 sky130_fd_sc_hd__nand2_1 _25224_ (.A(net504),
    .B(_10848_),
    .Y(_10849_));
 sky130_fd_sc_hd__a21oi_1 _25225_ (.A1(_10846_),
    .A2(_10849_),
    .B1(net496),
    .Y(_10850_));
 sky130_fd_sc_hd__a31oi_1 _25226_ (.A1(net496),
    .A2(net504),
    .A3(_10843_),
    .B1(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__a21oi_1 _25227_ (.A1(_10842_),
    .A2(_10851_),
    .B1(_10564_),
    .Y(_10852_));
 sky130_fd_sc_hd__a21oi_2 _25228_ (.A1(_10564_),
    .A2(_10840_),
    .B1(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__nand2_1 _25229_ (.A(net526),
    .B(\w[0][14] ),
    .Y(_10854_));
 sky130_fd_sc_hd__o21ai_4 _25230_ (.A1(net453),
    .A2(_10853_),
    .B1(_10854_),
    .Y(_00005_));
 sky130_fd_sc_hd__mux4_1 _25231_ (.A0(\w[50][15] ),
    .A1(\w[48][15] ),
    .A2(\w[54][15] ),
    .A3(\w[52][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10855_));
 sky130_fd_sc_hd__mux4_1 _25232_ (.A0(\w[58][15] ),
    .A1(\w[56][15] ),
    .A2(\w[62][15] ),
    .A3(\w[60][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10856_));
 sky130_fd_sc_hd__mux4_1 _25233_ (.A0(\w[34][15] ),
    .A1(\w[32][15] ),
    .A2(\w[38][15] ),
    .A3(\w[36][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10857_));
 sky130_fd_sc_hd__mux4_1 _25234_ (.A0(\w[42][15] ),
    .A1(\w[40][15] ),
    .A2(\w[46][15] ),
    .A3(\w[44][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10858_));
 sky130_fd_sc_hd__mux4_1 _25235_ (.A0(_10855_),
    .A1(_10856_),
    .A2(_10857_),
    .A3(_10858_),
    .S0(net505),
    .S1(net496),
    .X(_10859_));
 sky130_fd_sc_hd__mux4_1 _25236_ (.A0(\w[2][15] ),
    .A1(\w[0][15] ),
    .A2(\w[6][15] ),
    .A3(\w[4][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10860_));
 sky130_fd_sc_hd__nand2_1 _25237_ (.A(net460),
    .B(_10860_),
    .Y(_10861_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__mux4_1 _25239_ (.A0(\w[10][15] ),
    .A1(\w[8][15] ),
    .A2(\w[14][15] ),
    .A3(\w[12][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10863_));
 sky130_fd_sc_hd__mux4_1 _25240_ (.A0(\w[18][15] ),
    .A1(\w[16][15] ),
    .A2(\w[22][15] ),
    .A3(\w[20][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10864_));
 sky130_fd_sc_hd__nand2_1 _25241_ (.A(net491),
    .B(_10864_),
    .Y(_10865_));
 sky130_fd_sc_hd__mux4_1 _25242_ (.A0(\w[26][15] ),
    .A1(\w[24][15] ),
    .A2(\w[30][15] ),
    .A3(\w[28][15] ),
    .S0(net546),
    .S1(net480),
    .X(_10866_));
 sky130_fd_sc_hd__nand2_1 _25243_ (.A(net505),
    .B(_10866_),
    .Y(_10867_));
 sky130_fd_sc_hd__a21oi_1 _25244_ (.A1(_10865_),
    .A2(_10867_),
    .B1(net496),
    .Y(_10868_));
 sky130_fd_sc_hd__a31oi_1 _25245_ (.A1(net496),
    .A2(net505),
    .A3(_10863_),
    .B1(_10868_),
    .Y(_10869_));
 sky130_fd_sc_hd__a21oi_1 _25246_ (.A1(_10861_),
    .A2(_10869_),
    .B1(net456),
    .Y(_10870_));
 sky130_fd_sc_hd__a21oi_1 _25247_ (.A1(net456),
    .A2(_10859_),
    .B1(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__nand2_1 _25248_ (.A(net526),
    .B(\w[0][15] ),
    .Y(_10872_));
 sky130_fd_sc_hd__o21ai_4 _25249_ (.A1(net455),
    .A2(_10871_),
    .B1(_10872_),
    .Y(_00006_));
 sky130_fd_sc_hd__mux4_1 _25250_ (.A0(\w[2][16] ),
    .A1(\w[0][16] ),
    .A2(\w[6][16] ),
    .A3(\w[4][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10873_));
 sky130_fd_sc_hd__mux4_1 _25251_ (.A0(\w[34][16] ),
    .A1(\w[32][16] ),
    .A2(\w[38][16] ),
    .A3(\w[36][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10874_));
 sky130_fd_sc_hd__mux2i_1 _25252_ (.A0(_10873_),
    .A1(_10874_),
    .S(net457),
    .Y(_10875_));
 sky130_fd_sc_hd__mux4_1 _25253_ (.A0(\w[10][16] ),
    .A1(\w[8][16] ),
    .A2(\w[14][16] ),
    .A3(\w[12][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10876_));
 sky130_fd_sc_hd__mux4_1 _25254_ (.A0(\w[18][16] ),
    .A1(\w[16][16] ),
    .A2(\w[22][16] ),
    .A3(\w[20][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10877_));
 sky130_fd_sc_hd__nand2_1 _25255_ (.A(net491),
    .B(_10877_),
    .Y(_10878_));
 sky130_fd_sc_hd__mux4_1 _25256_ (.A0(\w[26][16] ),
    .A1(\w[24][16] ),
    .A2(\w[30][16] ),
    .A3(\w[28][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10879_));
 sky130_fd_sc_hd__nand2_1 _25257_ (.A(net502),
    .B(_10879_),
    .Y(_10880_));
 sky130_fd_sc_hd__a21oi_1 _25258_ (.A1(_10878_),
    .A2(_10880_),
    .B1(net497),
    .Y(_10881_));
 sky130_fd_sc_hd__a311oi_1 _25259_ (.A1(net497),
    .A2(net502),
    .A3(_10876_),
    .B1(_10881_),
    .C1(net457),
    .Y(_10882_));
 sky130_fd_sc_hd__mux4_1 _25260_ (.A0(\w[42][16] ),
    .A1(\w[40][16] ),
    .A2(\w[46][16] ),
    .A3(\w[44][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10883_));
 sky130_fd_sc_hd__mux4_1 _25261_ (.A0(\w[50][16] ),
    .A1(\w[48][16] ),
    .A2(\w[54][16] ),
    .A3(\w[52][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10884_));
 sky130_fd_sc_hd__nand2_1 _25262_ (.A(net491),
    .B(_10884_),
    .Y(_10885_));
 sky130_fd_sc_hd__mux4_1 _25263_ (.A0(\w[58][16] ),
    .A1(\w[56][16] ),
    .A2(\w[62][16] ),
    .A3(\w[60][16] ),
    .S0(net551),
    .S1(net479),
    .X(_10886_));
 sky130_fd_sc_hd__nand2_1 _25264_ (.A(net502),
    .B(_10886_),
    .Y(_10887_));
 sky130_fd_sc_hd__a21oi_1 _25265_ (.A1(_10885_),
    .A2(_10887_),
    .B1(net497),
    .Y(_10888_));
 sky130_fd_sc_hd__a311oi_2 _25266_ (.A1(net497),
    .A2(net500),
    .A3(_10883_),
    .B1(_10888_),
    .C1(net462),
    .Y(_10889_));
 sky130_fd_sc_hd__o22ai_1 _25267_ (.A1(_10575_),
    .A2(_10875_),
    .B1(_10882_),
    .B2(_10889_),
    .Y(_10890_));
 sky130_fd_sc_hd__a22o_2 _25268_ (.A1(net526),
    .A2(\w[0][16] ),
    .B1(_10573_),
    .B2(_10890_),
    .X(_00007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__mux4_1 _25270_ (.A0(\w[18][17] ),
    .A1(\w[16][17] ),
    .A2(\w[22][17] ),
    .A3(\w[20][17] ),
    .S0(net549),
    .S1(net477),
    .X(_10892_));
 sky130_fd_sc_hd__mux4_1 _25271_ (.A0(\w[26][17] ),
    .A1(\w[24][17] ),
    .A2(\w[30][17] ),
    .A3(\w[28][17] ),
    .S0(net549),
    .S1(net477),
    .X(_10893_));
 sky130_fd_sc_hd__mux4_1 _25272_ (.A0(\w[2][17] ),
    .A1(\w[0][17] ),
    .A2(\w[6][17] ),
    .A3(\w[4][17] ),
    .S0(net549),
    .S1(net477),
    .X(_10894_));
 sky130_fd_sc_hd__mux4_1 _25273_ (.A0(\w[10][17] ),
    .A1(\w[8][17] ),
    .A2(\w[14][17] ),
    .A3(\w[12][17] ),
    .S0(net549),
    .S1(net477),
    .X(_10895_));
 sky130_fd_sc_hd__mux4_4 _25274_ (.A0(_10892_),
    .A1(_10893_),
    .A2(_10894_),
    .A3(_10895_),
    .S0(net501),
    .S1(net493),
    .X(_10896_));
 sky130_fd_sc_hd__mux4_1 _25275_ (.A0(\w[34][17] ),
    .A1(\w[32][17] ),
    .A2(\w[38][17] ),
    .A3(\w[36][17] ),
    .S0(net552),
    .S1(net483),
    .X(_10897_));
 sky130_fd_sc_hd__nand2_1 _25276_ (.A(net460),
    .B(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__mux4_1 _25277_ (.A0(\w[42][17] ),
    .A1(\w[40][17] ),
    .A2(\w[46][17] ),
    .A3(\w[44][17] ),
    .S0(net552),
    .S1(net483),
    .X(_10899_));
 sky130_fd_sc_hd__mux4_1 _25278_ (.A0(\w[50][17] ),
    .A1(\w[48][17] ),
    .A2(\w[54][17] ),
    .A3(\w[52][17] ),
    .S0(net552),
    .S1(net483),
    .X(_10900_));
 sky130_fd_sc_hd__nand2_1 _25279_ (.A(net489),
    .B(_10900_),
    .Y(_10901_));
 sky130_fd_sc_hd__mux4_1 _25280_ (.A0(\w[58][17] ),
    .A1(\w[56][17] ),
    .A2(\w[62][17] ),
    .A3(\w[60][17] ),
    .S0(net552),
    .S1(net483),
    .X(_10902_));
 sky130_fd_sc_hd__nand2_1 _25281_ (.A(net500),
    .B(_10902_),
    .Y(_10903_));
 sky130_fd_sc_hd__a21oi_1 _25282_ (.A1(_10901_),
    .A2(_10903_),
    .B1(net495),
    .Y(_10904_));
 sky130_fd_sc_hd__a31oi_1 _25283_ (.A1(net495),
    .A2(net500),
    .A3(_10899_),
    .B1(_10904_),
    .Y(_10905_));
 sky130_fd_sc_hd__a21oi_1 _25284_ (.A1(_10898_),
    .A2(_10905_),
    .B1(net462),
    .Y(_10906_));
 sky130_fd_sc_hd__a21oi_1 _25285_ (.A1(net462),
    .A2(_10896_),
    .B1(_10906_),
    .Y(_10907_));
 sky130_fd_sc_hd__nand2_2 _25286_ (.A(net525),
    .B(\w[0][17] ),
    .Y(_10908_));
 sky130_fd_sc_hd__o21ai_4 _25287_ (.A1(net455),
    .A2(_10907_),
    .B1(_10908_),
    .Y(_00008_));
 sky130_fd_sc_hd__mux4_1 _25288_ (.A0(\w[18][18] ),
    .A1(\w[16][18] ),
    .A2(\w[22][18] ),
    .A3(\w[20][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10909_));
 sky130_fd_sc_hd__mux4_1 _25289_ (.A0(\w[26][18] ),
    .A1(\w[24][18] ),
    .A2(\w[30][18] ),
    .A3(\w[28][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10910_));
 sky130_fd_sc_hd__mux4_1 _25290_ (.A0(\w[2][18] ),
    .A1(\w[0][18] ),
    .A2(\w[6][18] ),
    .A3(\w[4][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10911_));
 sky130_fd_sc_hd__mux4_1 _25291_ (.A0(\w[10][18] ),
    .A1(\w[8][18] ),
    .A2(\w[14][18] ),
    .A3(\w[12][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10912_));
 sky130_fd_sc_hd__mux4_1 _25292_ (.A0(_10909_),
    .A1(_10910_),
    .A2(_10911_),
    .A3(_10912_),
    .S0(net504),
    .S1(net496),
    .X(_10913_));
 sky130_fd_sc_hd__mux4_1 _25293_ (.A0(\w[50][18] ),
    .A1(\w[48][18] ),
    .A2(\w[54][18] ),
    .A3(\w[52][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10914_));
 sky130_fd_sc_hd__mux4_1 _25294_ (.A0(\w[58][18] ),
    .A1(\w[56][18] ),
    .A2(\w[62][18] ),
    .A3(\w[60][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10915_));
 sky130_fd_sc_hd__mux4_1 _25295_ (.A0(\w[34][18] ),
    .A1(\w[32][18] ),
    .A2(\w[38][18] ),
    .A3(\w[36][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10916_));
 sky130_fd_sc_hd__mux4_1 _25296_ (.A0(\w[42][18] ),
    .A1(\w[40][18] ),
    .A2(\w[46][18] ),
    .A3(\w[44][18] ),
    .S0(net548),
    .S1(net482),
    .X(_10917_));
 sky130_fd_sc_hd__mux4_1 _25297_ (.A0(_10914_),
    .A1(_10915_),
    .A2(_10916_),
    .A3(_10917_),
    .S0(net504),
    .S1(net496),
    .X(_10918_));
 sky130_fd_sc_hd__mux2i_2 _25298_ (.A0(_10913_),
    .A1(_10918_),
    .S(_10564_),
    .Y(_10919_));
 sky130_fd_sc_hd__nand2_1 _25299_ (.A(net526),
    .B(\w[0][18] ),
    .Y(_10920_));
 sky130_fd_sc_hd__o21ai_4 _25300_ (.A1(net453),
    .A2(_10919_),
    .B1(_10920_),
    .Y(_00009_));
 sky130_fd_sc_hd__mux4_1 _25301_ (.A0(\w[50][19] ),
    .A1(\w[48][19] ),
    .A2(\w[54][19] ),
    .A3(\w[52][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10921_));
 sky130_fd_sc_hd__mux4_1 _25302_ (.A0(\w[58][19] ),
    .A1(\w[56][19] ),
    .A2(\w[62][19] ),
    .A3(\w[60][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10922_));
 sky130_fd_sc_hd__mux4_1 _25303_ (.A0(\w[34][19] ),
    .A1(\w[32][19] ),
    .A2(\w[38][19] ),
    .A3(\w[36][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10923_));
 sky130_fd_sc_hd__mux4_1 _25304_ (.A0(\w[42][19] ),
    .A1(\w[40][19] ),
    .A2(\w[46][19] ),
    .A3(\w[44][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10924_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__mux4_1 _25306_ (.A0(_10921_),
    .A1(_10922_),
    .A2(_10923_),
    .A3(_10924_),
    .S0(net504),
    .S1(net496),
    .X(_10926_));
 sky130_fd_sc_hd__mux4_1 _25307_ (.A0(\w[2][19] ),
    .A1(\w[0][19] ),
    .A2(\w[6][19] ),
    .A3(\w[4][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10927_));
 sky130_fd_sc_hd__nand2_1 _25308_ (.A(net460),
    .B(_10927_),
    .Y(_10928_));
 sky130_fd_sc_hd__mux4_1 _25309_ (.A0(\w[10][19] ),
    .A1(\w[8][19] ),
    .A2(\w[14][19] ),
    .A3(\w[12][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10929_));
 sky130_fd_sc_hd__mux4_1 _25310_ (.A0(\w[18][19] ),
    .A1(\w[16][19] ),
    .A2(\w[22][19] ),
    .A3(\w[20][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10930_));
 sky130_fd_sc_hd__nand2_1 _25311_ (.A(net491),
    .B(_10930_),
    .Y(_10931_));
 sky130_fd_sc_hd__mux4_1 _25312_ (.A0(\w[26][19] ),
    .A1(\w[24][19] ),
    .A2(\w[30][19] ),
    .A3(\w[28][19] ),
    .S0(net546),
    .S1(net480),
    .X(_10932_));
 sky130_fd_sc_hd__nand2_1 _25313_ (.A(net504),
    .B(_10932_),
    .Y(_10933_));
 sky130_fd_sc_hd__a21oi_1 _25314_ (.A1(_10931_),
    .A2(_10933_),
    .B1(net496),
    .Y(_10934_));
 sky130_fd_sc_hd__a31oi_1 _25315_ (.A1(net496),
    .A2(net504),
    .A3(_10929_),
    .B1(_10934_),
    .Y(_10935_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__a21oi_1 _25317_ (.A1(_10928_),
    .A2(_10935_),
    .B1(net456),
    .Y(_10937_));
 sky130_fd_sc_hd__a21oi_1 _25318_ (.A1(net456),
    .A2(_10926_),
    .B1(_10937_),
    .Y(_10938_));
 sky130_fd_sc_hd__nand2_1 _25319_ (.A(net526),
    .B(\w[0][19] ),
    .Y(_10939_));
 sky130_fd_sc_hd__o21ai_4 _25320_ (.A1(net455),
    .A2(_10938_),
    .B1(_10939_),
    .Y(_00010_));
 sky130_fd_sc_hd__mux4_1 _25321_ (.A0(\w[2][20] ),
    .A1(\w[0][20] ),
    .A2(\w[6][20] ),
    .A3(\w[4][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10940_));
 sky130_fd_sc_hd__mux4_1 _25322_ (.A0(\w[34][20] ),
    .A1(\w[32][20] ),
    .A2(\w[38][20] ),
    .A3(\w[36][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10941_));
 sky130_fd_sc_hd__mux2i_1 _25323_ (.A0(_10940_),
    .A1(_10941_),
    .S(net458),
    .Y(_10942_));
 sky130_fd_sc_hd__mux4_2 _25324_ (.A0(\w[10][20] ),
    .A1(\w[8][20] ),
    .A2(\w[14][20] ),
    .A3(\w[12][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10943_));
 sky130_fd_sc_hd__mux4_1 _25325_ (.A0(\w[18][20] ),
    .A1(\w[16][20] ),
    .A2(\w[22][20] ),
    .A3(\w[20][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10944_));
 sky130_fd_sc_hd__nand2_1 _25326_ (.A(net490),
    .B(_10944_),
    .Y(_10945_));
 sky130_fd_sc_hd__mux4_1 _25327_ (.A0(\w[26][20] ),
    .A1(\w[24][20] ),
    .A2(\w[30][20] ),
    .A3(\w[28][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10946_));
 sky130_fd_sc_hd__nand2_1 _25328_ (.A(net501),
    .B(_10946_),
    .Y(_10947_));
 sky130_fd_sc_hd__a21oi_1 _25329_ (.A1(_10945_),
    .A2(_10947_),
    .B1(net493),
    .Y(_10948_));
 sky130_fd_sc_hd__a311oi_2 _25330_ (.A1(net493),
    .A2(net501),
    .A3(_10943_),
    .B1(_10948_),
    .C1(net458),
    .Y(_10949_));
 sky130_fd_sc_hd__mux4_1 _25331_ (.A0(\w[42][20] ),
    .A1(\w[40][20] ),
    .A2(\w[46][20] ),
    .A3(\w[44][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10950_));
 sky130_fd_sc_hd__mux4_1 _25332_ (.A0(\w[50][20] ),
    .A1(\w[48][20] ),
    .A2(\w[54][20] ),
    .A3(\w[52][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10951_));
 sky130_fd_sc_hd__nand2_1 _25333_ (.A(net489),
    .B(_10951_),
    .Y(_10952_));
 sky130_fd_sc_hd__mux4_1 _25334_ (.A0(\w[58][20] ),
    .A1(\w[56][20] ),
    .A2(\w[62][20] ),
    .A3(\w[60][20] ),
    .S0(net549),
    .S1(net477),
    .X(_10953_));
 sky130_fd_sc_hd__nand2_1 _25335_ (.A(net503),
    .B(_10953_),
    .Y(_10954_));
 sky130_fd_sc_hd__a21oi_1 _25336_ (.A1(_10952_),
    .A2(_10954_),
    .B1(net494),
    .Y(_10955_));
 sky130_fd_sc_hd__a311oi_1 _25337_ (.A1(net494),
    .A2(net503),
    .A3(_10950_),
    .B1(_10955_),
    .C1(net461),
    .Y(_10956_));
 sky130_fd_sc_hd__o22ai_1 _25338_ (.A1(_10575_),
    .A2(_10942_),
    .B1(_10949_),
    .B2(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__a22o_2 _25339_ (.A1(net525),
    .A2(\w[0][20] ),
    .B1(_10573_),
    .B2(_10957_),
    .X(_00012_));
 sky130_fd_sc_hd__mux4_1 _25340_ (.A0(\w[50][21] ),
    .A1(\w[48][21] ),
    .A2(\w[54][21] ),
    .A3(\w[52][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10958_));
 sky130_fd_sc_hd__mux4_1 _25341_ (.A0(\w[58][21] ),
    .A1(\w[56][21] ),
    .A2(\w[62][21] ),
    .A3(\w[60][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10959_));
 sky130_fd_sc_hd__mux4_1 _25342_ (.A0(\w[34][21] ),
    .A1(\w[32][21] ),
    .A2(\w[38][21] ),
    .A3(\w[36][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10960_));
 sky130_fd_sc_hd__mux4_1 _25343_ (.A0(\w[42][21] ),
    .A1(\w[40][21] ),
    .A2(\w[46][21] ),
    .A3(\w[44][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10961_));
 sky130_fd_sc_hd__mux4_2 _25344_ (.A0(_10958_),
    .A1(_10959_),
    .A2(_10960_),
    .A3(_10961_),
    .S0(net506),
    .S1(net498),
    .X(_10962_));
 sky130_fd_sc_hd__mux4_1 _25345_ (.A0(\w[2][21] ),
    .A1(\w[0][21] ),
    .A2(\w[6][21] ),
    .A3(\w[4][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10963_));
 sky130_fd_sc_hd__nand2_1 _25346_ (.A(net460),
    .B(_10963_),
    .Y(_10964_));
 sky130_fd_sc_hd__mux4_1 _25347_ (.A0(\w[10][21] ),
    .A1(\w[8][21] ),
    .A2(\w[14][21] ),
    .A3(\w[12][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10965_));
 sky130_fd_sc_hd__mux4_1 _25348_ (.A0(\w[18][21] ),
    .A1(\w[16][21] ),
    .A2(\w[22][21] ),
    .A3(\w[20][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10966_));
 sky130_fd_sc_hd__nand2_1 _25349_ (.A(net491),
    .B(_10966_),
    .Y(_10967_));
 sky130_fd_sc_hd__mux4_1 _25350_ (.A0(\w[26][21] ),
    .A1(\w[24][21] ),
    .A2(\w[30][21] ),
    .A3(\w[28][21] ),
    .S0(net547),
    .S1(net481),
    .X(_10968_));
 sky130_fd_sc_hd__nand2_1 _25351_ (.A(net505),
    .B(_10968_),
    .Y(_10969_));
 sky130_fd_sc_hd__a21oi_1 _25352_ (.A1(_10967_),
    .A2(_10969_),
    .B1(net497),
    .Y(_10970_));
 sky130_fd_sc_hd__a31oi_1 _25353_ (.A1(net497),
    .A2(net505),
    .A3(_10965_),
    .B1(_10970_),
    .Y(_10971_));
 sky130_fd_sc_hd__a21oi_1 _25354_ (.A1(_10964_),
    .A2(_10971_),
    .B1(net456),
    .Y(_10972_));
 sky130_fd_sc_hd__a21oi_1 _25355_ (.A1(net456),
    .A2(_10962_),
    .B1(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__nand2_1 _25356_ (.A(net526),
    .B(\w[0][21] ),
    .Y(_10974_));
 sky130_fd_sc_hd__o21ai_4 _25357_ (.A1(net455),
    .A2(_10973_),
    .B1(_10974_),
    .Y(_00013_));
 sky130_fd_sc_hd__mux4_1 _25358_ (.A0(\w[18][22] ),
    .A1(\w[16][22] ),
    .A2(\w[22][22] ),
    .A3(\w[20][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10975_));
 sky130_fd_sc_hd__mux4_1 _25359_ (.A0(\w[26][22] ),
    .A1(\w[24][22] ),
    .A2(\w[30][22] ),
    .A3(\w[28][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10976_));
 sky130_fd_sc_hd__mux4_1 _25360_ (.A0(\w[2][22] ),
    .A1(\w[0][22] ),
    .A2(\w[6][22] ),
    .A3(\w[4][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10977_));
 sky130_fd_sc_hd__mux4_1 _25361_ (.A0(\w[10][22] ),
    .A1(\w[8][22] ),
    .A2(\w[14][22] ),
    .A3(\w[12][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10978_));
 sky130_fd_sc_hd__mux4_1 _25362_ (.A0(_10975_),
    .A1(_10976_),
    .A2(_10977_),
    .A3(_10978_),
    .S0(net505),
    .S1(net497),
    .X(_10979_));
 sky130_fd_sc_hd__mux4_1 _25363_ (.A0(\w[34][22] ),
    .A1(\w[32][22] ),
    .A2(\w[38][22] ),
    .A3(\w[36][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10980_));
 sky130_fd_sc_hd__nand2_1 _25364_ (.A(net460),
    .B(_10980_),
    .Y(_10981_));
 sky130_fd_sc_hd__mux4_1 _25365_ (.A0(\w[42][22] ),
    .A1(\w[40][22] ),
    .A2(\w[46][22] ),
    .A3(\w[44][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10982_));
 sky130_fd_sc_hd__mux4_1 _25366_ (.A0(\w[50][22] ),
    .A1(\w[48][22] ),
    .A2(\w[54][22] ),
    .A3(\w[52][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10983_));
 sky130_fd_sc_hd__nand2_1 _25367_ (.A(net491),
    .B(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__mux4_1 _25368_ (.A0(\w[58][22] ),
    .A1(\w[56][22] ),
    .A2(\w[62][22] ),
    .A3(\w[60][22] ),
    .S0(net547),
    .S1(net481),
    .X(_10985_));
 sky130_fd_sc_hd__nand2_1 _25369_ (.A(net505),
    .B(_10985_),
    .Y(_10986_));
 sky130_fd_sc_hd__a21oi_1 _25370_ (.A1(_10984_),
    .A2(_10986_),
    .B1(net498),
    .Y(_10987_));
 sky130_fd_sc_hd__a31oi_1 _25371_ (.A1(net498),
    .A2(net505),
    .A3(_10982_),
    .B1(_10987_),
    .Y(_10988_));
 sky130_fd_sc_hd__a21oi_1 _25372_ (.A1(_10981_),
    .A2(_10988_),
    .B1(net462),
    .Y(_10989_));
 sky130_fd_sc_hd__a21oi_1 _25373_ (.A1(net462),
    .A2(_10979_),
    .B1(_10989_),
    .Y(_10990_));
 sky130_fd_sc_hd__nand2_1 _25374_ (.A(net526),
    .B(\w[0][22] ),
    .Y(_10991_));
 sky130_fd_sc_hd__o21ai_4 _25375_ (.A1(net455),
    .A2(_10990_),
    .B1(_10991_),
    .Y(_00014_));
 sky130_fd_sc_hd__mux4_1 _25376_ (.A0(\w[18][23] ),
    .A1(\w[16][23] ),
    .A2(\w[22][23] ),
    .A3(\w[20][23] ),
    .S0(net548),
    .S1(net482),
    .X(_10992_));
 sky130_fd_sc_hd__mux4_1 _25377_ (.A0(\w[26][23] ),
    .A1(\w[24][23] ),
    .A2(\w[30][23] ),
    .A3(\w[28][23] ),
    .S0(net548),
    .S1(net482),
    .X(_10993_));
 sky130_fd_sc_hd__mux4_1 _25378_ (.A0(\w[2][23] ),
    .A1(\w[0][23] ),
    .A2(\w[6][23] ),
    .A3(\w[4][23] ),
    .S0(net548),
    .S1(net482),
    .X(_10994_));
 sky130_fd_sc_hd__mux4_1 _25379_ (.A0(\w[10][23] ),
    .A1(\w[8][23] ),
    .A2(\w[14][23] ),
    .A3(\w[12][23] ),
    .S0(net548),
    .S1(net482),
    .X(_10995_));
 sky130_fd_sc_hd__mux4_2 _25380_ (.A0(_10992_),
    .A1(_10993_),
    .A2(_10994_),
    .A3(_10995_),
    .S0(net504),
    .S1(net496),
    .X(_10996_));
 sky130_fd_sc_hd__mux4_1 _25381_ (.A0(\w[34][23] ),
    .A1(\w[32][23] ),
    .A2(\w[38][23] ),
    .A3(\w[36][23] ),
    .S0(net548),
    .S1(net482),
    .X(_10997_));
 sky130_fd_sc_hd__nand2_1 _25382_ (.A(net460),
    .B(_10997_),
    .Y(_10998_));
 sky130_fd_sc_hd__mux4_1 _25383_ (.A0(\w[42][23] ),
    .A1(\w[40][23] ),
    .A2(\w[46][23] ),
    .A3(\w[44][23] ),
    .S0(net548),
    .S1(net482),
    .X(_10999_));
 sky130_fd_sc_hd__mux4_1 _25384_ (.A0(\w[50][23] ),
    .A1(\w[48][23] ),
    .A2(\w[54][23] ),
    .A3(\w[52][23] ),
    .S0(net548),
    .S1(net482),
    .X(_11000_));
 sky130_fd_sc_hd__nand2_1 _25385_ (.A(net492),
    .B(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__mux4_1 _25386_ (.A0(\w[58][23] ),
    .A1(\w[56][23] ),
    .A2(\w[62][23] ),
    .A3(\w[60][23] ),
    .S0(net548),
    .S1(net482),
    .X(_11002_));
 sky130_fd_sc_hd__nand2_1 _25387_ (.A(net504),
    .B(_11002_),
    .Y(_11003_));
 sky130_fd_sc_hd__a21oi_1 _25388_ (.A1(_11001_),
    .A2(_11003_),
    .B1(net499),
    .Y(_11004_));
 sky130_fd_sc_hd__a31oi_1 _25389_ (.A1(net499),
    .A2(net504),
    .A3(_10999_),
    .B1(_11004_),
    .Y(_11005_));
 sky130_fd_sc_hd__a21oi_2 _25390_ (.A1(_10998_),
    .A2(_11005_),
    .B1(_10508_),
    .Y(_11006_));
 sky130_fd_sc_hd__a21oi_1 _25391_ (.A1(_10508_),
    .A2(_10996_),
    .B1(_11006_),
    .Y(_11007_));
 sky130_fd_sc_hd__nand2_1 _25392_ (.A(net526),
    .B(\w[0][23] ),
    .Y(_11008_));
 sky130_fd_sc_hd__o21ai_4 _25393_ (.A1(net453),
    .A2(_11007_),
    .B1(_11008_),
    .Y(_00015_));
 sky130_fd_sc_hd__mux4_2 _25394_ (.A0(\w[2][24] ),
    .A1(\w[0][24] ),
    .A2(\w[6][24] ),
    .A3(\w[4][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11009_));
 sky130_fd_sc_hd__mux4_1 _25395_ (.A0(\w[34][24] ),
    .A1(\w[32][24] ),
    .A2(\w[38][24] ),
    .A3(\w[36][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11010_));
 sky130_fd_sc_hd__mux2i_1 _25396_ (.A0(_11009_),
    .A1(_11010_),
    .S(net458),
    .Y(_11011_));
 sky130_fd_sc_hd__mux4_1 _25397_ (.A0(\w[10][24] ),
    .A1(\w[8][24] ),
    .A2(\w[14][24] ),
    .A3(\w[12][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11012_));
 sky130_fd_sc_hd__mux4_1 _25398_ (.A0(\w[18][24] ),
    .A1(\w[16][24] ),
    .A2(\w[22][24] ),
    .A3(\w[20][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11013_));
 sky130_fd_sc_hd__nand2_1 _25399_ (.A(net490),
    .B(_11013_),
    .Y(_11014_));
 sky130_fd_sc_hd__mux4_1 _25400_ (.A0(\w[26][24] ),
    .A1(\w[24][24] ),
    .A2(\w[30][24] ),
    .A3(\w[28][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11015_));
 sky130_fd_sc_hd__nand2_1 _25401_ (.A(net501),
    .B(_11015_),
    .Y(_11016_));
 sky130_fd_sc_hd__a21oi_1 _25402_ (.A1(_11014_),
    .A2(_11016_),
    .B1(net493),
    .Y(_11017_));
 sky130_fd_sc_hd__a311oi_1 _25403_ (.A1(net493),
    .A2(net501),
    .A3(_11012_),
    .B1(_11017_),
    .C1(net458),
    .Y(_11018_));
 sky130_fd_sc_hd__mux4_1 _25404_ (.A0(\w[42][24] ),
    .A1(\w[40][24] ),
    .A2(\w[46][24] ),
    .A3(\w[44][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11019_));
 sky130_fd_sc_hd__mux4_1 _25405_ (.A0(\w[50][24] ),
    .A1(\w[48][24] ),
    .A2(\w[54][24] ),
    .A3(\w[52][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11020_));
 sky130_fd_sc_hd__nand2_1 _25406_ (.A(net490),
    .B(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__mux4_1 _25407_ (.A0(\w[58][24] ),
    .A1(\w[56][24] ),
    .A2(\w[62][24] ),
    .A3(\w[60][24] ),
    .S0(net550),
    .S1(net478),
    .X(_11022_));
 sky130_fd_sc_hd__nand2_1 _25408_ (.A(net501),
    .B(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__a21oi_1 _25409_ (.A1(_11021_),
    .A2(_11023_),
    .B1(net493),
    .Y(_11024_));
 sky130_fd_sc_hd__a311oi_2 _25410_ (.A1(net493),
    .A2(net501),
    .A3(_11019_),
    .B1(_11024_),
    .C1(net461),
    .Y(_11025_));
 sky130_fd_sc_hd__o22ai_1 _25411_ (.A1(_10575_),
    .A2(_11011_),
    .B1(_11018_),
    .B2(_11025_),
    .Y(_11026_));
 sky130_fd_sc_hd__a22o_1 _25412_ (.A1(net525),
    .A2(\w[0][24] ),
    .B1(_10573_),
    .B2(_11026_),
    .X(_00016_));
 sky130_fd_sc_hd__mux4_1 _25413_ (.A0(\w[50][25] ),
    .A1(\w[48][25] ),
    .A2(\w[54][25] ),
    .A3(\w[52][25] ),
    .S0(net552),
    .S1(net483),
    .X(_11027_));
 sky130_fd_sc_hd__mux4_1 _25414_ (.A0(\w[58][25] ),
    .A1(\w[56][25] ),
    .A2(\w[62][25] ),
    .A3(\w[60][25] ),
    .S0(net552),
    .S1(net483),
    .X(_11028_));
 sky130_fd_sc_hd__mux4_1 _25415_ (.A0(\w[34][25] ),
    .A1(\w[32][25] ),
    .A2(\w[38][25] ),
    .A3(\w[36][25] ),
    .S0(net552),
    .S1(net483),
    .X(_11029_));
 sky130_fd_sc_hd__mux4_1 _25416_ (.A0(\w[42][25] ),
    .A1(\w[40][25] ),
    .A2(\w[46][25] ),
    .A3(\w[44][25] ),
    .S0(net552),
    .S1(net483),
    .X(_11030_));
 sky130_fd_sc_hd__mux4_4 _25417_ (.A0(_11027_),
    .A1(_11028_),
    .A2(_11029_),
    .A3(_11030_),
    .S0(net502),
    .S1(net495),
    .X(_11031_));
 sky130_fd_sc_hd__mux4_1 _25418_ (.A0(\w[2][25] ),
    .A1(\w[0][25] ),
    .A2(\w[6][25] ),
    .A3(\w[4][25] ),
    .S0(net551),
    .S1(net479),
    .X(_11032_));
 sky130_fd_sc_hd__nand2_1 _25419_ (.A(net460),
    .B(_11032_),
    .Y(_11033_));
 sky130_fd_sc_hd__mux4_1 _25420_ (.A0(\w[10][25] ),
    .A1(\w[8][25] ),
    .A2(\w[14][25] ),
    .A3(\w[12][25] ),
    .S0(net551),
    .S1(net479),
    .X(_11034_));
 sky130_fd_sc_hd__mux4_1 _25421_ (.A0(\w[18][25] ),
    .A1(\w[16][25] ),
    .A2(\w[22][25] ),
    .A3(\w[20][25] ),
    .S0(net551),
    .S1(net479),
    .X(_11035_));
 sky130_fd_sc_hd__nand2_1 _25422_ (.A(net489),
    .B(_11035_),
    .Y(_11036_));
 sky130_fd_sc_hd__mux4_1 _25423_ (.A0(\w[26][25] ),
    .A1(\w[24][25] ),
    .A2(\w[30][25] ),
    .A3(\w[28][25] ),
    .S0(net551),
    .S1(net479),
    .X(_11037_));
 sky130_fd_sc_hd__nand2_1 _25424_ (.A(net502),
    .B(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__a21oi_1 _25425_ (.A1(_11036_),
    .A2(_11038_),
    .B1(net497),
    .Y(_11039_));
 sky130_fd_sc_hd__a31oi_1 _25426_ (.A1(net497),
    .A2(net502),
    .A3(_11034_),
    .B1(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__a21oi_1 _25427_ (.A1(_11033_),
    .A2(_11040_),
    .B1(net457),
    .Y(_11041_));
 sky130_fd_sc_hd__a21oi_1 _25428_ (.A1(net457),
    .A2(_11031_),
    .B1(_11041_),
    .Y(_11042_));
 sky130_fd_sc_hd__nand2_1 _25429_ (.A(net526),
    .B(\w[0][25] ),
    .Y(_11043_));
 sky130_fd_sc_hd__o21ai_4 _25430_ (.A1(net455),
    .A2(_11042_),
    .B1(_11043_),
    .Y(_00017_));
 sky130_fd_sc_hd__mux4_1 _25431_ (.A0(\w[18][26] ),
    .A1(\w[16][26] ),
    .A2(\w[22][26] ),
    .A3(\w[20][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11044_));
 sky130_fd_sc_hd__mux4_1 _25432_ (.A0(\w[26][26] ),
    .A1(\w[24][26] ),
    .A2(\w[30][26] ),
    .A3(\w[28][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11045_));
 sky130_fd_sc_hd__mux4_1 _25433_ (.A0(\w[2][26] ),
    .A1(\w[0][26] ),
    .A2(\w[6][26] ),
    .A3(\w[4][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11046_));
 sky130_fd_sc_hd__mux4_1 _25434_ (.A0(\w[10][26] ),
    .A1(\w[8][26] ),
    .A2(\w[14][26] ),
    .A3(\w[12][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11047_));
 sky130_fd_sc_hd__mux4_1 _25435_ (.A0(_11044_),
    .A1(_11045_),
    .A2(_11046_),
    .A3(_11047_),
    .S0(net506),
    .S1(net497),
    .X(_11048_));
 sky130_fd_sc_hd__mux4_1 _25436_ (.A0(\w[34][26] ),
    .A1(\w[32][26] ),
    .A2(\w[38][26] ),
    .A3(\w[36][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11049_));
 sky130_fd_sc_hd__nand2_1 _25437_ (.A(net460),
    .B(_11049_),
    .Y(_11050_));
 sky130_fd_sc_hd__mux4_1 _25438_ (.A0(\w[42][26] ),
    .A1(\w[40][26] ),
    .A2(\w[46][26] ),
    .A3(\w[44][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11051_));
 sky130_fd_sc_hd__mux4_1 _25439_ (.A0(\w[50][26] ),
    .A1(\w[48][26] ),
    .A2(\w[54][26] ),
    .A3(\w[52][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11052_));
 sky130_fd_sc_hd__nand2_1 _25440_ (.A(net492),
    .B(_11052_),
    .Y(_11053_));
 sky130_fd_sc_hd__mux4_1 _25441_ (.A0(\w[58][26] ),
    .A1(\w[56][26] ),
    .A2(\w[62][26] ),
    .A3(\w[60][26] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11054_));
 sky130_fd_sc_hd__nand2_1 _25442_ (.A(_10499_),
    .B(_11054_),
    .Y(_11055_));
 sky130_fd_sc_hd__a21oi_1 _25443_ (.A1(_11053_),
    .A2(_11055_),
    .B1(net499),
    .Y(_11056_));
 sky130_fd_sc_hd__a31oi_1 _25444_ (.A1(net498),
    .A2(_10499_),
    .A3(_11051_),
    .B1(_11056_),
    .Y(_11057_));
 sky130_fd_sc_hd__a21oi_1 _25445_ (.A1(_11050_),
    .A2(_11057_),
    .B1(_10508_),
    .Y(_11058_));
 sky130_fd_sc_hd__a21oi_1 _25446_ (.A1(net462),
    .A2(_11048_),
    .B1(_11058_),
    .Y(_11059_));
 sky130_fd_sc_hd__nand2_1 _25447_ (.A(net526),
    .B(\w[0][26] ),
    .Y(_11060_));
 sky130_fd_sc_hd__o21ai_4 _25448_ (.A1(net455),
    .A2(_11059_),
    .B1(_11060_),
    .Y(_00018_));
 sky130_fd_sc_hd__mux4_1 _25449_ (.A0(\w[2][27] ),
    .A1(\w[0][27] ),
    .A2(\w[6][27] ),
    .A3(\w[4][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11061_));
 sky130_fd_sc_hd__mux4_1 _25450_ (.A0(\w[34][27] ),
    .A1(\w[32][27] ),
    .A2(\w[38][27] ),
    .A3(\w[36][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11062_));
 sky130_fd_sc_hd__mux2i_1 _25451_ (.A0(_11061_),
    .A1(_11062_),
    .S(net458),
    .Y(_11063_));
 sky130_fd_sc_hd__mux4_2 _25452_ (.A0(\w[10][27] ),
    .A1(\w[8][27] ),
    .A2(\w[14][27] ),
    .A3(\w[12][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11064_));
 sky130_fd_sc_hd__mux4_1 _25453_ (.A0(\w[18][27] ),
    .A1(\w[16][27] ),
    .A2(\w[22][27] ),
    .A3(\w[20][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11065_));
 sky130_fd_sc_hd__nand2_1 _25454_ (.A(net490),
    .B(_11065_),
    .Y(_11066_));
 sky130_fd_sc_hd__mux4_1 _25455_ (.A0(\w[26][27] ),
    .A1(\w[24][27] ),
    .A2(\w[30][27] ),
    .A3(\w[28][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11067_));
 sky130_fd_sc_hd__nand2_1 _25456_ (.A(net501),
    .B(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__a21oi_1 _25457_ (.A1(_11066_),
    .A2(_11068_),
    .B1(net493),
    .Y(_11069_));
 sky130_fd_sc_hd__a311oi_1 _25458_ (.A1(net493),
    .A2(net501),
    .A3(_11064_),
    .B1(_11069_),
    .C1(net458),
    .Y(_11070_));
 sky130_fd_sc_hd__mux4_1 _25459_ (.A0(\w[42][27] ),
    .A1(\w[40][27] ),
    .A2(\w[46][27] ),
    .A3(\w[44][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11071_));
 sky130_fd_sc_hd__mux4_1 _25460_ (.A0(\w[50][27] ),
    .A1(\w[48][27] ),
    .A2(\w[54][27] ),
    .A3(\w[52][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11072_));
 sky130_fd_sc_hd__nand2_1 _25461_ (.A(net490),
    .B(_11072_),
    .Y(_11073_));
 sky130_fd_sc_hd__mux4_1 _25462_ (.A0(\w[58][27] ),
    .A1(\w[56][27] ),
    .A2(\w[62][27] ),
    .A3(\w[60][27] ),
    .S0(net550),
    .S1(net478),
    .X(_11074_));
 sky130_fd_sc_hd__nand2_1 _25463_ (.A(net503),
    .B(_11074_),
    .Y(_11075_));
 sky130_fd_sc_hd__a21oi_1 _25464_ (.A1(_11073_),
    .A2(_11075_),
    .B1(net493),
    .Y(_11076_));
 sky130_fd_sc_hd__a311oi_2 _25465_ (.A1(net493),
    .A2(net503),
    .A3(_11071_),
    .B1(_11076_),
    .C1(net461),
    .Y(_11077_));
 sky130_fd_sc_hd__o22ai_1 _25466_ (.A1(_10575_),
    .A2(_11063_),
    .B1(_11070_),
    .B2(_11077_),
    .Y(_11078_));
 sky130_fd_sc_hd__a22o_1 _25467_ (.A1(net525),
    .A2(\w[0][27] ),
    .B1(_10573_),
    .B2(_11078_),
    .X(_00019_));
 sky130_fd_sc_hd__mux4_2 _25468_ (.A0(\w[2][28] ),
    .A1(\w[0][28] ),
    .A2(\w[6][28] ),
    .A3(\w[4][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11079_));
 sky130_fd_sc_hd__mux4_1 _25469_ (.A0(\w[34][28] ),
    .A1(\w[32][28] ),
    .A2(\w[38][28] ),
    .A3(\w[36][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11080_));
 sky130_fd_sc_hd__mux2i_1 _25470_ (.A0(_11079_),
    .A1(_11080_),
    .S(net458),
    .Y(_11081_));
 sky130_fd_sc_hd__mux4_1 _25471_ (.A0(\w[10][28] ),
    .A1(\w[8][28] ),
    .A2(\w[14][28] ),
    .A3(\w[12][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11082_));
 sky130_fd_sc_hd__mux4_1 _25472_ (.A0(\w[18][28] ),
    .A1(\w[16][28] ),
    .A2(\w[22][28] ),
    .A3(\w[20][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11083_));
 sky130_fd_sc_hd__nand2_1 _25473_ (.A(net490),
    .B(_11083_),
    .Y(_11084_));
 sky130_fd_sc_hd__mux4_1 _25474_ (.A0(\w[26][28] ),
    .A1(\w[24][28] ),
    .A2(\w[30][28] ),
    .A3(\w[28][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11085_));
 sky130_fd_sc_hd__nand2_1 _25475_ (.A(net501),
    .B(_11085_),
    .Y(_11086_));
 sky130_fd_sc_hd__a21oi_1 _25476_ (.A1(_11084_),
    .A2(_11086_),
    .B1(net493),
    .Y(_11087_));
 sky130_fd_sc_hd__a311oi_2 _25477_ (.A1(net493),
    .A2(net501),
    .A3(_11082_),
    .B1(_11087_),
    .C1(net458),
    .Y(_11088_));
 sky130_fd_sc_hd__mux4_1 _25478_ (.A0(\w[42][28] ),
    .A1(\w[40][28] ),
    .A2(\w[46][28] ),
    .A3(\w[44][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11089_));
 sky130_fd_sc_hd__mux4_1 _25479_ (.A0(\w[50][28] ),
    .A1(\w[48][28] ),
    .A2(\w[54][28] ),
    .A3(\w[52][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11090_));
 sky130_fd_sc_hd__nand2_1 _25480_ (.A(net490),
    .B(_11090_),
    .Y(_11091_));
 sky130_fd_sc_hd__mux4_1 _25481_ (.A0(\w[58][28] ),
    .A1(\w[56][28] ),
    .A2(\w[62][28] ),
    .A3(\w[60][28] ),
    .S0(net550),
    .S1(net478),
    .X(_11092_));
 sky130_fd_sc_hd__nand2_1 _25482_ (.A(net501),
    .B(_11092_),
    .Y(_11093_));
 sky130_fd_sc_hd__a21oi_1 _25483_ (.A1(_11091_),
    .A2(_11093_),
    .B1(net493),
    .Y(_11094_));
 sky130_fd_sc_hd__a311oi_1 _25484_ (.A1(net493),
    .A2(net501),
    .A3(_11089_),
    .B1(_11094_),
    .C1(net461),
    .Y(_11095_));
 sky130_fd_sc_hd__o22ai_1 _25485_ (.A1(_10575_),
    .A2(_11081_),
    .B1(_11088_),
    .B2(_11095_),
    .Y(_11096_));
 sky130_fd_sc_hd__a22o_1 _25486_ (.A1(net525),
    .A2(\w[0][28] ),
    .B1(_10573_),
    .B2(_11096_),
    .X(_00020_));
 sky130_fd_sc_hd__mux4_1 _25487_ (.A0(\w[18][29] ),
    .A1(\w[16][29] ),
    .A2(\w[22][29] ),
    .A3(\w[20][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11097_));
 sky130_fd_sc_hd__mux4_1 _25488_ (.A0(\w[26][29] ),
    .A1(\w[24][29] ),
    .A2(\w[30][29] ),
    .A3(\w[28][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11098_));
 sky130_fd_sc_hd__mux4_1 _25489_ (.A0(\w[2][29] ),
    .A1(\w[0][29] ),
    .A2(\w[6][29] ),
    .A3(\w[4][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11099_));
 sky130_fd_sc_hd__mux4_1 _25490_ (.A0(\w[10][29] ),
    .A1(\w[8][29] ),
    .A2(\w[14][29] ),
    .A3(\w[12][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11100_));
 sky130_fd_sc_hd__mux4_1 _25491_ (.A0(_11097_),
    .A1(_11098_),
    .A2(_11099_),
    .A3(_11100_),
    .S0(net506),
    .S1(net497),
    .X(_11101_));
 sky130_fd_sc_hd__mux4_1 _25492_ (.A0(\w[34][29] ),
    .A1(\w[32][29] ),
    .A2(\w[38][29] ),
    .A3(\w[36][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11102_));
 sky130_fd_sc_hd__nand2_1 _25493_ (.A(net460),
    .B(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__mux4_1 _25494_ (.A0(\w[42][29] ),
    .A1(\w[40][29] ),
    .A2(\w[46][29] ),
    .A3(\w[44][29] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_11104_));
 sky130_fd_sc_hd__mux4_1 _25495_ (.A0(\w[50][29] ),
    .A1(\w[48][29] ),
    .A2(\w[54][29] ),
    .A3(\w[52][29] ),
    .S0(\count_hash1[1] ),
    .S1(net481),
    .X(_11105_));
 sky130_fd_sc_hd__nand2_1 _25496_ (.A(net491),
    .B(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__mux4_1 _25497_ (.A0(\w[58][29] ),
    .A1(\w[56][29] ),
    .A2(\w[62][29] ),
    .A3(\w[60][29] ),
    .S0(\count_hash1[1] ),
    .S1(net481),
    .X(_11107_));
 sky130_fd_sc_hd__nand2_1 _25498_ (.A(net506),
    .B(_11107_),
    .Y(_11108_));
 sky130_fd_sc_hd__a21oi_1 _25499_ (.A1(_11106_),
    .A2(_11108_),
    .B1(net498),
    .Y(_11109_));
 sky130_fd_sc_hd__a31oi_1 _25500_ (.A1(net498),
    .A2(net506),
    .A3(_11104_),
    .B1(_11109_),
    .Y(_11110_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__a21oi_1 _25503_ (.A1(_11103_),
    .A2(_11110_),
    .B1(net462),
    .Y(_11113_));
 sky130_fd_sc_hd__a21oi_1 _25504_ (.A1(net462),
    .A2(_11101_),
    .B1(_11113_),
    .Y(_11114_));
 sky130_fd_sc_hd__nand2_1 _25505_ (.A(net526),
    .B(\w[0][29] ),
    .Y(_11115_));
 sky130_fd_sc_hd__o21ai_4 _25506_ (.A1(net455),
    .A2(_11114_),
    .B1(_11115_),
    .Y(_00021_));
 sky130_fd_sc_hd__mux4_1 _25507_ (.A0(\w[18][30] ),
    .A1(\w[16][30] ),
    .A2(\w[22][30] ),
    .A3(\w[20][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11116_));
 sky130_fd_sc_hd__mux4_1 _25508_ (.A0(\w[26][30] ),
    .A1(\w[24][30] ),
    .A2(\w[30][30] ),
    .A3(\w[28][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11117_));
 sky130_fd_sc_hd__mux4_1 _25509_ (.A0(\w[2][30] ),
    .A1(\w[0][30] ),
    .A2(\w[6][30] ),
    .A3(\w[4][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11118_));
 sky130_fd_sc_hd__mux4_1 _25510_ (.A0(\w[10][30] ),
    .A1(\w[8][30] ),
    .A2(\w[14][30] ),
    .A3(\w[12][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11119_));
 sky130_fd_sc_hd__mux4_1 _25511_ (.A0(_11116_),
    .A1(_11117_),
    .A2(_11118_),
    .A3(_11119_),
    .S0(net504),
    .S1(net496),
    .X(_11120_));
 sky130_fd_sc_hd__mux4_1 _25512_ (.A0(\w[50][30] ),
    .A1(\w[48][30] ),
    .A2(\w[54][30] ),
    .A3(\w[52][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11121_));
 sky130_fd_sc_hd__mux4_1 _25513_ (.A0(\w[58][30] ),
    .A1(\w[56][30] ),
    .A2(\w[62][30] ),
    .A3(\w[60][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11122_));
 sky130_fd_sc_hd__mux4_1 _25514_ (.A0(\w[34][30] ),
    .A1(\w[32][30] ),
    .A2(\w[38][30] ),
    .A3(\w[36][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11123_));
 sky130_fd_sc_hd__mux4_1 _25515_ (.A0(\w[42][30] ),
    .A1(\w[40][30] ),
    .A2(\w[46][30] ),
    .A3(\w[44][30] ),
    .S0(net546),
    .S1(net480),
    .X(_11124_));
 sky130_fd_sc_hd__mux4_1 _25516_ (.A0(_11121_),
    .A1(_11122_),
    .A2(_11123_),
    .A3(_11124_),
    .S0(net504),
    .S1(net499),
    .X(_11125_));
 sky130_fd_sc_hd__mux2i_2 _25517_ (.A0(_11120_),
    .A1(_11125_),
    .S(net456),
    .Y(_11126_));
 sky130_fd_sc_hd__nand2_1 _25518_ (.A(net526),
    .B(\w[0][30] ),
    .Y(_11127_));
 sky130_fd_sc_hd__o21ai_4 _25519_ (.A1(net453),
    .A2(_11126_),
    .B1(_11127_),
    .Y(_00023_));
 sky130_fd_sc_hd__mux4_2 _25520_ (.A0(\w[2][31] ),
    .A1(\w[0][31] ),
    .A2(\w[6][31] ),
    .A3(\w[4][31] ),
    .S0(net550),
    .S1(net478),
    .X(_11128_));
 sky130_fd_sc_hd__mux4_1 _25521_ (.A0(\w[34][31] ),
    .A1(\w[32][31] ),
    .A2(\w[38][31] ),
    .A3(\w[36][31] ),
    .S0(net549),
    .S1(net477),
    .X(_11129_));
 sky130_fd_sc_hd__mux2i_1 _25522_ (.A0(_11128_),
    .A1(_11129_),
    .S(net458),
    .Y(_11130_));
 sky130_fd_sc_hd__mux4_1 _25523_ (.A0(\w[10][31] ),
    .A1(\w[8][31] ),
    .A2(\w[14][31] ),
    .A3(\w[12][31] ),
    .S0(net550),
    .S1(net478),
    .X(_11131_));
 sky130_fd_sc_hd__mux4_1 _25524_ (.A0(\w[18][31] ),
    .A1(\w[16][31] ),
    .A2(\w[22][31] ),
    .A3(\w[20][31] ),
    .S0(net550),
    .S1(net478),
    .X(_11132_));
 sky130_fd_sc_hd__nand2_1 _25525_ (.A(net490),
    .B(_11132_),
    .Y(_11133_));
 sky130_fd_sc_hd__mux4_1 _25526_ (.A0(\w[26][31] ),
    .A1(\w[24][31] ),
    .A2(\w[30][31] ),
    .A3(\w[28][31] ),
    .S0(net550),
    .S1(net478),
    .X(_11134_));
 sky130_fd_sc_hd__nand2_1 _25527_ (.A(net501),
    .B(_11134_),
    .Y(_11135_));
 sky130_fd_sc_hd__a21oi_1 _25528_ (.A1(_11133_),
    .A2(_11135_),
    .B1(net493),
    .Y(_11136_));
 sky130_fd_sc_hd__a311oi_2 _25529_ (.A1(net493),
    .A2(net501),
    .A3(_11131_),
    .B1(_11136_),
    .C1(net458),
    .Y(_11137_));
 sky130_fd_sc_hd__mux4_1 _25530_ (.A0(\w[42][31] ),
    .A1(\w[40][31] ),
    .A2(\w[46][31] ),
    .A3(\w[44][31] ),
    .S0(net549),
    .S1(net477),
    .X(_11138_));
 sky130_fd_sc_hd__mux4_1 _25531_ (.A0(\w[50][31] ),
    .A1(\w[48][31] ),
    .A2(\w[54][31] ),
    .A3(\w[52][31] ),
    .S0(net549),
    .S1(net477),
    .X(_11139_));
 sky130_fd_sc_hd__nand2_1 _25532_ (.A(net489),
    .B(_11139_),
    .Y(_11140_));
 sky130_fd_sc_hd__mux4_1 _25533_ (.A0(\w[58][31] ),
    .A1(\w[56][31] ),
    .A2(\w[62][31] ),
    .A3(\w[60][31] ),
    .S0(net549),
    .S1(net477),
    .X(_11141_));
 sky130_fd_sc_hd__nand2_1 _25534_ (.A(net503),
    .B(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__a21oi_1 _25535_ (.A1(_11140_),
    .A2(_11142_),
    .B1(net494),
    .Y(_11143_));
 sky130_fd_sc_hd__a311oi_4 _25536_ (.A1(net494),
    .A2(net503),
    .A3(_11138_),
    .B1(_11143_),
    .C1(net461),
    .Y(_11144_));
 sky130_fd_sc_hd__o22ai_1 _25537_ (.A1(_10575_),
    .A2(_11130_),
    .B1(_11137_),
    .B2(_11144_),
    .Y(_11145_));
 sky130_fd_sc_hd__a22o_2 _25538_ (.A1(net525),
    .A2(\w[0][31] ),
    .B1(_10573_),
    .B2(_11145_),
    .X(_00024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_386 ();
 sky130_fd_sc_hd__mux4_1 _25548_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(\count15_1[2] ),
    .S1(net697),
    .X(_11155_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_382 ();
 sky130_fd_sc_hd__mux4_1 _25553_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11160_));
 sky130_fd_sc_hd__mux4_1 _25554_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(\count15_1[2] ),
    .S1(net697),
    .X(_11161_));
 sky130_fd_sc_hd__mux4_1 _25555_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(\count15_1[2] ),
    .S1(net697),
    .X(_11162_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_377 ();
 sky130_fd_sc_hd__mux4_4 _25561_ (.A0(_11155_),
    .A1(_11160_),
    .A2(_11161_),
    .A3(_11162_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11168_));
 sky130_fd_sc_hd__mux4_1 _25562_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net692),
    .S1(net699),
    .X(_11169_));
 sky130_fd_sc_hd__mux4_1 _25563_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net692),
    .S1(net699),
    .X(_11170_));
 sky130_fd_sc_hd__mux4_1 _25564_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net692),
    .S1(\count15_1[1] ),
    .X(_11171_));
 sky130_fd_sc_hd__mux4_1 _25565_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net692),
    .S1(\count15_1[1] ),
    .X(_11172_));
 sky130_fd_sc_hd__mux4_1 _25566_ (.A0(_11169_),
    .A1(_11170_),
    .A2(_11171_),
    .A3(_11172_),
    .S0(net687),
    .S1(net685),
    .X(_11173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_375 ();
 sky130_fd_sc_hd__mux2i_4 _25569_ (.A0(_11168_),
    .A1(_11173_),
    .S(net683),
    .Y(_11176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_372 ();
 sky130_fd_sc_hd__mux4_1 _25573_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net693),
    .S1(net698),
    .X(_11180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_370 ();
 sky130_fd_sc_hd__mux4_1 _25576_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net693),
    .S1(net698),
    .X(_11183_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_368 ();
 sky130_fd_sc_hd__mux4_1 _25579_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net693),
    .S1(net698),
    .X(_11186_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_366 ();
 sky130_fd_sc_hd__mux4_1 _25582_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net693),
    .S1(net698),
    .X(_11189_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_364 ();
 sky130_fd_sc_hd__mux4_4 _25585_ (.A0(_11180_),
    .A1(_11183_),
    .A2(_11186_),
    .A3(_11189_),
    .S0(net688),
    .S1(net686),
    .X(_11192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_363 ();
 sky130_fd_sc_hd__mux4_1 _25587_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net694),
    .S1(net699),
    .X(_11194_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_361 ();
 sky130_fd_sc_hd__mux4_1 _25590_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net694),
    .S1(net699),
    .X(_11197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_359 ();
 sky130_fd_sc_hd__mux4_1 _25593_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net694),
    .S1(net699),
    .X(_11200_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 ();
 sky130_fd_sc_hd__mux4_1 _25596_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net694),
    .S1(net699),
    .X(_11203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 ();
 sky130_fd_sc_hd__mux4_1 _25599_ (.A0(_11194_),
    .A1(_11197_),
    .A2(_11200_),
    .A3(_11203_),
    .S0(net688),
    .S1(net686),
    .X(_11206_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 ();
 sky130_fd_sc_hd__mux2i_4 _25601_ (.A0(_11192_),
    .A1(_11206_),
    .S(net684),
    .Y(_11208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 ();
 sky130_fd_sc_hd__mux4_1 _25604_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net690),
    .S1(net697),
    .X(_11211_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_351 ();
 sky130_fd_sc_hd__mux4_1 _25606_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net690),
    .S1(\count15_1[1] ),
    .X(_11213_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_349 ();
 sky130_fd_sc_hd__mux4_1 _25609_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net690),
    .S1(net697),
    .X(_11216_));
 sky130_fd_sc_hd__mux4_1 _25610_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net690),
    .S1(net697),
    .X(_11217_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_348 ();
 sky130_fd_sc_hd__mux4_4 _25612_ (.A0(_11211_),
    .A1(_11213_),
    .A2(_11216_),
    .A3(_11217_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11219_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_346 ();
 sky130_fd_sc_hd__mux4_1 _25615_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net691),
    .S1(net700),
    .X(_11222_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_344 ();
 sky130_fd_sc_hd__mux4_1 _25618_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net691),
    .S1(net700),
    .X(_11225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_343 ();
 sky130_fd_sc_hd__mux4_1 _25620_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net691),
    .S1(net700),
    .X(_11227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_341 ();
 sky130_fd_sc_hd__mux4_1 _25623_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net691),
    .S1(net700),
    .X(_11230_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_339 ();
 sky130_fd_sc_hd__mux4_1 _25626_ (.A0(_11222_),
    .A1(_11225_),
    .A2(_11227_),
    .A3(_11230_),
    .S0(net687),
    .S1(net685),
    .X(_11233_));
 sky130_fd_sc_hd__mux2i_4 _25627_ (.A0(_11219_),
    .A1(_11233_),
    .S(net683),
    .Y(_11234_));
 sky130_fd_sc_hd__xnor2_1 _25628_ (.A(_11208_),
    .B(_11234_),
    .Y(_11235_));
 sky130_fd_sc_hd__xnor2_2 _25629_ (.A(_11176_),
    .B(_11235_),
    .Y(_11750_));
 sky130_fd_sc_hd__mux4_1 _25630_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net693),
    .S1(net698),
    .X(_11236_));
 sky130_fd_sc_hd__mux4_1 _25631_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net693),
    .S1(net698),
    .X(_11237_));
 sky130_fd_sc_hd__mux4_1 _25632_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net693),
    .S1(net698),
    .X(_11238_));
 sky130_fd_sc_hd__mux4_1 _25633_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net693),
    .S1(net698),
    .X(_11239_));
 sky130_fd_sc_hd__mux4_4 _25634_ (.A0(_11236_),
    .A1(_11237_),
    .A2(_11238_),
    .A3(_11239_),
    .S0(net688),
    .S1(net686),
    .X(_11240_));
 sky130_fd_sc_hd__mux4_1 _25635_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net696),
    .S1(net701),
    .X(_11241_));
 sky130_fd_sc_hd__mux4_1 _25636_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net696),
    .S1(net701),
    .X(_11242_));
 sky130_fd_sc_hd__mux4_1 _25637_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net696),
    .S1(net701),
    .X(_11243_));
 sky130_fd_sc_hd__mux4_1 _25638_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net696),
    .S1(net701),
    .X(_11244_));
 sky130_fd_sc_hd__mux4_1 _25639_ (.A0(_11241_),
    .A1(_11242_),
    .A2(_11243_),
    .A3(_11244_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11245_));
 sky130_fd_sc_hd__mux2i_4 _25640_ (.A0(_11240_),
    .A1(_11245_),
    .S(net684),
    .Y(_11246_));
 sky130_fd_sc_hd__mux4_1 _25641_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11247_));
 sky130_fd_sc_hd__mux4_1 _25642_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11248_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_338 ();
 sky130_fd_sc_hd__mux4_1 _25644_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11250_));
 sky130_fd_sc_hd__mux4_1 _25645_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11251_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_337 ();
 sky130_fd_sc_hd__mux4_4 _25647_ (.A0(_11247_),
    .A1(_11248_),
    .A2(_11250_),
    .A3(_11251_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11253_));
 sky130_fd_sc_hd__mux4_1 _25648_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(\count15_1[2] ),
    .S1(net701),
    .X(_11254_));
 sky130_fd_sc_hd__mux4_1 _25649_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net692),
    .S1(net701),
    .X(_11255_));
 sky130_fd_sc_hd__mux4_1 _25650_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(\count15_1[2] ),
    .S1(net701),
    .X(_11256_));
 sky130_fd_sc_hd__mux4_1 _25651_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(\count15_1[2] ),
    .S1(net701),
    .X(_11257_));
 sky130_fd_sc_hd__mux4_1 _25652_ (.A0(_11254_),
    .A1(_11255_),
    .A2(_11256_),
    .A3(_11257_),
    .S0(net687),
    .S1(net685),
    .X(_11258_));
 sky130_fd_sc_hd__mux2i_4 _25653_ (.A0(_11253_),
    .A1(_11258_),
    .S(net683),
    .Y(_11259_));
 sky130_fd_sc_hd__mux4_1 _25654_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net691),
    .S1(net697),
    .X(_11260_));
 sky130_fd_sc_hd__mux4_1 _25655_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net691),
    .S1(net697),
    .X(_11261_));
 sky130_fd_sc_hd__mux4_1 _25656_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net691),
    .S1(net697),
    .X(_11262_));
 sky130_fd_sc_hd__mux4_1 _25657_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net691),
    .S1(net697),
    .X(_11263_));
 sky130_fd_sc_hd__mux4_4 _25658_ (.A0(_11260_),
    .A1(_11261_),
    .A2(_11262_),
    .A3(_11263_),
    .S0(net688),
    .S1(net686),
    .X(_11264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_336 ();
 sky130_fd_sc_hd__mux4_1 _25660_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net692),
    .S1(net699),
    .X(_11266_));
 sky130_fd_sc_hd__mux4_1 _25661_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net692),
    .S1(net699),
    .X(_11267_));
 sky130_fd_sc_hd__mux4_1 _25662_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net692),
    .S1(net699),
    .X(_11268_));
 sky130_fd_sc_hd__mux4_1 _25663_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net692),
    .S1(net699),
    .X(_11269_));
 sky130_fd_sc_hd__mux4_1 _25664_ (.A0(_11266_),
    .A1(_11267_),
    .A2(_11268_),
    .A3(_11269_),
    .S0(net687),
    .S1(net685),
    .X(_11270_));
 sky130_fd_sc_hd__mux2i_4 _25665_ (.A0(_11264_),
    .A1(_11270_),
    .S(net683),
    .Y(_11271_));
 sky130_fd_sc_hd__xnor2_1 _25666_ (.A(_11259_),
    .B(_11271_),
    .Y(_11272_));
 sky130_fd_sc_hd__xnor2_2 _25667_ (.A(_11246_),
    .B(_11272_),
    .Y(_11755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_326 ();
 sky130_fd_sc_hd__mux4_1 _25678_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11283_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_324 ();
 sky130_fd_sc_hd__mux4_1 _25681_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11286_));
 sky130_fd_sc_hd__mux4_1 _25682_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_322 ();
 sky130_fd_sc_hd__mux4_1 _25685_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_317 ();
 sky130_fd_sc_hd__mux4_4 _25691_ (.A0(_11283_),
    .A1(_11286_),
    .A2(_11287_),
    .A3(_11290_),
    .S0(net617),
    .S1(net613),
    .X(_11296_));
 sky130_fd_sc_hd__mux4_1 _25692_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_315 ();
 sky130_fd_sc_hd__mux4_1 _25695_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11300_));
 sky130_fd_sc_hd__mux4_1 _25696_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11301_));
 sky130_fd_sc_hd__mux4_1 _25697_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net621),
    .S1(net625),
    .X(_11302_));
 sky130_fd_sc_hd__mux4_1 _25698_ (.A0(_11297_),
    .A1(_11300_),
    .A2(_11301_),
    .A3(_11302_),
    .S0(net617),
    .S1(net613),
    .X(_11303_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_313 ();
 sky130_fd_sc_hd__mux2i_4 _25701_ (.A0(_11296_),
    .A1(_11303_),
    .S(net610),
    .Y(_11306_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_310 ();
 sky130_fd_sc_hd__mux4_1 _25705_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net618),
    .S1(net626),
    .X(_11310_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_308 ();
 sky130_fd_sc_hd__mux4_1 _25708_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net618),
    .S1(net626),
    .X(_11313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_306 ();
 sky130_fd_sc_hd__mux4_1 _25711_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net618),
    .S1(net626),
    .X(_11316_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_304 ();
 sky130_fd_sc_hd__mux4_1 _25714_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net618),
    .S1(net626),
    .X(_11319_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_302 ();
 sky130_fd_sc_hd__mux4_4 _25717_ (.A0(_11310_),
    .A1(_11313_),
    .A2(_11316_),
    .A3(_11319_),
    .S0(net615),
    .S1(net612),
    .X(_11322_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_300 ();
 sky130_fd_sc_hd__mux4_1 _25720_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net619),
    .S1(net627),
    .X(_11325_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_299 ();
 sky130_fd_sc_hd__mux4_1 _25722_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net619),
    .S1(net627),
    .X(_11327_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_297 ();
 sky130_fd_sc_hd__mux4_1 _25725_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net619),
    .S1(net627),
    .X(_11330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_295 ();
 sky130_fd_sc_hd__mux4_1 _25728_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net619),
    .S1(net627),
    .X(_11333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_293 ();
 sky130_fd_sc_hd__mux4_1 _25731_ (.A0(_11325_),
    .A1(_11327_),
    .A2(_11330_),
    .A3(_11333_),
    .S0(net615),
    .S1(net612),
    .X(_11336_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_292 ();
 sky130_fd_sc_hd__mux2i_4 _25733_ (.A0(_11322_),
    .A1(_11336_),
    .S(net610),
    .Y(_11338_));
 sky130_fd_sc_hd__mux4_1 _25734_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11339_));
 sky130_fd_sc_hd__mux4_1 _25735_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11340_));
 sky130_fd_sc_hd__mux4_1 _25736_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11341_));
 sky130_fd_sc_hd__mux4_1 _25737_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11342_));
 sky130_fd_sc_hd__mux4_4 _25738_ (.A0(_11339_),
    .A1(_11340_),
    .A2(_11341_),
    .A3(_11342_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11343_));
 sky130_fd_sc_hd__mux4_1 _25739_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11344_));
 sky130_fd_sc_hd__mux4_1 _25740_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11345_));
 sky130_fd_sc_hd__mux4_1 _25741_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11346_));
 sky130_fd_sc_hd__mux4_1 _25742_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11347_));
 sky130_fd_sc_hd__mux4_1 _25743_ (.A0(_11344_),
    .A1(_11345_),
    .A2(_11346_),
    .A3(_11347_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11348_));
 sky130_fd_sc_hd__mux2i_4 _25744_ (.A0(_11343_),
    .A1(_11348_),
    .S(\count2_1[5] ),
    .Y(_11349_));
 sky130_fd_sc_hd__xnor2_1 _25745_ (.A(_11338_),
    .B(_11349_),
    .Y(_11350_));
 sky130_fd_sc_hd__xnor2_1 _25746_ (.A(_11306_),
    .B(_11350_),
    .Y(_11760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_291 ();
 sky130_fd_sc_hd__mux4_1 _25748_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11352_));
 sky130_fd_sc_hd__mux4_1 _25749_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11353_));
 sky130_fd_sc_hd__mux4_1 _25750_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11354_));
 sky130_fd_sc_hd__mux4_1 _25751_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11355_));
 sky130_fd_sc_hd__mux4_2 _25752_ (.A0(_11352_),
    .A1(_11353_),
    .A2(_11354_),
    .A3(_11355_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11356_));
 sky130_fd_sc_hd__mux4_1 _25753_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11357_));
 sky130_fd_sc_hd__mux4_1 _25754_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11358_));
 sky130_fd_sc_hd__mux4_1 _25755_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11359_));
 sky130_fd_sc_hd__mux4_1 _25756_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net696),
    .S1(net701),
    .X(_11360_));
 sky130_fd_sc_hd__mux4_1 _25757_ (.A0(_11357_),
    .A1(_11358_),
    .A2(_11359_),
    .A3(_11360_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11361_));
 sky130_fd_sc_hd__mux2i_4 _25758_ (.A0(_11356_),
    .A1(_11361_),
    .S(net684),
    .Y(_11362_));
 sky130_fd_sc_hd__mux4_1 _25759_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net690),
    .S1(net697),
    .X(_11363_));
 sky130_fd_sc_hd__mux4_1 _25760_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net690),
    .S1(\count15_1[1] ),
    .X(_11364_));
 sky130_fd_sc_hd__mux4_1 _25761_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net690),
    .S1(net697),
    .X(_11365_));
 sky130_fd_sc_hd__mux4_1 _25762_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net690),
    .S1(net697),
    .X(_11366_));
 sky130_fd_sc_hd__mux4_4 _25763_ (.A0(_11363_),
    .A1(_11364_),
    .A2(_11365_),
    .A3(_11366_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11367_));
 sky130_fd_sc_hd__mux4_1 _25764_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net692),
    .S1(net700),
    .X(_11368_));
 sky130_fd_sc_hd__mux4_1 _25765_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net692),
    .S1(net700),
    .X(_11369_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_290 ();
 sky130_fd_sc_hd__mux4_1 _25767_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net690),
    .S1(net700),
    .X(_11371_));
 sky130_fd_sc_hd__mux4_1 _25768_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net692),
    .S1(net700),
    .X(_11372_));
 sky130_fd_sc_hd__mux4_1 _25769_ (.A0(_11368_),
    .A1(_11369_),
    .A2(_11371_),
    .A3(_11372_),
    .S0(net687),
    .S1(net685),
    .X(_11373_));
 sky130_fd_sc_hd__mux2i_4 _25770_ (.A0(_11367_),
    .A1(_11373_),
    .S(net683),
    .Y(_11374_));
 sky130_fd_sc_hd__mux4_1 _25771_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net695),
    .S1(net699),
    .X(_11375_));
 sky130_fd_sc_hd__mux4_1 _25772_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net695),
    .S1(net699),
    .X(_11376_));
 sky130_fd_sc_hd__mux4_1 _25773_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net695),
    .S1(net699),
    .X(_11377_));
 sky130_fd_sc_hd__mux4_1 _25774_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net695),
    .S1(net699),
    .X(_11378_));
 sky130_fd_sc_hd__mux4_4 _25775_ (.A0(_11375_),
    .A1(_11376_),
    .A2(_11377_),
    .A3(_11378_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11379_));
 sky130_fd_sc_hd__mux4_1 _25776_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net695),
    .S1(net701),
    .X(_11380_));
 sky130_fd_sc_hd__mux4_1 _25777_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net695),
    .S1(net701),
    .X(_11381_));
 sky130_fd_sc_hd__mux4_1 _25778_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net695),
    .S1(net701),
    .X(_11382_));
 sky130_fd_sc_hd__mux4_1 _25779_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net695),
    .S1(net701),
    .X(_11383_));
 sky130_fd_sc_hd__mux4_1 _25780_ (.A0(_11380_),
    .A1(_11381_),
    .A2(_11382_),
    .A3(_11383_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11384_));
 sky130_fd_sc_hd__mux2i_4 _25781_ (.A0(_11379_),
    .A1(_11384_),
    .S(net684),
    .Y(_11385_));
 sky130_fd_sc_hd__xnor2_1 _25782_ (.A(_11374_),
    .B(_11385_),
    .Y(_11386_));
 sky130_fd_sc_hd__xnor2_2 _25783_ (.A(_11362_),
    .B(_11386_),
    .Y(_11763_));
 sky130_fd_sc_hd__mux4_1 _25784_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11387_));
 sky130_fd_sc_hd__mux4_1 _25785_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11388_));
 sky130_fd_sc_hd__mux4_1 _25786_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11389_));
 sky130_fd_sc_hd__mux4_1 _25787_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11390_));
 sky130_fd_sc_hd__mux4_4 _25788_ (.A0(_11387_),
    .A1(_11388_),
    .A2(_11389_),
    .A3(_11390_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11391_));
 sky130_fd_sc_hd__mux4_1 _25789_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net620),
    .S1(net624),
    .X(_11392_));
 sky130_fd_sc_hd__mux4_1 _25790_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net620),
    .S1(net624),
    .X(_11393_));
 sky130_fd_sc_hd__mux4_1 _25791_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net620),
    .S1(net624),
    .X(_11394_));
 sky130_fd_sc_hd__mux4_1 _25792_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net620),
    .S1(net624),
    .X(_11395_));
 sky130_fd_sc_hd__mux4_1 _25793_ (.A0(_11392_),
    .A1(_11393_),
    .A2(_11394_),
    .A3(_11395_),
    .S0(net616),
    .S1(\count2_1[4] ),
    .X(_11396_));
 sky130_fd_sc_hd__mux2i_4 _25794_ (.A0(_11391_),
    .A1(_11396_),
    .S(\count2_1[5] ),
    .Y(_11397_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_289 ();
 sky130_fd_sc_hd__mux4_1 _25796_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net620),
    .S1(net627),
    .X(_11399_));
 sky130_fd_sc_hd__mux4_1 _25797_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net620),
    .S1(net627),
    .X(_11400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_288 ();
 sky130_fd_sc_hd__mux4_1 _25799_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net620),
    .S1(net627),
    .X(_11402_));
 sky130_fd_sc_hd__mux4_1 _25800_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net620),
    .S1(net627),
    .X(_11403_));
 sky130_fd_sc_hd__mux4_4 _25801_ (.A0(_11399_),
    .A1(_11400_),
    .A2(_11402_),
    .A3(_11403_),
    .S0(net616),
    .S1(net614),
    .X(_11404_));
 sky130_fd_sc_hd__mux4_1 _25802_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net619),
    .S1(net627),
    .X(_11405_));
 sky130_fd_sc_hd__mux4_1 _25803_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net620),
    .S1(net627),
    .X(_11406_));
 sky130_fd_sc_hd__mux4_1 _25804_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net620),
    .S1(net627),
    .X(_11407_));
 sky130_fd_sc_hd__mux4_1 _25805_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net620),
    .S1(net627),
    .X(_11408_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_287 ();
 sky130_fd_sc_hd__mux4_1 _25807_ (.A0(_11405_),
    .A1(_11406_),
    .A2(_11407_),
    .A3(_11408_),
    .S0(net616),
    .S1(net614),
    .X(_11410_));
 sky130_fd_sc_hd__mux2i_4 _25808_ (.A0(_11404_),
    .A1(_11410_),
    .S(net611),
    .Y(_11411_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_286 ();
 sky130_fd_sc_hd__mux4_1 _25810_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net618),
    .S1(net626),
    .X(_11413_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_285 ();
 sky130_fd_sc_hd__mux4_1 _25812_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net618),
    .S1(net626),
    .X(_11415_));
 sky130_fd_sc_hd__mux4_1 _25813_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net618),
    .S1(net626),
    .X(_11416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_283 ();
 sky130_fd_sc_hd__mux4_1 _25816_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net618),
    .S1(net626),
    .X(_11419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_281 ();
 sky130_fd_sc_hd__mux4_4 _25819_ (.A0(_11413_),
    .A1(_11415_),
    .A2(_11416_),
    .A3(_11419_),
    .S0(net616),
    .S1(net614),
    .X(_11422_));
 sky130_fd_sc_hd__mux4_1 _25820_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net619),
    .S1(net627),
    .X(_11423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_279 ();
 sky130_fd_sc_hd__mux4_1 _25823_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net619),
    .S1(net627),
    .X(_11426_));
 sky130_fd_sc_hd__mux4_1 _25824_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net619),
    .S1(net627),
    .X(_11427_));
 sky130_fd_sc_hd__mux4_1 _25825_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net619),
    .S1(net627),
    .X(_11428_));
 sky130_fd_sc_hd__mux4_1 _25826_ (.A0(_11423_),
    .A1(_11426_),
    .A2(_11427_),
    .A3(_11428_),
    .S0(net615),
    .S1(net612),
    .X(_11429_));
 sky130_fd_sc_hd__mux2i_4 _25827_ (.A0(_11422_),
    .A1(_11429_),
    .S(net611),
    .Y(_11430_));
 sky130_fd_sc_hd__xnor2_1 _25828_ (.A(_11411_),
    .B(_11430_),
    .Y(_11431_));
 sky130_fd_sc_hd__xnor2_1 _25829_ (.A(_11397_),
    .B(_11431_),
    .Y(_11768_));
 sky130_fd_sc_hd__mux4_1 _25830_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net693),
    .S1(net698),
    .X(_11432_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_278 ();
 sky130_fd_sc_hd__mux4_1 _25832_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net693),
    .S1(net698),
    .X(_11434_));
 sky130_fd_sc_hd__mux4_1 _25833_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net693),
    .S1(net698),
    .X(_11435_));
 sky130_fd_sc_hd__mux4_1 _25834_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net693),
    .S1(net698),
    .X(_11436_));
 sky130_fd_sc_hd__mux4_4 _25835_ (.A0(_11432_),
    .A1(_11434_),
    .A2(_11435_),
    .A3(_11436_),
    .S0(net688),
    .S1(net686),
    .X(_11437_));
 sky130_fd_sc_hd__mux4_1 _25836_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net696),
    .S1(net701),
    .X(_11438_));
 sky130_fd_sc_hd__mux4_1 _25837_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net694),
    .S1(net701),
    .X(_11439_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_277 ();
 sky130_fd_sc_hd__mux4_1 _25839_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net696),
    .S1(net701),
    .X(_11441_));
 sky130_fd_sc_hd__mux4_1 _25840_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net696),
    .S1(net701),
    .X(_11442_));
 sky130_fd_sc_hd__mux4_1 _25841_ (.A0(_11438_),
    .A1(_11439_),
    .A2(_11441_),
    .A3(_11442_),
    .S0(net688),
    .S1(net686),
    .X(_11443_));
 sky130_fd_sc_hd__mux2i_4 _25842_ (.A0(_11437_),
    .A1(_11443_),
    .S(net684),
    .Y(_11444_));
 sky130_fd_sc_hd__mux4_1 _25843_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net694),
    .S1(net698),
    .X(_11445_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_275 ();
 sky130_fd_sc_hd__mux4_1 _25846_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net694),
    .S1(net698),
    .X(_11448_));
 sky130_fd_sc_hd__mux4_1 _25847_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net694),
    .S1(net698),
    .X(_11449_));
 sky130_fd_sc_hd__mux4_1 _25848_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net694),
    .S1(net698),
    .X(_11450_));
 sky130_fd_sc_hd__mux4_4 _25849_ (.A0(_11445_),
    .A1(_11448_),
    .A2(_11449_),
    .A3(_11450_),
    .S0(net688),
    .S1(net686),
    .X(_11451_));
 sky130_fd_sc_hd__mux4_1 _25850_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net696),
    .S1(net699),
    .X(_11452_));
 sky130_fd_sc_hd__mux4_1 _25851_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net696),
    .S1(net699),
    .X(_11453_));
 sky130_fd_sc_hd__mux4_1 _25852_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net696),
    .S1(net699),
    .X(_11454_));
 sky130_fd_sc_hd__mux4_1 _25853_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net696),
    .S1(net699),
    .X(_11455_));
 sky130_fd_sc_hd__mux4_1 _25854_ (.A0(_11452_),
    .A1(_11453_),
    .A2(_11454_),
    .A3(_11455_),
    .S0(net688),
    .S1(net686),
    .X(_11456_));
 sky130_fd_sc_hd__mux2i_4 _25855_ (.A0(_11451_),
    .A1(_11456_),
    .S(net684),
    .Y(_11457_));
 sky130_fd_sc_hd__mux4_1 _25856_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net695),
    .S1(net699),
    .X(_11458_));
 sky130_fd_sc_hd__mux4_1 _25857_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net695),
    .S1(net699),
    .X(_11459_));
 sky130_fd_sc_hd__mux4_1 _25858_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net695),
    .S1(net699),
    .X(_11460_));
 sky130_fd_sc_hd__mux4_1 _25859_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net695),
    .S1(net699),
    .X(_11461_));
 sky130_fd_sc_hd__mux4_4 _25860_ (.A0(_11458_),
    .A1(_11459_),
    .A2(_11460_),
    .A3(_11461_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11462_));
 sky130_fd_sc_hd__mux4_1 _25861_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net693),
    .S1(net699),
    .X(_11463_));
 sky130_fd_sc_hd__mux4_1 _25862_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net693),
    .S1(net699),
    .X(_11464_));
 sky130_fd_sc_hd__mux4_1 _25863_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net693),
    .S1(net699),
    .X(_11465_));
 sky130_fd_sc_hd__mux4_1 _25864_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net693),
    .S1(net699),
    .X(_11466_));
 sky130_fd_sc_hd__mux4_1 _25865_ (.A0(_11463_),
    .A1(_11464_),
    .A2(_11465_),
    .A3(_11466_),
    .S0(net688),
    .S1(net686),
    .X(_11467_));
 sky130_fd_sc_hd__mux2i_4 _25866_ (.A0(_11462_),
    .A1(_11467_),
    .S(net684),
    .Y(_11468_));
 sky130_fd_sc_hd__xnor2_1 _25867_ (.A(_11457_),
    .B(_11468_),
    .Y(_11469_));
 sky130_fd_sc_hd__xnor2_2 _25868_ (.A(_11444_),
    .B(_11469_),
    .Y(_11774_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_274 ();
 sky130_fd_sc_hd__mux4_1 _25870_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11471_));
 sky130_fd_sc_hd__mux4_1 _25871_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11472_));
 sky130_fd_sc_hd__mux4_1 _25872_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11473_));
 sky130_fd_sc_hd__mux4_1 _25873_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11474_));
 sky130_fd_sc_hd__mux4_4 _25874_ (.A0(_11471_),
    .A1(_11472_),
    .A2(_11473_),
    .A3(_11474_),
    .S0(net615),
    .S1(net612),
    .X(_11475_));
 sky130_fd_sc_hd__mux4_1 _25875_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_272 ();
 sky130_fd_sc_hd__mux4_1 _25878_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11479_));
 sky130_fd_sc_hd__mux4_1 _25879_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_271 ();
 sky130_fd_sc_hd__mux4_1 _25881_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net621),
    .S1(net625),
    .X(_11482_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_270 ();
 sky130_fd_sc_hd__mux4_1 _25883_ (.A0(_11476_),
    .A1(_11479_),
    .A2(_11480_),
    .A3(_11482_),
    .S0(net617),
    .S1(net613),
    .X(_11484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_269 ();
 sky130_fd_sc_hd__mux2i_4 _25885_ (.A0(_11475_),
    .A1(_11484_),
    .S(net610),
    .Y(_11486_));
 sky130_fd_sc_hd__mux4_1 _25886_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net619),
    .S1(net627),
    .X(_11487_));
 sky130_fd_sc_hd__mux4_1 _25887_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net619),
    .S1(net627),
    .X(_11488_));
 sky130_fd_sc_hd__mux4_1 _25888_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net619),
    .S1(net627),
    .X(_11489_));
 sky130_fd_sc_hd__mux4_1 _25889_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net619),
    .S1(net627),
    .X(_11490_));
 sky130_fd_sc_hd__mux4_4 _25890_ (.A0(_11487_),
    .A1(_11488_),
    .A2(_11489_),
    .A3(_11490_),
    .S0(net616),
    .S1(net614),
    .X(_11491_));
 sky130_fd_sc_hd__mux4_1 _25891_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net618),
    .S1(net626),
    .X(_11492_));
 sky130_fd_sc_hd__mux4_1 _25892_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net618),
    .S1(net626),
    .X(_11493_));
 sky130_fd_sc_hd__mux4_1 _25893_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net618),
    .S1(net626),
    .X(_11494_));
 sky130_fd_sc_hd__mux4_1 _25894_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net618),
    .S1(net626),
    .X(_11495_));
 sky130_fd_sc_hd__mux4_1 _25895_ (.A0(_11492_),
    .A1(_11493_),
    .A2(_11494_),
    .A3(_11495_),
    .S0(net616),
    .S1(net614),
    .X(_11496_));
 sky130_fd_sc_hd__mux2i_4 _25896_ (.A0(_11491_),
    .A1(_11496_),
    .S(net611),
    .Y(_11497_));
 sky130_fd_sc_hd__xnor2_1 _25897_ (.A(_11486_),
    .B(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__xnor2_1 _25898_ (.A(_11306_),
    .B(_11498_),
    .Y(_11779_));
 sky130_fd_sc_hd__mux4_1 _25899_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net695),
    .S1(net699),
    .X(_11499_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_268 ();
 sky130_fd_sc_hd__mux4_1 _25901_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net695),
    .S1(net699),
    .X(_11501_));
 sky130_fd_sc_hd__mux4_1 _25902_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net695),
    .S1(net699),
    .X(_11502_));
 sky130_fd_sc_hd__mux4_1 _25903_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net695),
    .S1(net699),
    .X(_11503_));
 sky130_fd_sc_hd__mux4_4 _25904_ (.A0(_11499_),
    .A1(_11501_),
    .A2(_11502_),
    .A3(_11503_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11504_));
 sky130_fd_sc_hd__mux4_1 _25905_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net693),
    .S1(net699),
    .X(_11505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_267 ();
 sky130_fd_sc_hd__mux4_1 _25907_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net693),
    .S1(net699),
    .X(_11507_));
 sky130_fd_sc_hd__mux4_1 _25908_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net693),
    .S1(net699),
    .X(_11508_));
 sky130_fd_sc_hd__mux4_1 _25909_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net693),
    .S1(net699),
    .X(_11509_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_266 ();
 sky130_fd_sc_hd__mux4_1 _25911_ (.A0(_11505_),
    .A1(_11507_),
    .A2(_11508_),
    .A3(_11509_),
    .S0(net688),
    .S1(net686),
    .X(_11511_));
 sky130_fd_sc_hd__mux2i_4 _25912_ (.A0(_11504_),
    .A1(_11511_),
    .S(net684),
    .Y(_11512_));
 sky130_fd_sc_hd__mux4_1 _25913_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net695),
    .S1(net699),
    .X(_11513_));
 sky130_fd_sc_hd__mux4_1 _25914_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net695),
    .S1(net699),
    .X(_11514_));
 sky130_fd_sc_hd__mux4_1 _25915_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net695),
    .S1(net699),
    .X(_11515_));
 sky130_fd_sc_hd__mux4_1 _25916_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net695),
    .S1(net699),
    .X(_11516_));
 sky130_fd_sc_hd__mux4_4 _25917_ (.A0(_11513_),
    .A1(_11514_),
    .A2(_11515_),
    .A3(_11516_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11517_));
 sky130_fd_sc_hd__mux4_1 _25918_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net696),
    .S1(net701),
    .X(_11518_));
 sky130_fd_sc_hd__mux4_1 _25919_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net696),
    .S1(net701),
    .X(_11519_));
 sky130_fd_sc_hd__mux4_1 _25920_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net696),
    .S1(net701),
    .X(_11520_));
 sky130_fd_sc_hd__mux4_1 _25921_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net696),
    .S1(net701),
    .X(_11521_));
 sky130_fd_sc_hd__mux4_2 _25922_ (.A0(_11518_),
    .A1(_11519_),
    .A2(_11520_),
    .A3(_11521_),
    .S0(net688),
    .S1(net686),
    .X(_11522_));
 sky130_fd_sc_hd__mux2i_4 _25923_ (.A0(_11517_),
    .A1(_11522_),
    .S(net684),
    .Y(_11523_));
 sky130_fd_sc_hd__xnor2_2 _25924_ (.A(_11512_),
    .B(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__xnor2_4 _25925_ (.A(_11234_),
    .B(_11524_),
    .Y(_11782_));
 sky130_fd_sc_hd__mux4_1 _25926_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11525_));
 sky130_fd_sc_hd__mux4_1 _25927_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11526_));
 sky130_fd_sc_hd__mux4_1 _25928_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11527_));
 sky130_fd_sc_hd__mux4_1 _25929_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11528_));
 sky130_fd_sc_hd__mux4_4 _25930_ (.A0(_11525_),
    .A1(_11526_),
    .A2(_11527_),
    .A3(_11528_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11529_));
 sky130_fd_sc_hd__mux4_1 _25931_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net623),
    .S1(net628),
    .X(_11530_));
 sky130_fd_sc_hd__mux4_1 _25932_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net623),
    .S1(net628),
    .X(_11531_));
 sky130_fd_sc_hd__mux4_1 _25933_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net623),
    .S1(net628),
    .X(_11532_));
 sky130_fd_sc_hd__mux4_1 _25934_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net623),
    .S1(net628),
    .X(_11533_));
 sky130_fd_sc_hd__mux4_1 _25935_ (.A0(_11530_),
    .A1(_11531_),
    .A2(_11532_),
    .A3(_11533_),
    .S0(net617),
    .S1(net613),
    .X(_11534_));
 sky130_fd_sc_hd__mux2i_4 _25936_ (.A0(_11529_),
    .A1(_11534_),
    .S(\count2_1[5] ),
    .Y(_11535_));
 sky130_fd_sc_hd__mux4_1 _25937_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11536_));
 sky130_fd_sc_hd__mux4_1 _25938_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11537_));
 sky130_fd_sc_hd__mux4_1 _25939_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11538_));
 sky130_fd_sc_hd__mux4_1 _25940_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11539_));
 sky130_fd_sc_hd__mux4_2 _25941_ (.A0(_11536_),
    .A1(_11537_),
    .A2(_11538_),
    .A3(_11539_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11540_));
 sky130_fd_sc_hd__mux4_1 _25942_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11541_));
 sky130_fd_sc_hd__mux4_1 _25943_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11542_));
 sky130_fd_sc_hd__mux4_1 _25944_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11543_));
 sky130_fd_sc_hd__mux4_1 _25945_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_11544_));
 sky130_fd_sc_hd__mux4_1 _25946_ (.A0(_11541_),
    .A1(_11542_),
    .A2(_11543_),
    .A3(_11544_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11545_));
 sky130_fd_sc_hd__mux2i_4 _25947_ (.A0(_11540_),
    .A1(_11545_),
    .S(\count2_1[5] ),
    .Y(_11546_));
 sky130_fd_sc_hd__xnor2_1 _25948_ (.A(_11535_),
    .B(_11546_),
    .Y(_11547_));
 sky130_fd_sc_hd__xnor2_1 _25949_ (.A(_11430_),
    .B(_11547_),
    .Y(_11787_));
 sky130_fd_sc_hd__mux4_1 _25950_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net690),
    .S1(net697),
    .X(_11548_));
 sky130_fd_sc_hd__mux4_1 _25951_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net690),
    .S1(\count15_1[1] ),
    .X(_11549_));
 sky130_fd_sc_hd__mux4_1 _25952_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net690),
    .S1(net697),
    .X(_11550_));
 sky130_fd_sc_hd__mux4_1 _25953_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net690),
    .S1(net697),
    .X(_11551_));
 sky130_fd_sc_hd__mux4_4 _25954_ (.A0(_11548_),
    .A1(_11549_),
    .A2(_11550_),
    .A3(_11551_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11552_));
 sky130_fd_sc_hd__mux4_1 _25955_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net692),
    .S1(net699),
    .X(_11553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_265 ();
 sky130_fd_sc_hd__mux4_1 _25957_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net691),
    .S1(net699),
    .X(_11555_));
 sky130_fd_sc_hd__mux4_1 _25958_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net691),
    .S1(net699),
    .X(_11556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_263 ();
 sky130_fd_sc_hd__mux4_1 _25961_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net692),
    .S1(net699),
    .X(_11559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_262 ();
 sky130_fd_sc_hd__mux4_2 _25963_ (.A0(_11553_),
    .A1(_11555_),
    .A2(_11556_),
    .A3(_11559_),
    .S0(net687),
    .S1(net685),
    .X(_11561_));
 sky130_fd_sc_hd__mux2i_4 _25964_ (.A0(_11552_),
    .A1(_11561_),
    .S(net683),
    .Y(_11562_));
 sky130_fd_sc_hd__mux4_1 _25965_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net694),
    .S1(net700),
    .X(_11563_));
 sky130_fd_sc_hd__mux4_1 _25966_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net691),
    .S1(net697),
    .X(_11564_));
 sky130_fd_sc_hd__mux4_1 _25967_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net694),
    .S1(net700),
    .X(_11565_));
 sky130_fd_sc_hd__mux4_1 _25968_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net694),
    .S1(net700),
    .X(_11566_));
 sky130_fd_sc_hd__mux4_4 _25969_ (.A0(_11563_),
    .A1(_11564_),
    .A2(_11565_),
    .A3(_11566_),
    .S0(net688),
    .S1(net686),
    .X(_11567_));
 sky130_fd_sc_hd__mux4_1 _25970_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net696),
    .S1(net698),
    .X(_11568_));
 sky130_fd_sc_hd__mux4_1 _25971_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net696),
    .S1(net698),
    .X(_11569_));
 sky130_fd_sc_hd__mux4_1 _25972_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net696),
    .S1(net698),
    .X(_11570_));
 sky130_fd_sc_hd__mux4_1 _25973_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net696),
    .S1(net698),
    .X(_11571_));
 sky130_fd_sc_hd__mux4_1 _25974_ (.A0(_11568_),
    .A1(_11569_),
    .A2(_11570_),
    .A3(_11571_),
    .S0(net688),
    .S1(net686),
    .X(_11572_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_261 ();
 sky130_fd_sc_hd__mux2i_4 _25976_ (.A0(_11567_),
    .A1(_11572_),
    .S(net684),
    .Y(_11574_));
 sky130_fd_sc_hd__xnor2_1 _25977_ (.A(_11562_),
    .B(_11574_),
    .Y(_11575_));
 sky130_fd_sc_hd__xnor2_2 _25978_ (.A(_11271_),
    .B(_11575_),
    .Y(_11790_));
 sky130_fd_sc_hd__mux4_1 _25979_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11576_));
 sky130_fd_sc_hd__mux4_1 _25980_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11577_));
 sky130_fd_sc_hd__mux4_1 _25981_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11578_));
 sky130_fd_sc_hd__mux4_1 _25982_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11579_));
 sky130_fd_sc_hd__mux4_4 _25983_ (.A0(_11576_),
    .A1(_11577_),
    .A2(_11578_),
    .A3(_11579_),
    .S0(net616),
    .S1(\count2_1[4] ),
    .X(_11580_));
 sky130_fd_sc_hd__mux4_1 _25984_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11581_));
 sky130_fd_sc_hd__mux4_1 _25985_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11582_));
 sky130_fd_sc_hd__mux4_1 _25986_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11583_));
 sky130_fd_sc_hd__mux4_1 _25987_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net620),
    .S1(net624),
    .X(_11584_));
 sky130_fd_sc_hd__mux4_1 _25988_ (.A0(_11581_),
    .A1(_11582_),
    .A2(_11583_),
    .A3(_11584_),
    .S0(net616),
    .S1(\count2_1[4] ),
    .X(_11585_));
 sky130_fd_sc_hd__mux2i_4 _25989_ (.A0(_11580_),
    .A1(_11585_),
    .S(\count2_1[5] ),
    .Y(_11586_));
 sky130_fd_sc_hd__mux4_1 _25990_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11587_));
 sky130_fd_sc_hd__mux4_1 _25991_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11588_));
 sky130_fd_sc_hd__mux4_1 _25992_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11589_));
 sky130_fd_sc_hd__mux4_1 _25993_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11590_));
 sky130_fd_sc_hd__mux4_4 _25994_ (.A0(_11587_),
    .A1(_11588_),
    .A2(_11589_),
    .A3(_11590_),
    .S0(net617),
    .S1(net613),
    .X(_11591_));
 sky130_fd_sc_hd__mux4_1 _25995_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11592_));
 sky130_fd_sc_hd__mux4_1 _25996_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11593_));
 sky130_fd_sc_hd__mux4_1 _25997_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11594_));
 sky130_fd_sc_hd__mux4_1 _25998_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net622),
    .S1(net628),
    .X(_11595_));
 sky130_fd_sc_hd__mux4_1 _25999_ (.A0(_11592_),
    .A1(_11593_),
    .A2(_11594_),
    .A3(_11595_),
    .S0(net617),
    .S1(net613),
    .X(_11596_));
 sky130_fd_sc_hd__mux2i_4 _26000_ (.A0(_11591_),
    .A1(_11596_),
    .S(net611),
    .Y(_11597_));
 sky130_fd_sc_hd__xnor2_1 _26001_ (.A(_11586_),
    .B(_11597_),
    .Y(_11598_));
 sky130_fd_sc_hd__xnor2_1 _26002_ (.A(_11497_),
    .B(_11598_),
    .Y(_11795_));
 sky130_fd_sc_hd__mux4_1 _26003_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net690),
    .S1(net697),
    .X(_11599_));
 sky130_fd_sc_hd__mux4_1 _26004_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net690),
    .S1(net697),
    .X(_11600_));
 sky130_fd_sc_hd__mux4_1 _26005_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net690),
    .S1(net697),
    .X(_11601_));
 sky130_fd_sc_hd__mux4_1 _26006_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net690),
    .S1(net697),
    .X(_11602_));
 sky130_fd_sc_hd__mux4_4 _26007_ (.A0(_11599_),
    .A1(_11600_),
    .A2(_11601_),
    .A3(_11602_),
    .S0(net687),
    .S1(net685),
    .X(_11603_));
 sky130_fd_sc_hd__mux4_1 _26008_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net691),
    .S1(net697),
    .X(_11604_));
 sky130_fd_sc_hd__mux4_1 _26009_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net691),
    .S1(net697),
    .X(_11605_));
 sky130_fd_sc_hd__mux4_1 _26010_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net691),
    .S1(net697),
    .X(_11606_));
 sky130_fd_sc_hd__mux4_1 _26011_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net691),
    .S1(net697),
    .X(_11607_));
 sky130_fd_sc_hd__mux4_1 _26012_ (.A0(_11604_),
    .A1(_11605_),
    .A2(_11606_),
    .A3(_11607_),
    .S0(net687),
    .S1(net685),
    .X(_11608_));
 sky130_fd_sc_hd__mux2i_4 _26013_ (.A0(_11603_),
    .A1(_11608_),
    .S(net683),
    .Y(_11609_));
 sky130_fd_sc_hd__mux4_1 _26014_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net695),
    .S1(net699),
    .X(_11610_));
 sky130_fd_sc_hd__mux4_1 _26015_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net695),
    .S1(net699),
    .X(_11611_));
 sky130_fd_sc_hd__mux4_1 _26016_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net695),
    .S1(net699),
    .X(_11612_));
 sky130_fd_sc_hd__mux4_1 _26017_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net695),
    .S1(net699),
    .X(_11613_));
 sky130_fd_sc_hd__mux4_4 _26018_ (.A0(_11610_),
    .A1(_11611_),
    .A2(_11612_),
    .A3(_11613_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11614_));
 sky130_fd_sc_hd__mux4_1 _26019_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net695),
    .S1(net701),
    .X(_11615_));
 sky130_fd_sc_hd__mux4_1 _26020_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net695),
    .S1(net701),
    .X(_11616_));
 sky130_fd_sc_hd__mux4_1 _26021_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net695),
    .S1(net701),
    .X(_11617_));
 sky130_fd_sc_hd__mux4_1 _26022_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net695),
    .S1(net701),
    .X(_11618_));
 sky130_fd_sc_hd__mux4_1 _26023_ (.A0(_11615_),
    .A1(_11616_),
    .A2(_11617_),
    .A3(_11618_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_11619_));
 sky130_fd_sc_hd__mux2i_4 _26024_ (.A0(_11614_),
    .A1(_11619_),
    .S(net684),
    .Y(_11620_));
 sky130_fd_sc_hd__xnor2_2 _26025_ (.A(_11609_),
    .B(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__xnor2_4 _26026_ (.A(_11385_),
    .B(_11621_),
    .Y(_11798_));
 sky130_fd_sc_hd__mux4_1 _26027_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11622_));
 sky130_fd_sc_hd__mux4_1 _26028_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11623_));
 sky130_fd_sc_hd__mux4_1 _26029_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11624_));
 sky130_fd_sc_hd__mux4_1 _26030_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11625_));
 sky130_fd_sc_hd__mux4_4 _26031_ (.A0(_11622_),
    .A1(_11623_),
    .A2(_11624_),
    .A3(_11625_),
    .S0(net615),
    .S1(net612),
    .X(_11626_));
 sky130_fd_sc_hd__mux4_1 _26032_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11627_));
 sky130_fd_sc_hd__mux4_1 _26033_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11628_));
 sky130_fd_sc_hd__mux4_1 _26034_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11629_));
 sky130_fd_sc_hd__mux4_1 _26035_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net619),
    .S1(net627),
    .X(_11630_));
 sky130_fd_sc_hd__mux4_1 _26036_ (.A0(_11627_),
    .A1(_11628_),
    .A2(_11629_),
    .A3(_11630_),
    .S0(net615),
    .S1(net612),
    .X(_11631_));
 sky130_fd_sc_hd__mux2i_4 _26037_ (.A0(_11626_),
    .A1(_11631_),
    .S(net610),
    .Y(_11632_));
 sky130_fd_sc_hd__mux4_1 _26038_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net618),
    .S1(net626),
    .X(_11633_));
 sky130_fd_sc_hd__mux4_1 _26039_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net618),
    .S1(net626),
    .X(_11634_));
 sky130_fd_sc_hd__mux4_1 _26040_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net618),
    .S1(net626),
    .X(_11635_));
 sky130_fd_sc_hd__mux4_1 _26041_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net618),
    .S1(net626),
    .X(_11636_));
 sky130_fd_sc_hd__mux4_4 _26042_ (.A0(_11633_),
    .A1(_11634_),
    .A2(_11635_),
    .A3(_11636_),
    .S0(net615),
    .S1(net612),
    .X(_11637_));
 sky130_fd_sc_hd__mux4_1 _26043_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net623),
    .S1(net625),
    .X(_11638_));
 sky130_fd_sc_hd__mux4_1 _26044_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net623),
    .S1(net625),
    .X(_11639_));
 sky130_fd_sc_hd__mux4_1 _26045_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net623),
    .S1(net625),
    .X(_11640_));
 sky130_fd_sc_hd__mux4_1 _26046_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net623),
    .S1(net625),
    .X(_11641_));
 sky130_fd_sc_hd__mux4_1 _26047_ (.A0(_11638_),
    .A1(_11639_),
    .A2(_11640_),
    .A3(_11641_),
    .S0(net617),
    .S1(net613),
    .X(_11642_));
 sky130_fd_sc_hd__mux2i_4 _26048_ (.A0(_11637_),
    .A1(_11642_),
    .S(net611),
    .Y(_11643_));
 sky130_fd_sc_hd__xnor2_1 _26049_ (.A(_11632_),
    .B(_11643_),
    .Y(_11644_));
 sky130_fd_sc_hd__xnor2_1 _26050_ (.A(_11535_),
    .B(_11644_),
    .Y(_11803_));
 sky130_fd_sc_hd__mux4_1 _26051_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net690),
    .S1(net697),
    .X(_11645_));
 sky130_fd_sc_hd__mux4_1 _26052_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net690),
    .S1(net697),
    .X(_11646_));
 sky130_fd_sc_hd__mux4_1 _26053_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net690),
    .S1(net697),
    .X(_11647_));
 sky130_fd_sc_hd__mux4_1 _26054_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net690),
    .S1(net697),
    .X(_11648_));
 sky130_fd_sc_hd__mux4_2 _26055_ (.A0(_11645_),
    .A1(_11646_),
    .A2(_11647_),
    .A3(_11648_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11649_));
 sky130_fd_sc_hd__mux4_1 _26056_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net692),
    .S1(net700),
    .X(_11650_));
 sky130_fd_sc_hd__mux4_1 _26057_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net692),
    .S1(net700),
    .X(_11651_));
 sky130_fd_sc_hd__mux4_1 _26058_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net692),
    .S1(net700),
    .X(_11652_));
 sky130_fd_sc_hd__mux4_1 _26059_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net692),
    .S1(net700),
    .X(_11653_));
 sky130_fd_sc_hd__mux4_1 _26060_ (.A0(_11650_),
    .A1(_11651_),
    .A2(_11652_),
    .A3(_11653_),
    .S0(net687),
    .S1(net685),
    .X(_11654_));
 sky130_fd_sc_hd__mux2i_4 _26061_ (.A0(_11649_),
    .A1(_11654_),
    .S(net683),
    .Y(_11655_));
 sky130_fd_sc_hd__mux4_1 _26062_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net691),
    .S1(net697),
    .X(_11656_));
 sky130_fd_sc_hd__mux4_1 _26063_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net691),
    .S1(net697),
    .X(_11657_));
 sky130_fd_sc_hd__mux4_1 _26064_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net691),
    .S1(net697),
    .X(_11658_));
 sky130_fd_sc_hd__mux4_1 _26065_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net691),
    .S1(net697),
    .X(_11659_));
 sky130_fd_sc_hd__mux4_4 _26066_ (.A0(_11656_),
    .A1(_11657_),
    .A2(_11658_),
    .A3(_11659_),
    .S0(net687),
    .S1(net685),
    .X(_11660_));
 sky130_fd_sc_hd__mux4_1 _26067_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net691),
    .S1(net700),
    .X(_11661_));
 sky130_fd_sc_hd__mux4_1 _26068_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net691),
    .S1(net700),
    .X(_11662_));
 sky130_fd_sc_hd__mux4_1 _26069_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net691),
    .S1(net700),
    .X(_11663_));
 sky130_fd_sc_hd__mux4_1 _26070_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net691),
    .S1(net700),
    .X(_11664_));
 sky130_fd_sc_hd__mux4_1 _26071_ (.A0(_11661_),
    .A1(_11662_),
    .A2(_11663_),
    .A3(_11664_),
    .S0(net687),
    .S1(net685),
    .X(_11665_));
 sky130_fd_sc_hd__mux2i_4 _26072_ (.A0(_11660_),
    .A1(_11665_),
    .S(net683),
    .Y(_11666_));
 sky130_fd_sc_hd__xnor2_1 _26073_ (.A(_11655_),
    .B(_11666_),
    .Y(_11667_));
 sky130_fd_sc_hd__xnor2_2 _26074_ (.A(_11468_),
    .B(_11667_),
    .Y(_11806_));
 sky130_fd_sc_hd__mux4_1 _26075_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net619),
    .S1(net627),
    .X(_11668_));
 sky130_fd_sc_hd__mux4_1 _26076_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net619),
    .S1(net627),
    .X(_11669_));
 sky130_fd_sc_hd__mux4_1 _26077_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net619),
    .S1(net627),
    .X(_11670_));
 sky130_fd_sc_hd__mux4_1 _26078_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net619),
    .S1(net627),
    .X(_11671_));
 sky130_fd_sc_hd__mux4_4 _26079_ (.A0(_11668_),
    .A1(_11669_),
    .A2(_11670_),
    .A3(_11671_),
    .S0(net615),
    .S1(net612),
    .X(_11672_));
 sky130_fd_sc_hd__mux4_1 _26080_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net623),
    .S1(net628),
    .X(_11673_));
 sky130_fd_sc_hd__mux4_1 _26081_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net623),
    .S1(net628),
    .X(_11674_));
 sky130_fd_sc_hd__mux4_1 _26082_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net623),
    .S1(net628),
    .X(_11675_));
 sky130_fd_sc_hd__mux4_1 _26083_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net623),
    .S1(net628),
    .X(_11676_));
 sky130_fd_sc_hd__mux4_1 _26084_ (.A0(_11673_),
    .A1(_11674_),
    .A2(_11675_),
    .A3(_11676_),
    .S0(net617),
    .S1(net613),
    .X(_11677_));
 sky130_fd_sc_hd__mux2i_4 _26085_ (.A0(_11672_),
    .A1(_11677_),
    .S(net611),
    .Y(_11678_));
 sky130_fd_sc_hd__mux4_1 _26086_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net621),
    .S1(net625),
    .X(_11679_));
 sky130_fd_sc_hd__mux4_1 _26087_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net621),
    .S1(net625),
    .X(_11680_));
 sky130_fd_sc_hd__mux4_1 _26088_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net621),
    .S1(net625),
    .X(_11681_));
 sky130_fd_sc_hd__mux4_1 _26089_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net621),
    .S1(net625),
    .X(_11682_));
 sky130_fd_sc_hd__mux4_4 _26090_ (.A0(_11679_),
    .A1(_11680_),
    .A2(_11681_),
    .A3(_11682_),
    .S0(net617),
    .S1(net613),
    .X(_11683_));
 sky130_fd_sc_hd__mux4_1 _26091_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net623),
    .S1(net625),
    .X(_11684_));
 sky130_fd_sc_hd__mux4_1 _26092_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net623),
    .S1(net625),
    .X(_11685_));
 sky130_fd_sc_hd__mux4_1 _26093_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net623),
    .S1(net625),
    .X(_11686_));
 sky130_fd_sc_hd__mux4_1 _26094_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net623),
    .S1(net625),
    .X(_11687_));
 sky130_fd_sc_hd__mux4_1 _26095_ (.A0(_11684_),
    .A1(_11685_),
    .A2(_11686_),
    .A3(_11687_),
    .S0(net615),
    .S1(net612),
    .X(_11688_));
 sky130_fd_sc_hd__mux2i_4 _26096_ (.A0(_11683_),
    .A1(_11688_),
    .S(net610),
    .Y(_11689_));
 sky130_fd_sc_hd__xnor2_1 _26097_ (.A(_11678_),
    .B(_11689_),
    .Y(_11690_));
 sky130_fd_sc_hd__xnor2_1 _26098_ (.A(_11597_),
    .B(_11690_),
    .Y(_11811_));
 sky130_fd_sc_hd__mux4_1 _26099_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net691),
    .S1(net697),
    .X(_11691_));
 sky130_fd_sc_hd__mux4_1 _26100_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net691),
    .S1(net697),
    .X(_11692_));
 sky130_fd_sc_hd__mux4_1 _26101_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net691),
    .S1(net697),
    .X(_11693_));
 sky130_fd_sc_hd__mux4_1 _26102_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net691),
    .S1(net697),
    .X(_11694_));
 sky130_fd_sc_hd__mux4_4 _26103_ (.A0(_11691_),
    .A1(_11692_),
    .A2(_11693_),
    .A3(_11694_),
    .S0(net688),
    .S1(net686),
    .X(_11695_));
 sky130_fd_sc_hd__mux4_1 _26104_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net696),
    .S1(net700),
    .X(_11696_));
 sky130_fd_sc_hd__mux4_1 _26105_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net696),
    .S1(net700),
    .X(_11697_));
 sky130_fd_sc_hd__mux4_1 _26106_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net696),
    .S1(net700),
    .X(_11698_));
 sky130_fd_sc_hd__mux4_1 _26107_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net696),
    .S1(net700),
    .X(_11699_));
 sky130_fd_sc_hd__mux4_1 _26108_ (.A0(_11696_),
    .A1(_11697_),
    .A2(_11698_),
    .A3(_11699_),
    .S0(net688),
    .S1(net686),
    .X(_11700_));
 sky130_fd_sc_hd__mux2i_4 _26109_ (.A0(_11695_),
    .A1(_11700_),
    .S(net683),
    .Y(_11701_));
 sky130_fd_sc_hd__mux4_1 _26110_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net690),
    .S1(net697),
    .X(_11702_));
 sky130_fd_sc_hd__mux4_1 _26111_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net690),
    .S1(\count15_1[1] ),
    .X(_11703_));
 sky130_fd_sc_hd__mux4_1 _26112_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net690),
    .S1(net697),
    .X(_11704_));
 sky130_fd_sc_hd__mux4_1 _26113_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net690),
    .S1(net697),
    .X(_11705_));
 sky130_fd_sc_hd__mux4_2 _26114_ (.A0(_11702_),
    .A1(_11703_),
    .A2(_11704_),
    .A3(_11705_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11706_));
 sky130_fd_sc_hd__mux4_1 _26115_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net692),
    .S1(net700),
    .X(_11707_));
 sky130_fd_sc_hd__mux4_1 _26116_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net692),
    .S1(net700),
    .X(_11708_));
 sky130_fd_sc_hd__mux4_1 _26117_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net692),
    .S1(net700),
    .X(_11709_));
 sky130_fd_sc_hd__mux4_1 _26118_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net692),
    .S1(net700),
    .X(_11710_));
 sky130_fd_sc_hd__mux4_1 _26119_ (.A0(_11707_),
    .A1(_11708_),
    .A2(_11709_),
    .A3(_11710_),
    .S0(net687),
    .S1(net685),
    .X(_11711_));
 sky130_fd_sc_hd__mux2i_4 _26120_ (.A0(_11706_),
    .A1(_11711_),
    .S(net683),
    .Y(_11712_));
 sky130_fd_sc_hd__xnor2_1 _26121_ (.A(_11701_),
    .B(_11712_),
    .Y(_11713_));
 sky130_fd_sc_hd__xnor2_2 _26122_ (.A(_11523_),
    .B(_11713_),
    .Y(_11814_));
 sky130_fd_sc_hd__mux4_1 _26123_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11714_));
 sky130_fd_sc_hd__mux4_1 _26124_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11715_));
 sky130_fd_sc_hd__mux4_1 _26125_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11716_));
 sky130_fd_sc_hd__mux4_1 _26126_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11717_));
 sky130_fd_sc_hd__mux4_4 _26127_ (.A0(_11714_),
    .A1(_11715_),
    .A2(_11716_),
    .A3(_11717_),
    .S0(net617),
    .S1(net613),
    .X(_11718_));
 sky130_fd_sc_hd__mux4_1 _26128_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11719_));
 sky130_fd_sc_hd__mux4_1 _26129_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11720_));
 sky130_fd_sc_hd__mux4_1 _26130_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11721_));
 sky130_fd_sc_hd__mux4_1 _26131_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net622),
    .S1(net628),
    .X(_11722_));
 sky130_fd_sc_hd__mux4_1 _26132_ (.A0(_11719_),
    .A1(_11720_),
    .A2(_11721_),
    .A3(_11722_),
    .S0(net617),
    .S1(net613),
    .X(_11723_));
 sky130_fd_sc_hd__mux2i_4 _26133_ (.A0(_11718_),
    .A1(_11723_),
    .S(net611),
    .Y(_11724_));
 sky130_fd_sc_hd__xnor2_1 _26134_ (.A(_11643_),
    .B(_11724_),
    .Y(_11725_));
 sky130_fd_sc_hd__xnor2_1 _26135_ (.A(_11349_),
    .B(_11725_),
    .Y(_11819_));
 sky130_fd_sc_hd__mux4_1 _26136_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net691),
    .S1(net697),
    .X(_11726_));
 sky130_fd_sc_hd__mux4_1 _26137_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net691),
    .S1(net697),
    .X(_11727_));
 sky130_fd_sc_hd__mux4_1 _26138_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net691),
    .S1(net697),
    .X(_11728_));
 sky130_fd_sc_hd__mux4_1 _26139_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net691),
    .S1(net697),
    .X(_11729_));
 sky130_fd_sc_hd__mux4_4 _26140_ (.A0(_11726_),
    .A1(_11727_),
    .A2(_11728_),
    .A3(_11729_),
    .S0(net688),
    .S1(net686),
    .X(_11730_));
 sky130_fd_sc_hd__mux4_1 _26141_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net696),
    .S1(net700),
    .X(_11731_));
 sky130_fd_sc_hd__mux4_1 _26142_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net696),
    .S1(net700),
    .X(_11732_));
 sky130_fd_sc_hd__mux4_1 _26143_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net696),
    .S1(net700),
    .X(_11733_));
 sky130_fd_sc_hd__mux4_1 _26144_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net696),
    .S1(net700),
    .X(_11734_));
 sky130_fd_sc_hd__mux4_1 _26145_ (.A0(_11731_),
    .A1(_11732_),
    .A2(_11733_),
    .A3(_11734_),
    .S0(net687),
    .S1(net686),
    .X(_11735_));
 sky130_fd_sc_hd__mux2i_4 _26146_ (.A0(_11730_),
    .A1(_11735_),
    .S(net683),
    .Y(_11736_));
 sky130_fd_sc_hd__mux4_1 _26147_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net690),
    .S1(net697),
    .X(_11737_));
 sky130_fd_sc_hd__mux4_1 _26148_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net690),
    .S1(\count15_1[1] ),
    .X(_11738_));
 sky130_fd_sc_hd__mux4_1 _26149_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net690),
    .S1(net697),
    .X(_11739_));
 sky130_fd_sc_hd__mux4_1 _26150_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net690),
    .S1(net697),
    .X(_11740_));
 sky130_fd_sc_hd__mux4_4 _26151_ (.A0(_11737_),
    .A1(_11738_),
    .A2(_11739_),
    .A3(_11740_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_11741_));
 sky130_fd_sc_hd__mux4_1 _26152_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net692),
    .S1(net700),
    .X(_11742_));
 sky130_fd_sc_hd__mux4_1 _26153_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net692),
    .S1(net700),
    .X(_11743_));
 sky130_fd_sc_hd__mux4_1 _26154_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net692),
    .S1(net700),
    .X(_11744_));
 sky130_fd_sc_hd__mux4_1 _26155_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net692),
    .S1(net700),
    .X(_11745_));
 sky130_fd_sc_hd__mux4_1 _26156_ (.A0(_11742_),
    .A1(_11743_),
    .A2(_11744_),
    .A3(_11745_),
    .S0(net687),
    .S1(net685),
    .X(_02570_));
 sky130_fd_sc_hd__mux2i_4 _26157_ (.A0(_11741_),
    .A1(_02570_),
    .S(net683),
    .Y(_02571_));
 sky130_fd_sc_hd__xnor2_1 _26158_ (.A(_11736_),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__xnor2_2 _26159_ (.A(_11562_),
    .B(_02572_),
    .Y(_11822_));
 sky130_fd_sc_hd__mux4_1 _26160_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02573_));
 sky130_fd_sc_hd__mux4_1 _26161_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02574_));
 sky130_fd_sc_hd__mux4_1 _26162_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02575_));
 sky130_fd_sc_hd__mux4_1 _26163_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02576_));
 sky130_fd_sc_hd__mux4_4 _26164_ (.A0(_02573_),
    .A1(_02574_),
    .A2(_02575_),
    .A3(_02576_),
    .S0(net617),
    .S1(net613),
    .X(_02577_));
 sky130_fd_sc_hd__mux4_1 _26165_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02578_));
 sky130_fd_sc_hd__mux4_1 _26166_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02579_));
 sky130_fd_sc_hd__mux4_1 _26167_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02580_));
 sky130_fd_sc_hd__mux4_1 _26168_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net622),
    .S1(net628),
    .X(_02581_));
 sky130_fd_sc_hd__mux4_1 _26169_ (.A0(_02578_),
    .A1(_02579_),
    .A2(_02580_),
    .A3(_02581_),
    .S0(net617),
    .S1(net613),
    .X(_02582_));
 sky130_fd_sc_hd__mux2i_4 _26170_ (.A0(_02577_),
    .A1(_02582_),
    .S(net611),
    .Y(_02583_));
 sky130_fd_sc_hd__xnor2_1 _26171_ (.A(_11678_),
    .B(_02583_),
    .Y(_02584_));
 sky130_fd_sc_hd__xnor2_1 _26172_ (.A(_11397_),
    .B(_02584_),
    .Y(_11827_));
 sky130_fd_sc_hd__mux4_1 _26173_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net690),
    .S1(net697),
    .X(_02585_));
 sky130_fd_sc_hd__mux4_1 _26174_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net690),
    .S1(net697),
    .X(_02586_));
 sky130_fd_sc_hd__mux4_1 _26175_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net690),
    .S1(net697),
    .X(_02587_));
 sky130_fd_sc_hd__mux4_1 _26176_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net690),
    .S1(net697),
    .X(_02588_));
 sky130_fd_sc_hd__mux4_2 _26177_ (.A0(_02585_),
    .A1(_02586_),
    .A2(_02587_),
    .A3(_02588_),
    .S0(net687),
    .S1(net685),
    .X(_02589_));
 sky130_fd_sc_hd__mux4_1 _26178_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net692),
    .S1(net697),
    .X(_02590_));
 sky130_fd_sc_hd__mux4_1 _26179_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net692),
    .S1(net697),
    .X(_02591_));
 sky130_fd_sc_hd__mux4_1 _26180_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net692),
    .S1(net697),
    .X(_02592_));
 sky130_fd_sc_hd__mux4_1 _26181_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net692),
    .S1(net697),
    .X(_02593_));
 sky130_fd_sc_hd__mux4_1 _26182_ (.A0(_02590_),
    .A1(_02591_),
    .A2(_02592_),
    .A3(_02593_),
    .S0(net687),
    .S1(net685),
    .X(_02594_));
 sky130_fd_sc_hd__mux2i_4 _26183_ (.A0(_02589_),
    .A1(_02594_),
    .S(net683),
    .Y(_02595_));
 sky130_fd_sc_hd__mux4_1 _26184_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net694),
    .S1(net700),
    .X(_02596_));
 sky130_fd_sc_hd__mux4_1 _26185_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net694),
    .S1(net700),
    .X(_02597_));
 sky130_fd_sc_hd__mux4_1 _26186_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net694),
    .S1(net700),
    .X(_02598_));
 sky130_fd_sc_hd__mux4_1 _26187_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net694),
    .S1(net700),
    .X(_02599_));
 sky130_fd_sc_hd__mux4_4 _26188_ (.A0(_02596_),
    .A1(_02597_),
    .A2(_02598_),
    .A3(_02599_),
    .S0(net688),
    .S1(net686),
    .X(_02600_));
 sky130_fd_sc_hd__mux4_1 _26189_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net694),
    .S1(net698),
    .X(_02601_));
 sky130_fd_sc_hd__mux4_1 _26190_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net694),
    .S1(net698),
    .X(_02602_));
 sky130_fd_sc_hd__mux4_1 _26191_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net694),
    .S1(net698),
    .X(_02603_));
 sky130_fd_sc_hd__mux4_1 _26192_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net694),
    .S1(net698),
    .X(_02604_));
 sky130_fd_sc_hd__mux4_1 _26193_ (.A0(_02601_),
    .A1(_02602_),
    .A2(_02603_),
    .A3(_02604_),
    .S0(net688),
    .S1(net686),
    .X(_02605_));
 sky130_fd_sc_hd__mux2i_4 _26194_ (.A0(_02600_),
    .A1(_02605_),
    .S(net684),
    .Y(_02606_));
 sky130_fd_sc_hd__xnor2_1 _26195_ (.A(_02595_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__xnor2_2 _26196_ (.A(_11620_),
    .B(_02607_),
    .Y(_11830_));
 sky130_fd_sc_hd__mux4_1 _26197_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net618),
    .S1(net626),
    .X(_02608_));
 sky130_fd_sc_hd__mux4_1 _26198_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net618),
    .S1(net626),
    .X(_02609_));
 sky130_fd_sc_hd__mux4_1 _26199_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net618),
    .S1(net626),
    .X(_02610_));
 sky130_fd_sc_hd__mux4_1 _26200_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net618),
    .S1(net626),
    .X(_02611_));
 sky130_fd_sc_hd__mux4_4 _26201_ (.A0(_02608_),
    .A1(_02609_),
    .A2(_02610_),
    .A3(_02611_),
    .S0(net616),
    .S1(net614),
    .X(_02612_));
 sky130_fd_sc_hd__mux4_1 _26202_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net619),
    .S1(net627),
    .X(_02613_));
 sky130_fd_sc_hd__mux4_1 _26203_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net619),
    .S1(net627),
    .X(_02614_));
 sky130_fd_sc_hd__mux4_1 _26204_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net619),
    .S1(net627),
    .X(_02615_));
 sky130_fd_sc_hd__mux4_1 _26205_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net619),
    .S1(net627),
    .X(_02616_));
 sky130_fd_sc_hd__mux4_1 _26206_ (.A0(_02613_),
    .A1(_02614_),
    .A2(_02615_),
    .A3(_02616_),
    .S0(net615),
    .S1(net612),
    .X(_02617_));
 sky130_fd_sc_hd__mux2i_4 _26207_ (.A0(_02612_),
    .A1(_02617_),
    .S(net611),
    .Y(_02618_));
 sky130_fd_sc_hd__xnor2_1 _26208_ (.A(_11724_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__xnor2_1 _26209_ (.A(_11306_),
    .B(_02619_),
    .Y(_11835_));
 sky130_fd_sc_hd__mux4_1 _26210_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net695),
    .S1(net699),
    .X(_02620_));
 sky130_fd_sc_hd__mux4_1 _26211_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net695),
    .S1(net699),
    .X(_02621_));
 sky130_fd_sc_hd__mux4_1 _26212_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net695),
    .S1(net699),
    .X(_02622_));
 sky130_fd_sc_hd__mux4_1 _26213_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net695),
    .S1(net699),
    .X(_02623_));
 sky130_fd_sc_hd__mux4_2 _26214_ (.A0(_02620_),
    .A1(_02621_),
    .A2(_02622_),
    .A3(_02623_),
    .S0(net689),
    .S1(\count15_1[4] ),
    .X(_02624_));
 sky130_fd_sc_hd__mux4_1 _26215_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net693),
    .S1(net699),
    .X(_02625_));
 sky130_fd_sc_hd__mux4_1 _26216_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net693),
    .S1(net698),
    .X(_02626_));
 sky130_fd_sc_hd__mux4_1 _26217_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net693),
    .S1(net698),
    .X(_02627_));
 sky130_fd_sc_hd__mux4_1 _26218_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net693),
    .S1(net698),
    .X(_02628_));
 sky130_fd_sc_hd__mux4_1 _26219_ (.A0(_02625_),
    .A1(_02626_),
    .A2(_02627_),
    .A3(_02628_),
    .S0(net688),
    .S1(net686),
    .X(_02629_));
 sky130_fd_sc_hd__mux2i_4 _26220_ (.A0(_02624_),
    .A1(_02629_),
    .S(net684),
    .Y(_02630_));
 sky130_fd_sc_hd__xnor2_1 _26221_ (.A(_11655_),
    .B(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__xnor2_2 _26222_ (.A(_11208_),
    .B(_02631_),
    .Y(_11838_));
 sky130_fd_sc_hd__mux4_1 _26223_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02632_));
 sky130_fd_sc_hd__mux4_1 _26224_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02633_));
 sky130_fd_sc_hd__mux4_1 _26225_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02634_));
 sky130_fd_sc_hd__mux4_1 _26226_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02635_));
 sky130_fd_sc_hd__mux4_4 _26227_ (.A0(_02632_),
    .A1(_02633_),
    .A2(_02634_),
    .A3(_02635_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02636_));
 sky130_fd_sc_hd__mux4_1 _26228_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net620),
    .S1(net624),
    .X(_02637_));
 sky130_fd_sc_hd__mux4_1 _26229_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net620),
    .S1(net624),
    .X(_02638_));
 sky130_fd_sc_hd__mux4_1 _26230_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net620),
    .S1(net624),
    .X(_02639_));
 sky130_fd_sc_hd__mux4_1 _26231_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net620),
    .S1(net624),
    .X(_02640_));
 sky130_fd_sc_hd__mux4_1 _26232_ (.A0(_02637_),
    .A1(_02638_),
    .A2(_02639_),
    .A3(_02640_),
    .S0(net616),
    .S1(\count2_1[4] ),
    .X(_02641_));
 sky130_fd_sc_hd__mux2i_4 _26233_ (.A0(_02636_),
    .A1(_02641_),
    .S(\count2_1[5] ),
    .Y(_02642_));
 sky130_fd_sc_hd__xnor2_1 _26234_ (.A(_02583_),
    .B(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__xnor2_1 _26235_ (.A(_11430_),
    .B(_02643_),
    .Y(_11843_));
 sky130_fd_sc_hd__mux4_1 _26236_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02644_));
 sky130_fd_sc_hd__mux4_1 _26237_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02645_));
 sky130_fd_sc_hd__mux4_1 _26238_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02646_));
 sky130_fd_sc_hd__mux4_1 _26239_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02647_));
 sky130_fd_sc_hd__mux4_2 _26240_ (.A0(_02644_),
    .A1(_02645_),
    .A2(_02646_),
    .A3(_02647_),
    .S0(net688),
    .S1(net686),
    .X(_02648_));
 sky130_fd_sc_hd__mux4_1 _26241_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02649_));
 sky130_fd_sc_hd__mux4_1 _26242_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02650_));
 sky130_fd_sc_hd__mux4_1 _26243_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02651_));
 sky130_fd_sc_hd__mux4_1 _26244_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net693),
    .S1(net698),
    .X(_02652_));
 sky130_fd_sc_hd__mux4_1 _26245_ (.A0(_02649_),
    .A1(_02650_),
    .A2(_02651_),
    .A3(_02652_),
    .S0(net688),
    .S1(net686),
    .X(_02653_));
 sky130_fd_sc_hd__mux2i_4 _26246_ (.A0(_02648_),
    .A1(_02653_),
    .S(net684),
    .Y(_02654_));
 sky130_fd_sc_hd__xnor2_1 _26247_ (.A(_11712_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__xnor2_2 _26248_ (.A(_11246_),
    .B(_02655_),
    .Y(_11846_));
 sky130_fd_sc_hd__mux4_1 _26249_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net621),
    .S1(net625),
    .X(_02656_));
 sky130_fd_sc_hd__mux4_1 _26250_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net621),
    .S1(net625),
    .X(_02657_));
 sky130_fd_sc_hd__mux4_1 _26251_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net621),
    .S1(net625),
    .X(_02658_));
 sky130_fd_sc_hd__mux4_1 _26252_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net621),
    .S1(net625),
    .X(_02659_));
 sky130_fd_sc_hd__mux4_4 _26253_ (.A0(_02656_),
    .A1(_02657_),
    .A2(_02658_),
    .A3(_02659_),
    .S0(net617),
    .S1(net613),
    .X(_02660_));
 sky130_fd_sc_hd__mux4_1 _26254_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net622),
    .S1(net628),
    .X(_02661_));
 sky130_fd_sc_hd__mux4_1 _26255_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net621),
    .S1(net625),
    .X(_02662_));
 sky130_fd_sc_hd__mux4_1 _26256_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net621),
    .S1(net625),
    .X(_02663_));
 sky130_fd_sc_hd__mux4_1 _26257_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net621),
    .S1(net625),
    .X(_02664_));
 sky130_fd_sc_hd__mux4_1 _26258_ (.A0(_02661_),
    .A1(_02662_),
    .A2(_02663_),
    .A3(_02664_),
    .S0(net617),
    .S1(net613),
    .X(_02665_));
 sky130_fd_sc_hd__mux2i_4 _26259_ (.A0(_02660_),
    .A1(_02665_),
    .S(net611),
    .Y(_02666_));
 sky130_fd_sc_hd__xnor2_1 _26260_ (.A(_02618_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__xnor2_1 _26261_ (.A(_11497_),
    .B(_02667_),
    .Y(_11851_));
 sky130_fd_sc_hd__mux4_1 _26262_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net694),
    .S1(net700),
    .X(_02668_));
 sky130_fd_sc_hd__mux4_1 _26263_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net694),
    .S1(net700),
    .X(_02669_));
 sky130_fd_sc_hd__mux4_1 _26264_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net694),
    .S1(net700),
    .X(_02670_));
 sky130_fd_sc_hd__mux4_1 _26265_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net694),
    .S1(net700),
    .X(_02671_));
 sky130_fd_sc_hd__mux4_4 _26266_ (.A0(_02668_),
    .A1(_02669_),
    .A2(_02670_),
    .A3(_02671_),
    .S0(net688),
    .S1(net686),
    .X(_02672_));
 sky130_fd_sc_hd__mux4_1 _26267_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net694),
    .S1(net698),
    .X(_02673_));
 sky130_fd_sc_hd__mux4_1 _26268_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net694),
    .S1(net698),
    .X(_02674_));
 sky130_fd_sc_hd__mux4_1 _26269_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net694),
    .S1(net698),
    .X(_02675_));
 sky130_fd_sc_hd__mux4_1 _26270_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net694),
    .S1(net698),
    .X(_02676_));
 sky130_fd_sc_hd__mux4_1 _26271_ (.A0(_02673_),
    .A1(_02674_),
    .A2(_02675_),
    .A3(_02676_),
    .S0(net688),
    .S1(net686),
    .X(_02677_));
 sky130_fd_sc_hd__mux2i_4 _26272_ (.A0(_02672_),
    .A1(_02677_),
    .S(net684),
    .Y(_02678_));
 sky130_fd_sc_hd__xnor2_1 _26273_ (.A(_02571_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__xnor2_2 _26274_ (.A(_11362_),
    .B(_02679_),
    .Y(_11854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_259 ();
 sky130_fd_sc_hd__mux4_1 _26277_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02682_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_257 ();
 sky130_fd_sc_hd__mux4_1 _26280_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_255 ();
 sky130_fd_sc_hd__mux4_1 _26283_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_253 ();
 sky130_fd_sc_hd__mux4_1 _26286_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_251 ();
 sky130_fd_sc_hd__mux4_2 _26289_ (.A0(_02682_),
    .A1(_02685_),
    .A2(_02688_),
    .A3(_02691_),
    .S0(net616),
    .S1(net614),
    .X(_02694_));
 sky130_fd_sc_hd__mux4_1 _26290_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02695_));
 sky130_fd_sc_hd__mux4_1 _26291_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02696_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_249 ();
 sky130_fd_sc_hd__mux4_1 _26294_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_247 ();
 sky130_fd_sc_hd__mux4_1 _26297_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net618),
    .S1(net626),
    .X(_02702_));
 sky130_fd_sc_hd__mux4_1 _26298_ (.A0(_02695_),
    .A1(_02696_),
    .A2(_02699_),
    .A3(_02702_),
    .S0(net616),
    .S1(net614),
    .X(_02703_));
 sky130_fd_sc_hd__mux2i_4 _26299_ (.A0(_02694_),
    .A1(_02703_),
    .S(net611),
    .Y(_02704_));
 sky130_fd_sc_hd__xnor2_1 _26300_ (.A(_02642_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__xnor2_1 _26301_ (.A(_11535_),
    .B(_02705_),
    .Y(_11859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_245 ();
 sky130_fd_sc_hd__mux4_1 _26304_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_02708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_243 ();
 sky130_fd_sc_hd__mux4_1 _26307_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_02711_));
 sky130_fd_sc_hd__mux4_1 _26308_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_02712_));
 sky130_fd_sc_hd__mux4_1 _26309_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_02713_));
 sky130_fd_sc_hd__mux4_4 _26310_ (.A0(_02708_),
    .A1(_02711_),
    .A2(_02712_),
    .A3(_02713_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_02714_));
 sky130_fd_sc_hd__mux4_1 _26311_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(\count15_1[2] ),
    .S1(net701),
    .X(_02715_));
 sky130_fd_sc_hd__mux4_1 _26312_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(\count15_1[2] ),
    .S1(net701),
    .X(_02716_));
 sky130_fd_sc_hd__mux4_1 _26313_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(\count15_1[2] ),
    .S1(net701),
    .X(_02717_));
 sky130_fd_sc_hd__mux4_1 _26314_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(\count15_1[2] ),
    .S1(net701),
    .X(_02718_));
 sky130_fd_sc_hd__mux4_2 _26315_ (.A0(_02715_),
    .A1(_02716_),
    .A2(_02717_),
    .A3(_02718_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_02719_));
 sky130_fd_sc_hd__mux2i_4 _26316_ (.A0(_02714_),
    .A1(_02719_),
    .S(\count15_1[5] ),
    .Y(_02720_));
 sky130_fd_sc_hd__xnor2_1 _26317_ (.A(_02595_),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__xnor2_2 _26318_ (.A(_11444_),
    .B(_02721_),
    .Y(_11862_));
 sky130_fd_sc_hd__mux4_1 _26319_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net618),
    .S1(net626),
    .X(_02722_));
 sky130_fd_sc_hd__mux4_1 _26320_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net618),
    .S1(net626),
    .X(_02723_));
 sky130_fd_sc_hd__mux4_1 _26321_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net618),
    .S1(net626),
    .X(_02724_));
 sky130_fd_sc_hd__mux4_1 _26322_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net618),
    .S1(net626),
    .X(_02725_));
 sky130_fd_sc_hd__mux4_4 _26323_ (.A0(_02722_),
    .A1(_02723_),
    .A2(_02724_),
    .A3(_02725_),
    .S0(net615),
    .S1(net612),
    .X(_02726_));
 sky130_fd_sc_hd__mux4_1 _26324_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net623),
    .S1(net628),
    .X(_02727_));
 sky130_fd_sc_hd__mux4_1 _26325_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net623),
    .S1(net628),
    .X(_02728_));
 sky130_fd_sc_hd__mux4_1 _26326_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net623),
    .S1(net628),
    .X(_02729_));
 sky130_fd_sc_hd__mux4_1 _26327_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net623),
    .S1(net628),
    .X(_02730_));
 sky130_fd_sc_hd__mux4_1 _26328_ (.A0(_02727_),
    .A1(_02728_),
    .A2(_02729_),
    .A3(_02730_),
    .S0(net617),
    .S1(net613),
    .X(_02731_));
 sky130_fd_sc_hd__mux2i_4 _26329_ (.A0(_02726_),
    .A1(_02731_),
    .S(net611),
    .Y(_02732_));
 sky130_fd_sc_hd__xnor2_2 _26330_ (.A(_02666_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__xnor2_4 _26331_ (.A(_11597_),
    .B(_02733_),
    .Y(_11867_));
 sky130_fd_sc_hd__mux4_1 _26332_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(\count15_1[2] ),
    .S1(net697),
    .X(_02734_));
 sky130_fd_sc_hd__mux4_1 _26333_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_02735_));
 sky130_fd_sc_hd__mux4_1 _26334_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_02736_));
 sky130_fd_sc_hd__mux4_1 _26335_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_02737_));
 sky130_fd_sc_hd__mux4_4 _26336_ (.A0(_02734_),
    .A1(_02735_),
    .A2(_02736_),
    .A3(_02737_),
    .S0(\count15_1[3] ),
    .S1(net685),
    .X(_02738_));
 sky130_fd_sc_hd__mux4_1 _26337_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net692),
    .S1(\count15_1[1] ),
    .X(_02739_));
 sky130_fd_sc_hd__mux4_1 _26338_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net692),
    .S1(\count15_1[1] ),
    .X(_02740_));
 sky130_fd_sc_hd__mux4_1 _26339_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net692),
    .S1(\count15_1[1] ),
    .X(_02741_));
 sky130_fd_sc_hd__mux4_1 _26340_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net692),
    .S1(\count15_1[1] ),
    .X(_02742_));
 sky130_fd_sc_hd__mux4_1 _26341_ (.A0(_02739_),
    .A1(_02740_),
    .A2(_02741_),
    .A3(_02742_),
    .S0(net687),
    .S1(net685),
    .X(_02743_));
 sky130_fd_sc_hd__mux2i_4 _26342_ (.A0(_02738_),
    .A1(_02743_),
    .S(net683),
    .Y(_02744_));
 sky130_fd_sc_hd__xnor2_1 _26343_ (.A(_11512_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__xnor2_2 _26344_ (.A(_11208_),
    .B(_02745_),
    .Y(_11870_));
 sky130_fd_sc_hd__mux4_1 _26345_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net618),
    .S1(net626),
    .X(_02746_));
 sky130_fd_sc_hd__mux4_1 _26346_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net618),
    .S1(net626),
    .X(_02747_));
 sky130_fd_sc_hd__mux4_1 _26347_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net618),
    .S1(net626),
    .X(_02748_));
 sky130_fd_sc_hd__mux4_1 _26348_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net618),
    .S1(net626),
    .X(_02749_));
 sky130_fd_sc_hd__mux4_2 _26349_ (.A0(_02746_),
    .A1(_02747_),
    .A2(_02748_),
    .A3(_02749_),
    .S0(net615),
    .S1(net612),
    .X(_02750_));
 sky130_fd_sc_hd__mux4_1 _26350_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net623),
    .S1(net625),
    .X(_02751_));
 sky130_fd_sc_hd__mux4_1 _26351_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net623),
    .S1(net625),
    .X(_02752_));
 sky130_fd_sc_hd__mux4_1 _26352_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net623),
    .S1(net625),
    .X(_02753_));
 sky130_fd_sc_hd__mux4_1 _26353_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net623),
    .S1(net625),
    .X(_02754_));
 sky130_fd_sc_hd__mux4_1 _26354_ (.A0(_02751_),
    .A1(_02752_),
    .A2(_02753_),
    .A3(_02754_),
    .S0(net615),
    .S1(net612),
    .X(_02755_));
 sky130_fd_sc_hd__mux2i_4 _26355_ (.A0(_02750_),
    .A1(_02755_),
    .S(net610),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_1 _26356_ (.A(_02704_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__xnor2_2 _26357_ (.A(_11643_),
    .B(_02757_),
    .Y(_11875_));
 sky130_fd_sc_hd__mux4_1 _26358_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02758_));
 sky130_fd_sc_hd__mux4_1 _26359_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02759_));
 sky130_fd_sc_hd__mux4_1 _26360_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02760_));
 sky130_fd_sc_hd__mux4_1 _26361_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02761_));
 sky130_fd_sc_hd__mux4_4 _26362_ (.A0(_02758_),
    .A1(_02759_),
    .A2(_02760_),
    .A3(_02761_),
    .S0(net687),
    .S1(net685),
    .X(_02762_));
 sky130_fd_sc_hd__mux4_1 _26363_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02763_));
 sky130_fd_sc_hd__mux4_1 _26364_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02764_));
 sky130_fd_sc_hd__mux4_1 _26365_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02765_));
 sky130_fd_sc_hd__mux4_1 _26366_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net691),
    .S1(net700),
    .X(_02766_));
 sky130_fd_sc_hd__mux4_1 _26367_ (.A0(_02763_),
    .A1(_02764_),
    .A2(_02765_),
    .A3(_02766_),
    .S0(net687),
    .S1(net685),
    .X(_02767_));
 sky130_fd_sc_hd__mux2i_4 _26368_ (.A0(_02762_),
    .A1(_02767_),
    .S(net683),
    .Y(_02768_));
 sky130_fd_sc_hd__xnor2_1 _26369_ (.A(_11574_),
    .B(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__xnor2_1 _26370_ (.A(_11246_),
    .B(_02769_),
    .Y(_11878_));
 sky130_fd_sc_hd__mux4_1 _26371_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net618),
    .S1(net626),
    .X(_02770_));
 sky130_fd_sc_hd__mux4_1 _26372_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net618),
    .S1(net626),
    .X(_02771_));
 sky130_fd_sc_hd__mux4_1 _26373_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net618),
    .S1(net626),
    .X(_02772_));
 sky130_fd_sc_hd__mux4_1 _26374_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net618),
    .S1(net626),
    .X(_02773_));
 sky130_fd_sc_hd__mux4_2 _26375_ (.A0(_02770_),
    .A1(_02771_),
    .A2(_02772_),
    .A3(_02773_),
    .S0(net615),
    .S1(net612),
    .X(_02774_));
 sky130_fd_sc_hd__mux4_1 _26376_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net619),
    .S1(net627),
    .X(_02775_));
 sky130_fd_sc_hd__mux4_1 _26377_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net619),
    .S1(net627),
    .X(_02776_));
 sky130_fd_sc_hd__mux4_1 _26378_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net619),
    .S1(net627),
    .X(_02777_));
 sky130_fd_sc_hd__mux4_1 _26379_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net619),
    .S1(net627),
    .X(_02778_));
 sky130_fd_sc_hd__mux4_1 _26380_ (.A0(_02775_),
    .A1(_02776_),
    .A2(_02777_),
    .A3(_02778_),
    .S0(net615),
    .S1(net612),
    .X(_02779_));
 sky130_fd_sc_hd__mux2i_4 _26381_ (.A0(_02774_),
    .A1(_02779_),
    .S(net610),
    .Y(_02780_));
 sky130_fd_sc_hd__xnor2_2 _26382_ (.A(_02732_),
    .B(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__xnor2_4 _26383_ (.A(_11678_),
    .B(_02781_),
    .Y(_11883_));
 sky130_fd_sc_hd__xnor2_1 _26384_ (.A(_11362_),
    .B(_11609_),
    .Y(_02782_));
 sky130_fd_sc_hd__xnor2_1 _26385_ (.A(_11176_),
    .B(_02782_),
    .Y(_11886_));
 sky130_fd_sc_hd__mux4_1 _26386_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02783_));
 sky130_fd_sc_hd__mux4_1 _26387_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02784_));
 sky130_fd_sc_hd__mux4_1 _26388_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02785_));
 sky130_fd_sc_hd__mux4_1 _26389_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02786_));
 sky130_fd_sc_hd__mux4_2 _26390_ (.A0(_02783_),
    .A1(_02784_),
    .A2(_02785_),
    .A3(_02786_),
    .S0(net616),
    .S1(net614),
    .X(_02787_));
 sky130_fd_sc_hd__mux4_1 _26391_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02788_));
 sky130_fd_sc_hd__mux4_1 _26392_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02789_));
 sky130_fd_sc_hd__mux4_1 _26393_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02790_));
 sky130_fd_sc_hd__mux4_1 _26394_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net619),
    .S1(net627),
    .X(_02791_));
 sky130_fd_sc_hd__mux4_1 _26395_ (.A0(_02788_),
    .A1(_02789_),
    .A2(_02790_),
    .A3(_02791_),
    .S0(net616),
    .S1(net614),
    .X(_02792_));
 sky130_fd_sc_hd__mux2i_4 _26396_ (.A0(_02787_),
    .A1(_02792_),
    .S(net611),
    .Y(_02793_));
 sky130_fd_sc_hd__xnor2_2 _26397_ (.A(_02756_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__xnor2_2 _26398_ (.A(_11724_),
    .B(_02794_),
    .Y(_11891_));
 sky130_fd_sc_hd__xnor2_1 _26399_ (.A(_11444_),
    .B(_11666_),
    .Y(_02795_));
 sky130_fd_sc_hd__xnor2_1 _26400_ (.A(_11259_),
    .B(_02795_),
    .Y(_11894_));
 sky130_fd_sc_hd__mux4_1 _26401_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02796_));
 sky130_fd_sc_hd__mux4_1 _26402_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02797_));
 sky130_fd_sc_hd__mux4_1 _26403_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02798_));
 sky130_fd_sc_hd__mux4_1 _26404_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02799_));
 sky130_fd_sc_hd__mux4_4 _26405_ (.A0(_02796_),
    .A1(_02797_),
    .A2(_02798_),
    .A3(_02799_),
    .S0(net616),
    .S1(\count2_1[4] ),
    .X(_02800_));
 sky130_fd_sc_hd__mux4_1 _26406_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02801_));
 sky130_fd_sc_hd__mux4_1 _26407_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02802_));
 sky130_fd_sc_hd__mux4_1 _26408_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02803_));
 sky130_fd_sc_hd__mux4_1 _26409_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net620),
    .S1(net624),
    .X(_02804_));
 sky130_fd_sc_hd__mux4_1 _26410_ (.A0(_02801_),
    .A1(_02802_),
    .A2(_02803_),
    .A3(_02804_),
    .S0(net616),
    .S1(net614),
    .X(_02805_));
 sky130_fd_sc_hd__mux2i_4 _26411_ (.A0(_02800_),
    .A1(_02805_),
    .S(net611),
    .Y(_02806_));
 sky130_fd_sc_hd__xnor2_1 _26412_ (.A(_02780_),
    .B(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__xnor2_2 _26413_ (.A(_02583_),
    .B(_02807_),
    .Y(_11899_));
 sky130_fd_sc_hd__xnor2_1 _26414_ (.A(_11512_),
    .B(_11701_),
    .Y(_02808_));
 sky130_fd_sc_hd__xnor2_1 _26415_ (.A(_11374_),
    .B(_02808_),
    .Y(_11902_));
 sky130_fd_sc_hd__mux4_1 _26416_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02809_));
 sky130_fd_sc_hd__mux4_1 _26417_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02810_));
 sky130_fd_sc_hd__mux4_1 _26418_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02811_));
 sky130_fd_sc_hd__mux4_1 _26419_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02812_));
 sky130_fd_sc_hd__mux4_4 _26420_ (.A0(_02809_),
    .A1(_02810_),
    .A2(_02811_),
    .A3(_02812_),
    .S0(net616),
    .S1(\count2_1[4] ),
    .X(_02813_));
 sky130_fd_sc_hd__mux4_1 _26421_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02814_));
 sky130_fd_sc_hd__mux4_1 _26422_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02815_));
 sky130_fd_sc_hd__mux4_1 _26423_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02816_));
 sky130_fd_sc_hd__mux4_1 _26424_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net620),
    .S1(net624),
    .X(_02817_));
 sky130_fd_sc_hd__mux4_1 _26425_ (.A0(_02814_),
    .A1(_02815_),
    .A2(_02816_),
    .A3(_02817_),
    .S0(net616),
    .S1(net614),
    .X(_02818_));
 sky130_fd_sc_hd__mux2i_4 _26426_ (.A0(_02813_),
    .A1(_02818_),
    .S(net611),
    .Y(_02819_));
 sky130_fd_sc_hd__xnor2_1 _26427_ (.A(_02793_),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__xnor2_2 _26428_ (.A(_02618_),
    .B(_02820_),
    .Y(_11907_));
 sky130_fd_sc_hd__xnor2_1 _26429_ (.A(_11574_),
    .B(_11736_),
    .Y(_02821_));
 sky130_fd_sc_hd__xnor2_1 _26430_ (.A(_11457_),
    .B(_02821_),
    .Y(_11910_));
 sky130_fd_sc_hd__mux4_1 _26431_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net618),
    .S1(net626),
    .X(_02822_));
 sky130_fd_sc_hd__mux4_1 _26432_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net618),
    .S1(net626),
    .X(_02823_));
 sky130_fd_sc_hd__mux4_1 _26433_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net618),
    .S1(net626),
    .X(_02824_));
 sky130_fd_sc_hd__mux4_1 _26434_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net618),
    .S1(net626),
    .X(_02825_));
 sky130_fd_sc_hd__mux4_2 _26435_ (.A0(_02822_),
    .A1(_02823_),
    .A2(_02824_),
    .A3(_02825_),
    .S0(net615),
    .S1(net612),
    .X(_02826_));
 sky130_fd_sc_hd__mux4_1 _26436_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net623),
    .S1(net625),
    .X(_02827_));
 sky130_fd_sc_hd__mux4_1 _26437_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net621),
    .S1(net625),
    .X(_02828_));
 sky130_fd_sc_hd__mux4_1 _26438_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net623),
    .S1(net625),
    .X(_02829_));
 sky130_fd_sc_hd__mux4_1 _26439_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net621),
    .S1(net625),
    .X(_02830_));
 sky130_fd_sc_hd__mux4_1 _26440_ (.A0(_02827_),
    .A1(_02828_),
    .A2(_02829_),
    .A3(_02830_),
    .S0(net615),
    .S1(net612),
    .X(_02831_));
 sky130_fd_sc_hd__mux2i_4 _26441_ (.A0(_02826_),
    .A1(_02831_),
    .S(net610),
    .Y(_02832_));
 sky130_fd_sc_hd__xnor2_1 _26442_ (.A(_02806_),
    .B(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__xnor2_2 _26443_ (.A(_02642_),
    .B(_02833_),
    .Y(_11915_));
 sky130_fd_sc_hd__xnor2_1 _26444_ (.A(_11609_),
    .B(_02606_),
    .Y(_02834_));
 sky130_fd_sc_hd__xnor2_2 _26445_ (.A(_11234_),
    .B(_02834_),
    .Y(_11918_));
 sky130_fd_sc_hd__mux4_1 _26446_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02835_));
 sky130_fd_sc_hd__mux4_1 _26447_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02836_));
 sky130_fd_sc_hd__mux4_1 _26448_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02837_));
 sky130_fd_sc_hd__mux4_1 _26449_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02838_));
 sky130_fd_sc_hd__mux4_4 _26450_ (.A0(_02835_),
    .A1(_02836_),
    .A2(_02837_),
    .A3(_02838_),
    .S0(net615),
    .S1(net612),
    .X(_02839_));
 sky130_fd_sc_hd__mux4_1 _26451_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02840_));
 sky130_fd_sc_hd__mux4_1 _26452_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02841_));
 sky130_fd_sc_hd__mux4_1 _26453_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02842_));
 sky130_fd_sc_hd__mux4_1 _26454_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net621),
    .S1(net625),
    .X(_02843_));
 sky130_fd_sc_hd__mux4_1 _26455_ (.A0(_02840_),
    .A1(_02841_),
    .A2(_02842_),
    .A3(_02843_),
    .S0(net617),
    .S1(net613),
    .X(_02844_));
 sky130_fd_sc_hd__mux2i_4 _26456_ (.A0(_02839_),
    .A1(_02844_),
    .S(net610),
    .Y(_02845_));
 sky130_fd_sc_hd__xnor2_1 _26457_ (.A(_02819_),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__xnor2_2 _26458_ (.A(_02666_),
    .B(_02846_),
    .Y(_11923_));
 sky130_fd_sc_hd__xnor2_1 _26459_ (.A(_11666_),
    .B(_02630_),
    .Y(_02847_));
 sky130_fd_sc_hd__xnor2_1 _26460_ (.A(_11271_),
    .B(_02847_),
    .Y(_11926_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_242 ();
 sky130_fd_sc_hd__mux4_1 _26462_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02849_));
 sky130_fd_sc_hd__mux4_1 _26463_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02850_));
 sky130_fd_sc_hd__mux4_1 _26464_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02851_));
 sky130_fd_sc_hd__mux4_1 _26465_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count2_1[2] ),
    .S1(net624),
    .X(_02852_));
 sky130_fd_sc_hd__mux4_4 _26466_ (.A0(_02849_),
    .A1(_02850_),
    .A2(_02851_),
    .A3(_02852_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02853_));
 sky130_fd_sc_hd__mux4_1 _26467_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net620),
    .S1(net627),
    .X(_02854_));
 sky130_fd_sc_hd__mux4_1 _26468_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net620),
    .S1(net627),
    .X(_02855_));
 sky130_fd_sc_hd__mux4_1 _26469_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net620),
    .S1(\count2_1[1] ),
    .X(_02856_));
 sky130_fd_sc_hd__mux4_1 _26470_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net623),
    .S1(\count2_1[1] ),
    .X(_02857_));
 sky130_fd_sc_hd__mux4_1 _26471_ (.A0(_02854_),
    .A1(_02855_),
    .A2(_02856_),
    .A3(_02857_),
    .S0(net616),
    .S1(net614),
    .X(_02858_));
 sky130_fd_sc_hd__mux2i_4 _26472_ (.A0(_02853_),
    .A1(_02858_),
    .S(\count2_1[5] ),
    .Y(_02859_));
 sky130_fd_sc_hd__xnor2_1 _26473_ (.A(_02832_),
    .B(_02859_),
    .Y(_11931_));
 sky130_fd_sc_hd__xnor2_1 _26474_ (.A(_11701_),
    .B(_02654_),
    .Y(_02860_));
 sky130_fd_sc_hd__xnor2_2 _26475_ (.A(_11385_),
    .B(_02860_),
    .Y(_11934_));
 sky130_fd_sc_hd__mux4_1 _26476_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net622),
    .S1(net628),
    .X(_02861_));
 sky130_fd_sc_hd__mux4_1 _26477_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net622),
    .S1(net628),
    .X(_02862_));
 sky130_fd_sc_hd__mux4_1 _26478_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net622),
    .S1(net628),
    .X(_02863_));
 sky130_fd_sc_hd__mux4_1 _26479_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net622),
    .S1(net628),
    .X(_02864_));
 sky130_fd_sc_hd__mux4_4 _26480_ (.A0(_02861_),
    .A1(_02862_),
    .A2(_02863_),
    .A3(_02864_),
    .S0(net617),
    .S1(net613),
    .X(_02865_));
 sky130_fd_sc_hd__mux4_1 _26481_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net623),
    .S1(net628),
    .X(_02866_));
 sky130_fd_sc_hd__mux4_1 _26482_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net623),
    .S1(net628),
    .X(_02867_));
 sky130_fd_sc_hd__mux4_1 _26483_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net623),
    .S1(net628),
    .X(_02868_));
 sky130_fd_sc_hd__mux4_1 _26484_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net623),
    .S1(net628),
    .X(_02869_));
 sky130_fd_sc_hd__mux4_1 _26485_ (.A0(_02866_),
    .A1(_02867_),
    .A2(_02868_),
    .A3(_02869_),
    .S0(net617),
    .S1(net613),
    .X(_02870_));
 sky130_fd_sc_hd__mux2i_4 _26486_ (.A0(_02865_),
    .A1(_02870_),
    .S(net611),
    .Y(_02871_));
 sky130_fd_sc_hd__xnor2_1 _26487_ (.A(_02845_),
    .B(_02871_),
    .Y(_11939_));
 sky130_fd_sc_hd__xnor2_1 _26488_ (.A(_11736_),
    .B(_02678_),
    .Y(_02872_));
 sky130_fd_sc_hd__xnor2_1 _26489_ (.A(_11468_),
    .B(_02872_),
    .Y(_11942_));
 sky130_fd_sc_hd__xnor2_1 _26490_ (.A(_11338_),
    .B(_02859_),
    .Y(_11947_));
 sky130_fd_sc_hd__xnor2_1 _26491_ (.A(_02606_),
    .B(_02720_),
    .Y(_02873_));
 sky130_fd_sc_hd__xnor2_1 _26492_ (.A(_11523_),
    .B(_02873_),
    .Y(_11950_));
 sky130_fd_sc_hd__xnor2_1 _26493_ (.A(_11411_),
    .B(_02871_),
    .Y(_11955_));
 sky130_fd_sc_hd__xnor2_1 _26494_ (.A(_02630_),
    .B(_02744_),
    .Y(_02874_));
 sky130_fd_sc_hd__xnor2_2 _26495_ (.A(_11562_),
    .B(_02874_),
    .Y(_11958_));
 sky130_fd_sc_hd__xnor2_2 _26496_ (.A(_11338_),
    .B(_11486_),
    .Y(_11963_));
 sky130_fd_sc_hd__xnor2_1 _26497_ (.A(_02654_),
    .B(_02768_),
    .Y(_02875_));
 sky130_fd_sc_hd__xnor2_1 _26498_ (.A(_11620_),
    .B(_02875_),
    .Y(_11966_));
 sky130_fd_sc_hd__xnor2_1 _26499_ (.A(_11411_),
    .B(_11546_),
    .Y(_11971_));
 sky130_fd_sc_hd__xnor2_1 _26500_ (.A(_11655_),
    .B(_02678_),
    .Y(_02876_));
 sky130_fd_sc_hd__xnor2_1 _26501_ (.A(_11176_),
    .B(_02876_),
    .Y(_11974_));
 sky130_fd_sc_hd__xnor2_1 _26502_ (.A(_11486_),
    .B(_11586_),
    .Y(_11979_));
 sky130_fd_sc_hd__xnor2_1 _26503_ (.A(_11259_),
    .B(_11712_),
    .Y(_11982_));
 sky130_fd_sc_hd__xnor2_1 _26504_ (.A(_11546_),
    .B(_11632_),
    .Y(_11987_));
 sky130_fd_sc_hd__xnor2_1 _26505_ (.A(_11374_),
    .B(_02571_),
    .Y(_11990_));
 sky130_fd_sc_hd__xnor2_2 _26506_ (.A(_11586_),
    .B(_11689_),
    .Y(_11995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_233 ();
 sky130_fd_sc_hd__mux4_1 _26516_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net602),
    .S1(net605),
    .X(_02886_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_231 ();
 sky130_fd_sc_hd__mux4_1 _26519_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net602),
    .S1(net605),
    .X(_02889_));
 sky130_fd_sc_hd__mux4_1 _26520_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net602),
    .S1(net605),
    .X(_02890_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_228 ();
 sky130_fd_sc_hd__mux4_1 _26524_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net602),
    .S1(net605),
    .X(_02894_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_223 ();
 sky130_fd_sc_hd__mux4_4 _26530_ (.A0(_02886_),
    .A1(_02889_),
    .A2(_02890_),
    .A3(_02894_),
    .S0(net596),
    .S1(net595),
    .X(_02900_));
 sky130_fd_sc_hd__mux4_1 _26531_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_02901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_221 ();
 sky130_fd_sc_hd__mux4_1 _26534_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net604),
    .S1(net609),
    .X(_02904_));
 sky130_fd_sc_hd__mux4_1 _26535_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_02905_));
 sky130_fd_sc_hd__mux4_1 _26536_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net604),
    .S1(net609),
    .X(_02906_));
 sky130_fd_sc_hd__mux4_1 _26537_ (.A0(_02901_),
    .A1(_02904_),
    .A2(_02905_),
    .A3(_02906_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_02907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_219 ();
 sky130_fd_sc_hd__mux2i_4 _26540_ (.A0(_02900_),
    .A1(_02907_),
    .S(net593),
    .Y(_02910_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__mux4_1 _26544_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net604),
    .S1(net609),
    .X(_02914_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__mux4_1 _26547_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net604),
    .S1(net609),
    .X(_02917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__mux4_1 _26550_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net604),
    .S1(net609),
    .X(_02920_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__mux4_1 _26552_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net604),
    .S1(net609),
    .X(_02922_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_209 ();
 sky130_fd_sc_hd__mux4_4 _26555_ (.A0(_02914_),
    .A1(_02917_),
    .A2(_02920_),
    .A3(_02922_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_02925_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_208 ();
 sky130_fd_sc_hd__mux4_1 _26557_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net602),
    .S1(net609),
    .X(_02927_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_206 ();
 sky130_fd_sc_hd__mux4_1 _26560_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net602),
    .S1(net609),
    .X(_02930_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_204 ();
 sky130_fd_sc_hd__mux4_1 _26563_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net602),
    .S1(net609),
    .X(_02933_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_202 ();
 sky130_fd_sc_hd__mux4_1 _26566_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net602),
    .S1(net609),
    .X(_02936_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_200 ();
 sky130_fd_sc_hd__mux4_1 _26569_ (.A0(_02927_),
    .A1(_02930_),
    .A2(_02933_),
    .A3(_02936_),
    .S0(net596),
    .S1(\count2_2[4] ),
    .X(_02939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_199 ();
 sky130_fd_sc_hd__mux2i_4 _26571_ (.A0(_02925_),
    .A1(_02939_),
    .S(net593),
    .Y(_02941_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_198 ();
 sky130_fd_sc_hd__mux4_1 _26573_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net601),
    .S1(net608),
    .X(_02943_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_196 ();
 sky130_fd_sc_hd__mux4_1 _26576_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net601),
    .S1(net608),
    .X(_02946_));
 sky130_fd_sc_hd__mux4_1 _26577_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net601),
    .S1(net608),
    .X(_02947_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_194 ();
 sky130_fd_sc_hd__mux4_1 _26580_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net601),
    .S1(net608),
    .X(_02950_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_192 ();
 sky130_fd_sc_hd__mux4_2 _26583_ (.A0(_02943_),
    .A1(_02946_),
    .A2(_02947_),
    .A3(_02950_),
    .S0(net597),
    .S1(net594),
    .X(_02953_));
 sky130_fd_sc_hd__mux4_1 _26584_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_02954_));
 sky130_fd_sc_hd__mux4_1 _26585_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_02955_));
 sky130_fd_sc_hd__mux4_1 _26586_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_02956_));
 sky130_fd_sc_hd__mux4_1 _26587_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_02957_));
 sky130_fd_sc_hd__mux4_1 _26588_ (.A0(_02954_),
    .A1(_02955_),
    .A2(_02956_),
    .A3(_02957_),
    .S0(net597),
    .S1(net594),
    .X(_02958_));
 sky130_fd_sc_hd__mux2i_4 _26589_ (.A0(_02953_),
    .A1(_02958_),
    .S(net592),
    .Y(_02959_));
 sky130_fd_sc_hd__xnor2_1 _26590_ (.A(_02941_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__xnor2_1 _26591_ (.A(_02910_),
    .B(_02960_),
    .Y(_12000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_183 ();
 sky130_fd_sc_hd__mux4_1 _26601_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net672),
    .S1(net679),
    .X(_02970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_179 ();
 sky130_fd_sc_hd__mux4_1 _26606_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net672),
    .S1(net679),
    .X(_02975_));
 sky130_fd_sc_hd__mux4_1 _26607_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net672),
    .S1(net679),
    .X(_02976_));
 sky130_fd_sc_hd__mux4_1 _26608_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net672),
    .S1(net679),
    .X(_02977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_174 ();
 sky130_fd_sc_hd__mux4_2 _26614_ (.A0(_02970_),
    .A1(_02975_),
    .A2(_02976_),
    .A3(_02977_),
    .S0(net671),
    .S1(net667),
    .X(_02983_));
 sky130_fd_sc_hd__mux4_1 _26615_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net672),
    .S1(net679),
    .X(_02984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_170 ();
 sky130_fd_sc_hd__mux4_1 _26620_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net672),
    .S1(net679),
    .X(_02989_));
 sky130_fd_sc_hd__mux4_1 _26621_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net672),
    .S1(net679),
    .X(_02990_));
 sky130_fd_sc_hd__mux4_1 _26622_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net672),
    .S1(\count15_2[1] ),
    .X(_02991_));
 sky130_fd_sc_hd__mux4_1 _26623_ (.A0(_02984_),
    .A1(_02989_),
    .A2(_02990_),
    .A3(_02991_),
    .S0(net671),
    .S1(net668),
    .X(_02992_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_168 ();
 sky130_fd_sc_hd__mux2i_4 _26626_ (.A0(_02983_),
    .A1(_02992_),
    .S(net665),
    .Y(_02995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_166 ();
 sky130_fd_sc_hd__mux4_1 _26629_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net677),
    .S1(net679),
    .X(_02998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_164 ();
 sky130_fd_sc_hd__mux4_1 _26632_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net677),
    .S1(net679),
    .X(_03001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_162 ();
 sky130_fd_sc_hd__mux4_1 _26635_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net677),
    .S1(net679),
    .X(_03004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_160 ();
 sky130_fd_sc_hd__mux4_1 _26638_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net677),
    .S1(net679),
    .X(_03007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_158 ();
 sky130_fd_sc_hd__mux4_2 _26641_ (.A0(_02998_),
    .A1(_03001_),
    .A2(_03004_),
    .A3(_03007_),
    .S0(net669),
    .S1(net667),
    .X(_03010_));
 sky130_fd_sc_hd__mux4_1 _26642_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net677),
    .S1(net679),
    .X(_03011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_157 ();
 sky130_fd_sc_hd__mux4_1 _26644_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net675),
    .S1(net679),
    .X(_03013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_155 ();
 sky130_fd_sc_hd__mux4_1 _26647_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net677),
    .S1(net679),
    .X(_03016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_153 ();
 sky130_fd_sc_hd__mux4_1 _26650_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net675),
    .S1(net679),
    .X(_03019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_151 ();
 sky130_fd_sc_hd__mux4_1 _26653_ (.A0(_03011_),
    .A1(_03013_),
    .A2(_03016_),
    .A3(_03019_),
    .S0(net671),
    .S1(net668),
    .X(_03022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_150 ();
 sky130_fd_sc_hd__mux2i_4 _26655_ (.A0(_03010_),
    .A1(_03022_),
    .S(\count15_2[5] ),
    .Y(_03024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_148 ();
 sky130_fd_sc_hd__mux4_1 _26658_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03027_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_146 ();
 sky130_fd_sc_hd__mux4_1 _26661_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03030_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_145 ();
 sky130_fd_sc_hd__mux4_1 _26663_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03032_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_144 ();
 sky130_fd_sc_hd__mux4_1 _26665_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_142 ();
 sky130_fd_sc_hd__mux4_4 _26668_ (.A0(_03027_),
    .A1(_03030_),
    .A2(_03032_),
    .A3(_03034_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_140 ();
 sky130_fd_sc_hd__mux4_1 _26671_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_138 ();
 sky130_fd_sc_hd__mux4_1 _26674_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_136 ();
 sky130_fd_sc_hd__mux4_1 _26677_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_134 ();
 sky130_fd_sc_hd__mux4_1 _26680_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03049_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__mux4_1 _26683_ (.A0(_03040_),
    .A1(_03043_),
    .A2(_03046_),
    .A3(_03049_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03052_));
 sky130_fd_sc_hd__mux2i_4 _26684_ (.A0(_03037_),
    .A1(_03052_),
    .S(\count15_2[5] ),
    .Y(_03053_));
 sky130_fd_sc_hd__xnor2_1 _26685_ (.A(_03024_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__xnor2_2 _26686_ (.A(_02995_),
    .B(_03054_),
    .Y(_11999_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_124 ();
 sky130_fd_sc_hd__mux4_1 _26695_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net561),
    .S1(net572),
    .X(_03063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_120 ();
 sky130_fd_sc_hd__mux4_1 _26700_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net561),
    .S1(net572),
    .X(_03068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_118 ();
 sky130_fd_sc_hd__mux4_1 _26703_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net561),
    .S1(net572),
    .X(_03071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_115 ();
 sky130_fd_sc_hd__mux4_1 _26707_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net561),
    .S1(net572),
    .X(_03075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_110 ();
 sky130_fd_sc_hd__mux4_2 _26713_ (.A0(_03063_),
    .A1(_03068_),
    .A2(_03071_),
    .A3(_03075_),
    .S0(net559),
    .S1(net555),
    .X(_03081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_108 ();
 sky130_fd_sc_hd__mux4_1 _26716_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net566),
    .S1(net571),
    .X(_03084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_106 ();
 sky130_fd_sc_hd__mux4_1 _26719_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net566),
    .S1(net571),
    .X(_03087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__mux4_1 _26722_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net566),
    .S1(net571),
    .X(_03090_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__mux4_1 _26725_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net566),
    .S1(net571),
    .X(_03093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__mux4_1 _26728_ (.A0(_03084_),
    .A1(_03087_),
    .A2(_03090_),
    .A3(_03093_),
    .S0(net559),
    .S1(net555),
    .X(_03096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_98 ();
 sky130_fd_sc_hd__mux2i_4 _26731_ (.A0(_03081_),
    .A1(_03096_),
    .S(net553),
    .Y(_11998_));
 sky130_fd_sc_hd__mux4_1 _26732_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net604),
    .S1(net609),
    .X(_03099_));
 sky130_fd_sc_hd__mux4_1 _26733_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net604),
    .S1(net609),
    .X(_03100_));
 sky130_fd_sc_hd__mux4_1 _26734_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net604),
    .S1(net609),
    .X(_03101_));
 sky130_fd_sc_hd__mux4_1 _26735_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net604),
    .S1(net609),
    .X(_03102_));
 sky130_fd_sc_hd__mux4_4 _26736_ (.A0(_03099_),
    .A1(_03100_),
    .A2(_03101_),
    .A3(_03102_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03103_));
 sky130_fd_sc_hd__mux4_1 _26737_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net604),
    .S1(net609),
    .X(_03104_));
 sky130_fd_sc_hd__mux4_1 _26738_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net603),
    .S1(net609),
    .X(_03105_));
 sky130_fd_sc_hd__mux4_1 _26739_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net604),
    .S1(net609),
    .X(_03106_));
 sky130_fd_sc_hd__mux4_1 _26740_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net603),
    .S1(net609),
    .X(_03107_));
 sky130_fd_sc_hd__mux4_2 _26741_ (.A0(_03104_),
    .A1(_03105_),
    .A2(_03106_),
    .A3(_03107_),
    .S0(net596),
    .S1(net595),
    .X(_03108_));
 sky130_fd_sc_hd__mux2i_4 _26742_ (.A0(_03103_),
    .A1(_03108_),
    .S(net593),
    .Y(_03109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_97 ();
 sky130_fd_sc_hd__mux4_1 _26744_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03111_));
 sky130_fd_sc_hd__mux4_1 _26745_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03112_));
 sky130_fd_sc_hd__mux4_1 _26746_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_96 ();
 sky130_fd_sc_hd__mux4_1 _26748_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03115_));
 sky130_fd_sc_hd__mux4_2 _26749_ (.A0(_03111_),
    .A1(_03112_),
    .A2(_03113_),
    .A3(_03115_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03116_));
 sky130_fd_sc_hd__mux4_1 _26750_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_95 ();
 sky130_fd_sc_hd__mux4_1 _26752_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03119_));
 sky130_fd_sc_hd__mux4_1 _26753_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03120_));
 sky130_fd_sc_hd__mux4_1 _26754_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(\count2_2[2] ),
    .S1(\count2_2[1] ),
    .X(_03121_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_94 ();
 sky130_fd_sc_hd__mux4_1 _26756_ (.A0(_03117_),
    .A1(_03119_),
    .A2(_03120_),
    .A3(_03121_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03123_));
 sky130_fd_sc_hd__mux2i_4 _26757_ (.A0(_03116_),
    .A1(_03123_),
    .S(net593),
    .Y(_03124_));
 sky130_fd_sc_hd__mux4_1 _26758_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net602),
    .S1(net605),
    .X(_03125_));
 sky130_fd_sc_hd__mux4_1 _26759_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net602),
    .S1(net605),
    .X(_03126_));
 sky130_fd_sc_hd__mux4_1 _26760_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net602),
    .S1(net605),
    .X(_03127_));
 sky130_fd_sc_hd__mux4_1 _26761_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net602),
    .S1(net605),
    .X(_03128_));
 sky130_fd_sc_hd__mux4_4 _26762_ (.A0(_03125_),
    .A1(_03126_),
    .A2(_03127_),
    .A3(_03128_),
    .S0(net596),
    .S1(net595),
    .X(_03129_));
 sky130_fd_sc_hd__mux4_1 _26763_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net603),
    .S1(net607),
    .X(_03130_));
 sky130_fd_sc_hd__mux4_1 _26764_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net603),
    .S1(net607),
    .X(_03131_));
 sky130_fd_sc_hd__mux4_1 _26765_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net603),
    .S1(net607),
    .X(_03132_));
 sky130_fd_sc_hd__mux4_1 _26766_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net603),
    .S1(net607),
    .X(_03133_));
 sky130_fd_sc_hd__mux4_1 _26767_ (.A0(_03130_),
    .A1(_03131_),
    .A2(_03132_),
    .A3(_03133_),
    .S0(net596),
    .S1(net595),
    .X(_03134_));
 sky130_fd_sc_hd__mux2i_4 _26768_ (.A0(_03129_),
    .A1(_03134_),
    .S(net593),
    .Y(_03135_));
 sky130_fd_sc_hd__xnor2_1 _26769_ (.A(_03124_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__xnor2_1 _26770_ (.A(_03109_),
    .B(_03136_),
    .Y(_12005_));
 sky130_fd_sc_hd__mux4_1 _26771_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03137_));
 sky130_fd_sc_hd__mux4_1 _26772_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03138_));
 sky130_fd_sc_hd__mux4_1 _26773_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03139_));
 sky130_fd_sc_hd__mux4_1 _26774_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03140_));
 sky130_fd_sc_hd__mux4_2 _26775_ (.A0(_03137_),
    .A1(_03138_),
    .A2(_03139_),
    .A3(_03140_),
    .S0(net669),
    .S1(net667),
    .X(_03141_));
 sky130_fd_sc_hd__mux4_1 _26776_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03142_));
 sky130_fd_sc_hd__mux4_1 _26777_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03143_));
 sky130_fd_sc_hd__mux4_1 _26778_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03144_));
 sky130_fd_sc_hd__mux4_1 _26779_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net673),
    .S1(net680),
    .X(_03145_));
 sky130_fd_sc_hd__mux4_1 _26780_ (.A0(_03142_),
    .A1(_03143_),
    .A2(_03144_),
    .A3(_03145_),
    .S0(net669),
    .S1(net667),
    .X(_03146_));
 sky130_fd_sc_hd__mux2i_4 _26781_ (.A0(_03141_),
    .A1(_03146_),
    .S(net666),
    .Y(_03147_));
 sky130_fd_sc_hd__mux4_1 _26782_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03148_));
 sky130_fd_sc_hd__mux4_1 _26783_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03149_));
 sky130_fd_sc_hd__mux4_1 _26784_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03150_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_93 ();
 sky130_fd_sc_hd__mux4_1 _26786_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03152_));
 sky130_fd_sc_hd__mux4_4 _26787_ (.A0(_03148_),
    .A1(_03149_),
    .A2(_03150_),
    .A3(_03152_),
    .S0(net670),
    .S1(net668),
    .X(_03153_));
 sky130_fd_sc_hd__mux4_1 _26788_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03154_));
 sky130_fd_sc_hd__mux4_1 _26789_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03155_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_91 ();
 sky130_fd_sc_hd__mux4_1 _26792_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_89 ();
 sky130_fd_sc_hd__mux4_1 _26795_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net675),
    .S1(net681),
    .X(_03161_));
 sky130_fd_sc_hd__mux4_1 _26796_ (.A0(_03154_),
    .A1(_03155_),
    .A2(_03158_),
    .A3(_03161_),
    .S0(net670),
    .S1(net668),
    .X(_03162_));
 sky130_fd_sc_hd__mux2i_4 _26797_ (.A0(_03153_),
    .A1(_03162_),
    .S(\count15_2[5] ),
    .Y(_03163_));
 sky130_fd_sc_hd__mux4_1 _26798_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03164_));
 sky130_fd_sc_hd__mux4_1 _26799_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03165_));
 sky130_fd_sc_hd__mux4_1 _26800_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03166_));
 sky130_fd_sc_hd__mux4_1 _26801_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03167_));
 sky130_fd_sc_hd__mux4_2 _26802_ (.A0(_03164_),
    .A1(_03165_),
    .A2(_03166_),
    .A3(_03167_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03168_));
 sky130_fd_sc_hd__mux4_1 _26803_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net674),
    .S1(net678),
    .X(_03169_));
 sky130_fd_sc_hd__mux4_1 _26804_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net674),
    .S1(net678),
    .X(_03170_));
 sky130_fd_sc_hd__mux4_1 _26805_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net674),
    .S1(net678),
    .X(_03171_));
 sky130_fd_sc_hd__mux4_1 _26806_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net674),
    .S1(net678),
    .X(_03172_));
 sky130_fd_sc_hd__mux4_1 _26807_ (.A0(_03169_),
    .A1(_03170_),
    .A2(_03171_),
    .A3(_03172_),
    .S0(net669),
    .S1(net667),
    .X(_03173_));
 sky130_fd_sc_hd__mux2i_4 _26808_ (.A0(_03168_),
    .A1(_03173_),
    .S(net666),
    .Y(_03174_));
 sky130_fd_sc_hd__xnor2_1 _26809_ (.A(_03163_),
    .B(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__xnor2_2 _26810_ (.A(_03147_),
    .B(_03175_),
    .Y(_12004_));
 sky130_fd_sc_hd__mux4_1 _26811_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net560),
    .S1(net570),
    .X(_03176_));
 sky130_fd_sc_hd__mux4_1 _26812_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net560),
    .S1(net570),
    .X(_03177_));
 sky130_fd_sc_hd__mux4_1 _26813_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net560),
    .S1(net570),
    .X(_03178_));
 sky130_fd_sc_hd__mux4_1 _26814_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net560),
    .S1(net570),
    .X(_03179_));
 sky130_fd_sc_hd__mux4_4 _26815_ (.A0(_03176_),
    .A1(_03177_),
    .A2(_03178_),
    .A3(_03179_),
    .S0(net557),
    .S1(net555),
    .X(_03180_));
 sky130_fd_sc_hd__mux4_1 _26816_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net566),
    .S1(net571),
    .X(_03181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_88 ();
 sky130_fd_sc_hd__mux4_1 _26818_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net566),
    .S1(net571),
    .X(_03183_));
 sky130_fd_sc_hd__mux4_1 _26819_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net566),
    .S1(net571),
    .X(_03184_));
 sky130_fd_sc_hd__mux4_1 _26820_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net566),
    .S1(net571),
    .X(_03185_));
 sky130_fd_sc_hd__mux4_1 _26821_ (.A0(_03181_),
    .A1(_03183_),
    .A2(_03184_),
    .A3(_03185_),
    .S0(net557),
    .S1(net555),
    .X(_03186_));
 sky130_fd_sc_hd__mux2i_4 _26822_ (.A0(_03180_),
    .A1(_03186_),
    .S(net553),
    .Y(_12003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_80 ();
 sky130_fd_sc_hd__mux4_1 _26831_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net641),
    .S1(net647),
    .X(_03195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_76 ();
 sky130_fd_sc_hd__mux4_1 _26836_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net641),
    .S1(net647),
    .X(_03200_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_74 ();
 sky130_fd_sc_hd__mux4_1 _26839_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net641),
    .S1(net647),
    .X(_03203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__mux4_1 _26843_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net641),
    .S1(net647),
    .X(_03207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_66 ();
 sky130_fd_sc_hd__mux4_4 _26849_ (.A0(_03195_),
    .A1(_03200_),
    .A2(_03203_),
    .A3(_03207_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03213_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__mux4_1 _26852_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net639),
    .S1(\count16_2[1] ),
    .X(_03216_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__mux4_1 _26855_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net639),
    .S1(\count16_2[1] ),
    .X(_03219_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_60 ();
 sky130_fd_sc_hd__mux4_1 _26858_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net639),
    .S1(\count16_2[1] ),
    .X(_03222_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_58 ();
 sky130_fd_sc_hd__mux4_1 _26861_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net639),
    .S1(\count16_2[1] ),
    .X(_03225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_56 ();
 sky130_fd_sc_hd__mux4_1 _26864_ (.A0(_03216_),
    .A1(_03219_),
    .A2(_03222_),
    .A3(_03225_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03228_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_54 ();
 sky130_fd_sc_hd__mux2i_4 _26867_ (.A0(_03213_),
    .A1(_03228_),
    .S(\count16_2[5] ),
    .Y(_12008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_53 ();
 sky130_fd_sc_hd__mux4_1 _26869_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net601),
    .S1(net608),
    .X(_03232_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_51 ();
 sky130_fd_sc_hd__mux4_1 _26872_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net601),
    .S1(net608),
    .X(_03235_));
 sky130_fd_sc_hd__mux4_1 _26873_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net601),
    .S1(net608),
    .X(_03236_));
 sky130_fd_sc_hd__mux4_1 _26874_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net601),
    .S1(net608),
    .X(_03237_));
 sky130_fd_sc_hd__mux4_4 _26875_ (.A0(_03232_),
    .A1(_03235_),
    .A2(_03236_),
    .A3(_03237_),
    .S0(net597),
    .S1(net594),
    .X(_03238_));
 sky130_fd_sc_hd__mux4_1 _26876_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net600),
    .S1(net607),
    .X(_03239_));
 sky130_fd_sc_hd__mux4_1 _26877_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net599),
    .S1(net606),
    .X(_03240_));
 sky130_fd_sc_hd__mux4_1 _26878_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net599),
    .S1(net606),
    .X(_03241_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_49 ();
 sky130_fd_sc_hd__mux4_1 _26881_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net599),
    .S1(net606),
    .X(_03244_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_48 ();
 sky130_fd_sc_hd__mux4_1 _26883_ (.A0(_03239_),
    .A1(_03240_),
    .A2(_03241_),
    .A3(_03244_),
    .S0(net598),
    .S1(net594),
    .X(_03246_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__mux2i_4 _26885_ (.A0(_03238_),
    .A1(_03246_),
    .S(net592),
    .Y(_03248_));
 sky130_fd_sc_hd__mux4_1 _26886_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net602),
    .S1(net605),
    .X(_03249_));
 sky130_fd_sc_hd__mux4_1 _26887_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net602),
    .S1(net605),
    .X(_03250_));
 sky130_fd_sc_hd__mux4_1 _26888_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net602),
    .S1(net605),
    .X(_03251_));
 sky130_fd_sc_hd__mux4_1 _26889_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net602),
    .S1(net605),
    .X(_03252_));
 sky130_fd_sc_hd__mux4_4 _26890_ (.A0(_03249_),
    .A1(_03250_),
    .A2(_03251_),
    .A3(_03252_),
    .S0(net596),
    .S1(\count2_2[4] ),
    .X(_03253_));
 sky130_fd_sc_hd__mux4_1 _26891_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net603),
    .S1(net609),
    .X(_03254_));
 sky130_fd_sc_hd__mux4_1 _26892_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net603),
    .S1(net609),
    .X(_03255_));
 sky130_fd_sc_hd__mux4_1 _26893_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net603),
    .S1(net609),
    .X(_03256_));
 sky130_fd_sc_hd__mux4_1 _26894_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net603),
    .S1(net609),
    .X(_03257_));
 sky130_fd_sc_hd__mux4_1 _26895_ (.A0(_03254_),
    .A1(_03255_),
    .A2(_03256_),
    .A3(_03257_),
    .S0(net596),
    .S1(net595),
    .X(_03258_));
 sky130_fd_sc_hd__mux2i_4 _26896_ (.A0(_03253_),
    .A1(_03258_),
    .S(net593),
    .Y(_03259_));
 sky130_fd_sc_hd__xnor2_1 _26897_ (.A(_03248_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__xnor2_1 _26898_ (.A(_02910_),
    .B(_03260_),
    .Y(_12013_));
 sky130_fd_sc_hd__mux4_1 _26899_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03261_));
 sky130_fd_sc_hd__mux4_1 _26900_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03262_));
 sky130_fd_sc_hd__mux4_1 _26901_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03263_));
 sky130_fd_sc_hd__mux4_1 _26902_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03264_));
 sky130_fd_sc_hd__mux4_4 _26903_ (.A0(_03261_),
    .A1(_03262_),
    .A2(_03263_),
    .A3(_03264_),
    .S0(net669),
    .S1(net667),
    .X(_03265_));
 sky130_fd_sc_hd__mux4_1 _26904_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03266_));
 sky130_fd_sc_hd__mux4_1 _26905_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03267_));
 sky130_fd_sc_hd__mux4_1 _26906_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03268_));
 sky130_fd_sc_hd__mux4_1 _26907_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net674),
    .S1(net678),
    .X(_03269_));
 sky130_fd_sc_hd__mux4_1 _26908_ (.A0(_03266_),
    .A1(_03267_),
    .A2(_03268_),
    .A3(_03269_),
    .S0(net669),
    .S1(net667),
    .X(_03270_));
 sky130_fd_sc_hd__mux2i_4 _26909_ (.A0(_03265_),
    .A1(_03270_),
    .S(net666),
    .Y(_03271_));
 sky130_fd_sc_hd__mux4_1 _26910_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03272_));
 sky130_fd_sc_hd__mux4_1 _26911_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03273_));
 sky130_fd_sc_hd__mux4_1 _26912_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03274_));
 sky130_fd_sc_hd__mux4_1 _26913_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03275_));
 sky130_fd_sc_hd__mux4_4 _26914_ (.A0(_03272_),
    .A1(_03273_),
    .A2(_03274_),
    .A3(_03275_),
    .S0(net670),
    .S1(net668),
    .X(_03276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_45 ();
 sky130_fd_sc_hd__mux4_1 _26917_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03279_));
 sky130_fd_sc_hd__mux4_1 _26918_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03280_));
 sky130_fd_sc_hd__mux4_1 _26919_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03281_));
 sky130_fd_sc_hd__mux4_1 _26920_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net675),
    .S1(net681),
    .X(_03282_));
 sky130_fd_sc_hd__mux4_1 _26921_ (.A0(_03279_),
    .A1(_03280_),
    .A2(_03281_),
    .A3(_03282_),
    .S0(net670),
    .S1(net668),
    .X(_03283_));
 sky130_fd_sc_hd__mux2i_4 _26922_ (.A0(_03276_),
    .A1(_03283_),
    .S(\count15_2[5] ),
    .Y(_03284_));
 sky130_fd_sc_hd__mux4_1 _26923_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03285_));
 sky130_fd_sc_hd__mux4_1 _26924_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03286_));
 sky130_fd_sc_hd__mux4_1 _26925_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03287_));
 sky130_fd_sc_hd__mux4_1 _26926_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03288_));
 sky130_fd_sc_hd__mux4_4 _26927_ (.A0(_03285_),
    .A1(_03286_),
    .A2(_03287_),
    .A3(_03288_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03289_));
 sky130_fd_sc_hd__mux4_1 _26928_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03290_));
 sky130_fd_sc_hd__mux4_1 _26929_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03291_));
 sky130_fd_sc_hd__mux4_1 _26930_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net674),
    .S1(\count15_2[1] ),
    .X(_03292_));
 sky130_fd_sc_hd__mux4_1 _26931_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net674),
    .S1(\count15_2[1] ),
    .X(_03293_));
 sky130_fd_sc_hd__mux4_1 _26932_ (.A0(_03290_),
    .A1(_03291_),
    .A2(_03292_),
    .A3(_03293_),
    .S0(net669),
    .S1(net667),
    .X(_03294_));
 sky130_fd_sc_hd__mux2i_4 _26933_ (.A0(_03289_),
    .A1(_03294_),
    .S(net666),
    .Y(_03295_));
 sky130_fd_sc_hd__xnor2_1 _26934_ (.A(_03284_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__xnor2_2 _26935_ (.A(_03271_),
    .B(_03296_),
    .Y(_12012_));
 sky130_fd_sc_hd__mux4_1 _26936_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net560),
    .S1(net570),
    .X(_03297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_44 ();
 sky130_fd_sc_hd__mux4_1 _26938_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net560),
    .S1(net570),
    .X(_03299_));
 sky130_fd_sc_hd__mux4_1 _26939_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net560),
    .S1(net570),
    .X(_03300_));
 sky130_fd_sc_hd__mux4_1 _26940_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net560),
    .S1(net570),
    .X(_03301_));
 sky130_fd_sc_hd__mux4_2 _26941_ (.A0(_03297_),
    .A1(_03299_),
    .A2(_03300_),
    .A3(_03301_),
    .S0(net557),
    .S1(net555),
    .X(_03302_));
 sky130_fd_sc_hd__mux4_1 _26942_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net565),
    .S1(net569),
    .X(_03303_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__mux4_1 _26944_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net565),
    .S1(net569),
    .X(_03305_));
 sky130_fd_sc_hd__mux4_1 _26945_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net565),
    .S1(net569),
    .X(_03306_));
 sky130_fd_sc_hd__mux4_1 _26946_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net565),
    .S1(net569),
    .X(_03307_));
 sky130_fd_sc_hd__mux4_1 _26947_ (.A0(_03303_),
    .A1(_03305_),
    .A2(_03306_),
    .A3(_03307_),
    .S0(net557),
    .S1(net555),
    .X(_03308_));
 sky130_fd_sc_hd__mux2i_4 _26948_ (.A0(_03302_),
    .A1(_03308_),
    .S(net553),
    .Y(_12011_));
 sky130_fd_sc_hd__mux4_1 _26949_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03309_));
 sky130_fd_sc_hd__mux4_1 _26950_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03310_));
 sky130_fd_sc_hd__mux4_1 _26951_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03311_));
 sky130_fd_sc_hd__mux4_1 _26952_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03312_));
 sky130_fd_sc_hd__mux4_4 _26953_ (.A0(_03309_),
    .A1(_03310_),
    .A2(_03311_),
    .A3(_03312_),
    .S0(net633),
    .S1(net631),
    .X(_03313_));
 sky130_fd_sc_hd__mux4_1 _26954_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03314_));
 sky130_fd_sc_hd__mux4_1 _26955_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03315_));
 sky130_fd_sc_hd__mux4_1 _26956_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03316_));
 sky130_fd_sc_hd__mux4_1 _26957_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net637),
    .S1(net643),
    .X(_03317_));
 sky130_fd_sc_hd__mux4_1 _26958_ (.A0(_03314_),
    .A1(_03315_),
    .A2(_03316_),
    .A3(_03317_),
    .S0(net633),
    .S1(net631),
    .X(_03318_));
 sky130_fd_sc_hd__mux2i_4 _26959_ (.A0(_03313_),
    .A1(_03318_),
    .S(net629),
    .Y(_12016_));
 sky130_fd_sc_hd__mux4_1 _26960_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net604),
    .S1(net609),
    .X(_03319_));
 sky130_fd_sc_hd__mux4_1 _26961_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net604),
    .S1(net609),
    .X(_03320_));
 sky130_fd_sc_hd__mux4_1 _26962_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net604),
    .S1(net609),
    .X(_03321_));
 sky130_fd_sc_hd__mux4_1 _26963_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net604),
    .S1(net609),
    .X(_03322_));
 sky130_fd_sc_hd__mux4_4 _26964_ (.A0(_03319_),
    .A1(_03320_),
    .A2(_03321_),
    .A3(_03322_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03323_));
 sky130_fd_sc_hd__mux4_1 _26965_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net604),
    .S1(net609),
    .X(_03324_));
 sky130_fd_sc_hd__mux4_1 _26966_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net604),
    .S1(net609),
    .X(_03325_));
 sky130_fd_sc_hd__mux4_1 _26967_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net602),
    .S1(net609),
    .X(_03326_));
 sky130_fd_sc_hd__mux4_1 _26968_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net602),
    .S1(net609),
    .X(_03327_));
 sky130_fd_sc_hd__mux4_1 _26969_ (.A0(_03324_),
    .A1(_03325_),
    .A2(_03326_),
    .A3(_03327_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03328_));
 sky130_fd_sc_hd__mux2i_4 _26970_ (.A0(_03323_),
    .A1(_03328_),
    .S(net593),
    .Y(_03329_));
 sky130_fd_sc_hd__mux4_1 _26971_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net604),
    .S1(net609),
    .X(_03330_));
 sky130_fd_sc_hd__mux4_1 _26972_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net604),
    .S1(net609),
    .X(_03331_));
 sky130_fd_sc_hd__mux4_1 _26973_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net604),
    .S1(net609),
    .X(_03332_));
 sky130_fd_sc_hd__mux4_1 _26974_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net604),
    .S1(net609),
    .X(_03333_));
 sky130_fd_sc_hd__mux4_4 _26975_ (.A0(_03330_),
    .A1(_03331_),
    .A2(_03332_),
    .A3(_03333_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03334_));
 sky130_fd_sc_hd__mux4_1 _26976_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net602),
    .S1(net609),
    .X(_03335_));
 sky130_fd_sc_hd__mux4_1 _26977_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net602),
    .S1(net609),
    .X(_03336_));
 sky130_fd_sc_hd__mux4_1 _26978_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net602),
    .S1(net609),
    .X(_03337_));
 sky130_fd_sc_hd__mux4_1 _26979_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net602),
    .S1(net609),
    .X(_03338_));
 sky130_fd_sc_hd__mux4_1 _26980_ (.A0(_03335_),
    .A1(_03336_),
    .A2(_03337_),
    .A3(_03338_),
    .S0(net596),
    .S1(\count2_2[4] ),
    .X(_03339_));
 sky130_fd_sc_hd__mux2i_4 _26981_ (.A0(_03334_),
    .A1(_03339_),
    .S(net593),
    .Y(_03340_));
 sky130_fd_sc_hd__xnor2_1 _26982_ (.A(_03329_),
    .B(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__xnor2_1 _26983_ (.A(_03124_),
    .B(_03341_),
    .Y(_12024_));
 sky130_fd_sc_hd__mux4_1 _26984_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net673),
    .S1(net680),
    .X(_03342_));
 sky130_fd_sc_hd__mux4_1 _26985_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net673),
    .S1(net680),
    .X(_03343_));
 sky130_fd_sc_hd__mux4_1 _26986_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net673),
    .S1(net680),
    .X(_03344_));
 sky130_fd_sc_hd__mux4_1 _26987_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net673),
    .S1(net680),
    .X(_03345_));
 sky130_fd_sc_hd__mux4_4 _26988_ (.A0(_03342_),
    .A1(_03343_),
    .A2(_03344_),
    .A3(_03345_),
    .S0(net669),
    .S1(net667),
    .X(_03346_));
 sky130_fd_sc_hd__mux4_1 _26989_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__mux4_1 _26991_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03349_));
 sky130_fd_sc_hd__mux4_1 _26992_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03350_));
 sky130_fd_sc_hd__mux4_1 _26993_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03351_));
 sky130_fd_sc_hd__mux4_1 _26994_ (.A0(_03347_),
    .A1(_03349_),
    .A2(_03350_),
    .A3(_03351_),
    .S0(net669),
    .S1(net667),
    .X(_03352_));
 sky130_fd_sc_hd__mux2i_4 _26995_ (.A0(_03346_),
    .A1(_03352_),
    .S(net666),
    .Y(_03353_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_40 ();
 sky130_fd_sc_hd__mux4_1 _26998_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03356_));
 sky130_fd_sc_hd__mux4_1 _26999_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03357_));
 sky130_fd_sc_hd__mux4_1 _27000_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03358_));
 sky130_fd_sc_hd__mux4_1 _27001_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03359_));
 sky130_fd_sc_hd__mux4_4 _27002_ (.A0(_03356_),
    .A1(_03357_),
    .A2(_03358_),
    .A3(_03359_),
    .S0(net669),
    .S1(net667),
    .X(_03360_));
 sky130_fd_sc_hd__mux4_1 _27003_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03361_));
 sky130_fd_sc_hd__mux4_1 _27004_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03362_));
 sky130_fd_sc_hd__mux4_1 _27005_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03363_));
 sky130_fd_sc_hd__mux4_1 _27006_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net674),
    .S1(net678),
    .X(_03364_));
 sky130_fd_sc_hd__mux4_1 _27007_ (.A0(_03361_),
    .A1(_03362_),
    .A2(_03363_),
    .A3(_03364_),
    .S0(net669),
    .S1(net667),
    .X(_03365_));
 sky130_fd_sc_hd__mux2i_4 _27008_ (.A0(_03360_),
    .A1(_03365_),
    .S(net666),
    .Y(_03366_));
 sky130_fd_sc_hd__mux4_1 _27009_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net676),
    .S1(net682),
    .X(_03367_));
 sky130_fd_sc_hd__mux4_1 _27010_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net676),
    .S1(net682),
    .X(_03368_));
 sky130_fd_sc_hd__mux4_1 _27011_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net676),
    .S1(net682),
    .X(_03369_));
 sky130_fd_sc_hd__mux4_1 _27012_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net676),
    .S1(net682),
    .X(_03370_));
 sky130_fd_sc_hd__mux4_4 _27013_ (.A0(_03367_),
    .A1(_03368_),
    .A2(_03369_),
    .A3(_03370_),
    .S0(net670),
    .S1(net668),
    .X(_03371_));
 sky130_fd_sc_hd__mux4_1 _27014_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net677),
    .S1(net682),
    .X(_03372_));
 sky130_fd_sc_hd__mux4_1 _27015_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net677),
    .S1(net682),
    .X(_03373_));
 sky130_fd_sc_hd__mux4_1 _27016_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net677),
    .S1(net682),
    .X(_03374_));
 sky130_fd_sc_hd__mux4_1 _27017_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net677),
    .S1(net682),
    .X(_03375_));
 sky130_fd_sc_hd__mux4_1 _27018_ (.A0(_03372_),
    .A1(_03373_),
    .A2(_03374_),
    .A3(_03375_),
    .S0(net670),
    .S1(net668),
    .X(_03376_));
 sky130_fd_sc_hd__mux2i_4 _27019_ (.A0(_03371_),
    .A1(_03376_),
    .S(\count15_2[5] ),
    .Y(_03377_));
 sky130_fd_sc_hd__xnor2_1 _27020_ (.A(_03366_),
    .B(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__xnor2_1 _27021_ (.A(_03353_),
    .B(_03378_),
    .Y(_12023_));
 sky130_fd_sc_hd__mux4_1 _27022_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net560),
    .S1(net570),
    .X(_03379_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__mux4_1 _27024_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net560),
    .S1(net570),
    .X(_03381_));
 sky130_fd_sc_hd__mux4_1 _27025_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net560),
    .S1(net570),
    .X(_03382_));
 sky130_fd_sc_hd__mux4_1 _27026_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net560),
    .S1(net570),
    .X(_03383_));
 sky130_fd_sc_hd__mux4_2 _27027_ (.A0(_03379_),
    .A1(_03381_),
    .A2(_03382_),
    .A3(_03383_),
    .S0(net557),
    .S1(net555),
    .X(_03384_));
 sky130_fd_sc_hd__mux4_1 _27028_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net560),
    .S1(net570),
    .X(_03385_));
 sky130_fd_sc_hd__mux4_1 _27029_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net560),
    .S1(net569),
    .X(_03386_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__mux4_1 _27031_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net566),
    .S1(net571),
    .X(_03388_));
 sky130_fd_sc_hd__mux4_1 _27032_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net566),
    .S1(net571),
    .X(_03389_));
 sky130_fd_sc_hd__mux4_1 _27033_ (.A0(_03385_),
    .A1(_03386_),
    .A2(_03388_),
    .A3(_03389_),
    .S0(net557),
    .S1(net555),
    .X(_03390_));
 sky130_fd_sc_hd__mux2i_4 _27034_ (.A0(_03384_),
    .A1(_03390_),
    .S(net553),
    .Y(_12022_));
 sky130_fd_sc_hd__mux4_1 _27035_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net641),
    .S1(net646),
    .X(_03391_));
 sky130_fd_sc_hd__mux4_1 _27036_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net641),
    .S1(net647),
    .X(_03392_));
 sky130_fd_sc_hd__mux4_1 _27037_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net641),
    .S1(net647),
    .X(_03393_));
 sky130_fd_sc_hd__mux4_1 _27038_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net641),
    .S1(net647),
    .X(_03394_));
 sky130_fd_sc_hd__mux4_4 _27039_ (.A0(_03391_),
    .A1(_03392_),
    .A2(_03393_),
    .A3(_03394_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03395_));
 sky130_fd_sc_hd__mux4_1 _27040_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net639),
    .S1(\count16_2[1] ),
    .X(_03396_));
 sky130_fd_sc_hd__mux4_1 _27041_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net638),
    .S1(\count16_2[1] ),
    .X(_03397_));
 sky130_fd_sc_hd__mux4_1 _27042_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net639),
    .S1(\count16_2[1] ),
    .X(_03398_));
 sky130_fd_sc_hd__mux4_1 _27043_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net639),
    .S1(\count16_2[1] ),
    .X(_03399_));
 sky130_fd_sc_hd__mux4_1 _27044_ (.A0(_03396_),
    .A1(_03397_),
    .A2(_03398_),
    .A3(_03399_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03400_));
 sky130_fd_sc_hd__mux2i_2 _27045_ (.A0(_03395_),
    .A1(_03400_),
    .S(\count16_2[5] ),
    .Y(_12027_));
 sky130_fd_sc_hd__mux4_1 _27046_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net603),
    .S1(net607),
    .X(_03401_));
 sky130_fd_sc_hd__mux4_1 _27047_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net603),
    .S1(net606),
    .X(_03402_));
 sky130_fd_sc_hd__mux4_1 _27048_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net603),
    .S1(net607),
    .X(_03403_));
 sky130_fd_sc_hd__mux4_1 _27049_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net603),
    .S1(net607),
    .X(_03404_));
 sky130_fd_sc_hd__mux4_4 _27050_ (.A0(_03401_),
    .A1(_03402_),
    .A2(_03403_),
    .A3(_03404_),
    .S0(net596),
    .S1(net595),
    .X(_03405_));
 sky130_fd_sc_hd__mux4_1 _27051_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net600),
    .S1(net607),
    .X(_03406_));
 sky130_fd_sc_hd__mux4_1 _27052_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net600),
    .S1(net605),
    .X(_03407_));
 sky130_fd_sc_hd__mux4_1 _27053_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net600),
    .S1(net607),
    .X(_03408_));
 sky130_fd_sc_hd__mux4_1 _27054_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net600),
    .S1(net607),
    .X(_03409_));
 sky130_fd_sc_hd__mux4_1 _27055_ (.A0(_03406_),
    .A1(_03407_),
    .A2(_03408_),
    .A3(_03409_),
    .S0(net596),
    .S1(net595),
    .X(_03410_));
 sky130_fd_sc_hd__mux2i_4 _27056_ (.A0(_03405_),
    .A1(_03410_),
    .S(net593),
    .Y(_03411_));
 sky130_fd_sc_hd__mux4_1 _27057_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net601),
    .S1(net608),
    .X(_03412_));
 sky130_fd_sc_hd__mux4_1 _27058_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net601),
    .S1(net608),
    .X(_03413_));
 sky130_fd_sc_hd__mux4_1 _27059_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net601),
    .S1(net608),
    .X(_03414_));
 sky130_fd_sc_hd__mux4_1 _27060_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net601),
    .S1(net608),
    .X(_03415_));
 sky130_fd_sc_hd__mux4_2 _27061_ (.A0(_03412_),
    .A1(_03413_),
    .A2(_03414_),
    .A3(_03415_),
    .S0(net597),
    .S1(net594),
    .X(_03416_));
 sky130_fd_sc_hd__mux4_1 _27062_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03417_));
 sky130_fd_sc_hd__mux4_1 _27063_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03418_));
 sky130_fd_sc_hd__mux4_1 _27064_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03419_));
 sky130_fd_sc_hd__mux4_1 _27065_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03420_));
 sky130_fd_sc_hd__mux4_1 _27066_ (.A0(_03417_),
    .A1(_03418_),
    .A2(_03419_),
    .A3(_03420_),
    .S0(net597),
    .S1(net594),
    .X(_03421_));
 sky130_fd_sc_hd__mux2i_4 _27067_ (.A0(_03416_),
    .A1(_03421_),
    .S(net592),
    .Y(_03422_));
 sky130_fd_sc_hd__xnor2_1 _27068_ (.A(_03411_),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__xnor2_1 _27069_ (.A(_03259_),
    .B(_03423_),
    .Y(_12032_));
 sky130_fd_sc_hd__mux4_1 _27070_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03424_));
 sky130_fd_sc_hd__mux4_1 _27071_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03425_));
 sky130_fd_sc_hd__mux4_1 _27072_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03426_));
 sky130_fd_sc_hd__mux4_1 _27073_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03427_));
 sky130_fd_sc_hd__mux4_2 _27074_ (.A0(_03424_),
    .A1(_03425_),
    .A2(_03426_),
    .A3(_03427_),
    .S0(net669),
    .S1(net667),
    .X(_03428_));
 sky130_fd_sc_hd__mux4_1 _27075_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__mux4_1 _27077_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03431_));
 sky130_fd_sc_hd__mux4_1 _27078_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03432_));
 sky130_fd_sc_hd__mux4_1 _27079_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net673),
    .S1(net680),
    .X(_03433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__mux4_1 _27081_ (.A0(_03429_),
    .A1(_03431_),
    .A2(_03432_),
    .A3(_03433_),
    .S0(net669),
    .S1(net667),
    .X(_03435_));
 sky130_fd_sc_hd__mux2i_4 _27082_ (.A0(_03428_),
    .A1(_03435_),
    .S(net666),
    .Y(_03436_));
 sky130_fd_sc_hd__mux4_1 _27083_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03437_));
 sky130_fd_sc_hd__mux4_1 _27084_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03438_));
 sky130_fd_sc_hd__mux4_1 _27085_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03439_));
 sky130_fd_sc_hd__mux4_1 _27086_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03440_));
 sky130_fd_sc_hd__mux4_4 _27087_ (.A0(_03437_),
    .A1(_03438_),
    .A2(_03439_),
    .A3(_03440_),
    .S0(net669),
    .S1(net667),
    .X(_03441_));
 sky130_fd_sc_hd__mux4_1 _27088_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03442_));
 sky130_fd_sc_hd__mux4_1 _27089_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03443_));
 sky130_fd_sc_hd__mux4_1 _27090_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03444_));
 sky130_fd_sc_hd__mux4_1 _27091_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net672),
    .S1(net679),
    .X(_03445_));
 sky130_fd_sc_hd__mux4_1 _27092_ (.A0(_03442_),
    .A1(_03443_),
    .A2(_03444_),
    .A3(_03445_),
    .S0(net671),
    .S1(net668),
    .X(_03446_));
 sky130_fd_sc_hd__mux2i_4 _27093_ (.A0(_03441_),
    .A1(_03446_),
    .S(net665),
    .Y(_03447_));
 sky130_fd_sc_hd__xnor2_1 _27094_ (.A(_03436_),
    .B(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__xnor2_2 _27095_ (.A(_03024_),
    .B(_03448_),
    .Y(_12031_));
 sky130_fd_sc_hd__mux4_1 _27096_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03449_));
 sky130_fd_sc_hd__mux4_1 _27097_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03450_));
 sky130_fd_sc_hd__mux4_1 _27098_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03451_));
 sky130_fd_sc_hd__mux4_1 _27099_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03452_));
 sky130_fd_sc_hd__mux4_2 _27100_ (.A0(_03449_),
    .A1(_03450_),
    .A2(_03451_),
    .A3(_03452_),
    .S0(net559),
    .S1(net555),
    .X(_03453_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__mux4_1 _27102_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03455_));
 sky130_fd_sc_hd__mux4_1 _27103_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03456_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__mux4_1 _27105_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03458_));
 sky130_fd_sc_hd__mux4_1 _27106_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net561),
    .S1(net572),
    .X(_03459_));
 sky130_fd_sc_hd__mux4_1 _27107_ (.A0(_03455_),
    .A1(_03456_),
    .A2(_03458_),
    .A3(_03459_),
    .S0(net559),
    .S1(net555),
    .X(_03460_));
 sky130_fd_sc_hd__mux2i_4 _27108_ (.A0(_03453_),
    .A1(_03460_),
    .S(net553),
    .Y(_12030_));
 sky130_fd_sc_hd__mux4_1 _27109_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net641),
    .S1(\count16_2[1] ),
    .X(_03461_));
 sky130_fd_sc_hd__mux4_1 _27110_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net641),
    .S1(\count16_2[1] ),
    .X(_03462_));
 sky130_fd_sc_hd__mux4_1 _27111_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net641),
    .S1(net642),
    .X(_03463_));
 sky130_fd_sc_hd__mux4_1 _27112_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net641),
    .S1(\count16_2[1] ),
    .X(_03464_));
 sky130_fd_sc_hd__mux4_4 _27113_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03465_));
 sky130_fd_sc_hd__mux4_1 _27114_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net641),
    .S1(net642),
    .X(_03466_));
 sky130_fd_sc_hd__mux4_1 _27115_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net641),
    .S1(net642),
    .X(_03467_));
 sky130_fd_sc_hd__mux4_1 _27116_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net641),
    .S1(net642),
    .X(_03468_));
 sky130_fd_sc_hd__mux4_1 _27117_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net641),
    .S1(net642),
    .X(_03469_));
 sky130_fd_sc_hd__mux4_1 _27118_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03470_));
 sky130_fd_sc_hd__mux2i_4 _27119_ (.A0(_03465_),
    .A1(_03470_),
    .S(\count16_2[5] ),
    .Y(_12035_));
 sky130_fd_sc_hd__mux4_1 _27120_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net601),
    .S1(net608),
    .X(_03471_));
 sky130_fd_sc_hd__mux4_1 _27121_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net601),
    .S1(net608),
    .X(_03472_));
 sky130_fd_sc_hd__mux4_1 _27122_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net601),
    .S1(net608),
    .X(_03473_));
 sky130_fd_sc_hd__mux4_1 _27123_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net601),
    .S1(net608),
    .X(_03474_));
 sky130_fd_sc_hd__mux4_2 _27124_ (.A0(_03471_),
    .A1(_03472_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(net597),
    .S1(net594),
    .X(_03475_));
 sky130_fd_sc_hd__mux4_1 _27125_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net599),
    .S1(net606),
    .X(_03476_));
 sky130_fd_sc_hd__mux4_1 _27126_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03477_));
 sky130_fd_sc_hd__mux4_1 _27127_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03478_));
 sky130_fd_sc_hd__mux4_1 _27128_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03479_));
 sky130_fd_sc_hd__mux4_1 _27129_ (.A0(_03476_),
    .A1(_03477_),
    .A2(_03478_),
    .A3(_03479_),
    .S0(net597),
    .S1(net594),
    .X(_03480_));
 sky130_fd_sc_hd__mux2i_4 _27130_ (.A0(_03475_),
    .A1(_03480_),
    .S(net592),
    .Y(_03481_));
 sky130_fd_sc_hd__mux4_1 _27131_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net601),
    .S1(net608),
    .X(_03482_));
 sky130_fd_sc_hd__mux4_1 _27132_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net601),
    .S1(net608),
    .X(_03483_));
 sky130_fd_sc_hd__mux4_1 _27133_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net601),
    .S1(net608),
    .X(_03484_));
 sky130_fd_sc_hd__mux4_1 _27134_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net601),
    .S1(net608),
    .X(_03485_));
 sky130_fd_sc_hd__mux4_4 _27135_ (.A0(_03482_),
    .A1(_03483_),
    .A2(_03484_),
    .A3(_03485_),
    .S0(net597),
    .S1(net594),
    .X(_03486_));
 sky130_fd_sc_hd__mux4_1 _27136_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net599),
    .S1(net606),
    .X(_03487_));
 sky130_fd_sc_hd__mux4_1 _27137_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net599),
    .S1(net606),
    .X(_03488_));
 sky130_fd_sc_hd__mux4_1 _27138_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net599),
    .S1(net606),
    .X(_03489_));
 sky130_fd_sc_hd__mux4_1 _27139_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net599),
    .S1(net606),
    .X(_03490_));
 sky130_fd_sc_hd__mux4_1 _27140_ (.A0(_03487_),
    .A1(_03488_),
    .A2(_03489_),
    .A3(_03490_),
    .S0(net597),
    .S1(net594),
    .X(_03491_));
 sky130_fd_sc_hd__mux2i_4 _27141_ (.A0(_03486_),
    .A1(_03491_),
    .S(net592),
    .Y(_03492_));
 sky130_fd_sc_hd__xnor2_1 _27142_ (.A(_03481_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__xnor2_1 _27143_ (.A(_03340_),
    .B(_03493_),
    .Y(_12040_));
 sky130_fd_sc_hd__mux4_1 _27144_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net674),
    .S1(net680),
    .X(_03494_));
 sky130_fd_sc_hd__mux4_1 _27145_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net674),
    .S1(net680),
    .X(_03495_));
 sky130_fd_sc_hd__mux4_1 _27146_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net674),
    .S1(net680),
    .X(_03496_));
 sky130_fd_sc_hd__mux4_1 _27147_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net674),
    .S1(net680),
    .X(_03497_));
 sky130_fd_sc_hd__mux4_4 _27148_ (.A0(_03494_),
    .A1(_03495_),
    .A2(_03496_),
    .A3(_03497_),
    .S0(net669),
    .S1(net667),
    .X(_03498_));
 sky130_fd_sc_hd__mux4_1 _27149_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net673),
    .S1(net680),
    .X(_03499_));
 sky130_fd_sc_hd__mux4_1 _27150_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03500_));
 sky130_fd_sc_hd__mux4_1 _27151_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03501_));
 sky130_fd_sc_hd__mux4_1 _27152_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net673),
    .S1(\count15_2[1] ),
    .X(_03502_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__mux4_1 _27154_ (.A0(_03499_),
    .A1(_03500_),
    .A2(_03501_),
    .A3(_03502_),
    .S0(net669),
    .S1(net667),
    .X(_03504_));
 sky130_fd_sc_hd__mux2i_4 _27155_ (.A0(_03498_),
    .A1(_03504_),
    .S(net666),
    .Y(_03505_));
 sky130_fd_sc_hd__mux4_1 _27156_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03506_));
 sky130_fd_sc_hd__mux4_1 _27157_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03507_));
 sky130_fd_sc_hd__mux4_1 _27158_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03508_));
 sky130_fd_sc_hd__mux4_1 _27159_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03509_));
 sky130_fd_sc_hd__mux4_4 _27160_ (.A0(_03506_),
    .A1(_03507_),
    .A2(_03508_),
    .A3(_03509_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03510_));
 sky130_fd_sc_hd__mux4_1 _27161_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net677),
    .S1(net682),
    .X(_03511_));
 sky130_fd_sc_hd__mux4_1 _27162_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net677),
    .S1(net682),
    .X(_03512_));
 sky130_fd_sc_hd__mux4_1 _27163_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net677),
    .S1(net682),
    .X(_03513_));
 sky130_fd_sc_hd__mux4_1 _27164_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net677),
    .S1(net682),
    .X(_03514_));
 sky130_fd_sc_hd__mux4_1 _27165_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(net671),
    .S1(\count15_2[4] ),
    .X(_03515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__mux2i_4 _27167_ (.A0(_03510_),
    .A1(_03515_),
    .S(\count15_2[5] ),
    .Y(_03517_));
 sky130_fd_sc_hd__xnor2_1 _27168_ (.A(_03505_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__xnor2_2 _27169_ (.A(_03163_),
    .B(_03518_),
    .Y(_12039_));
 sky130_fd_sc_hd__mux4_1 _27170_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03519_));
 sky130_fd_sc_hd__mux4_1 _27171_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03520_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__mux4_1 _27173_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03522_));
 sky130_fd_sc_hd__mux4_1 _27174_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03523_));
 sky130_fd_sc_hd__mux4_4 _27175_ (.A0(_03519_),
    .A1(_03520_),
    .A2(_03522_),
    .A3(_03523_),
    .S0(net559),
    .S1(\count7_2[4] ),
    .X(_03524_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__mux4_1 _27177_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03526_));
 sky130_fd_sc_hd__mux4_1 _27178_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03527_));
 sky130_fd_sc_hd__mux4_1 _27179_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03528_));
 sky130_fd_sc_hd__mux4_1 _27180_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net562),
    .S1(net567),
    .X(_03529_));
 sky130_fd_sc_hd__mux4_1 _27181_ (.A0(_03526_),
    .A1(_03527_),
    .A2(_03528_),
    .A3(_03529_),
    .S0(net559),
    .S1(net555),
    .X(_03530_));
 sky130_fd_sc_hd__mux2i_4 _27182_ (.A0(_03524_),
    .A1(_03530_),
    .S(net553),
    .Y(_12038_));
 sky130_fd_sc_hd__mux4_1 _27183_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net636),
    .S1(net646),
    .X(_03531_));
 sky130_fd_sc_hd__mux4_1 _27184_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net636),
    .S1(net647),
    .X(_03532_));
 sky130_fd_sc_hd__mux4_1 _27185_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net636),
    .S1(net646),
    .X(_03533_));
 sky130_fd_sc_hd__mux4_1 _27186_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net636),
    .S1(net646),
    .X(_03534_));
 sky130_fd_sc_hd__mux4_4 _27187_ (.A0(_03531_),
    .A1(_03532_),
    .A2(_03533_),
    .A3(_03534_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03535_));
 sky130_fd_sc_hd__mux4_1 _27188_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net639),
    .S1(net645),
    .X(_03536_));
 sky130_fd_sc_hd__mux4_1 _27189_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net639),
    .S1(net647),
    .X(_03537_));
 sky130_fd_sc_hd__mux4_1 _27190_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net636),
    .S1(net647),
    .X(_03538_));
 sky130_fd_sc_hd__mux4_1 _27191_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net639),
    .S1(net647),
    .X(_03539_));
 sky130_fd_sc_hd__mux4_1 _27192_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03540_));
 sky130_fd_sc_hd__mux2i_4 _27193_ (.A0(_03535_),
    .A1(_03540_),
    .S(\count16_2[5] ),
    .Y(_12043_));
 sky130_fd_sc_hd__mux4_1 _27194_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net601),
    .S1(net608),
    .X(_03541_));
 sky130_fd_sc_hd__mux4_1 _27195_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net601),
    .S1(net608),
    .X(_03542_));
 sky130_fd_sc_hd__mux4_1 _27196_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net601),
    .S1(net608),
    .X(_03543_));
 sky130_fd_sc_hd__mux4_1 _27197_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net601),
    .S1(net608),
    .X(_03544_));
 sky130_fd_sc_hd__mux4_4 _27198_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(net597),
    .S1(net594),
    .X(_03545_));
 sky130_fd_sc_hd__mux4_1 _27199_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03546_));
 sky130_fd_sc_hd__mux4_1 _27200_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03547_));
 sky130_fd_sc_hd__mux4_1 _27201_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03548_));
 sky130_fd_sc_hd__mux4_1 _27202_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net600),
    .S1(\count2_2[1] ),
    .X(_03549_));
 sky130_fd_sc_hd__mux4_1 _27203_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(net597),
    .S1(net594),
    .X(_03550_));
 sky130_fd_sc_hd__mux2i_4 _27204_ (.A0(_03545_),
    .A1(_03550_),
    .S(net592),
    .Y(_03551_));
 sky130_fd_sc_hd__mux4_1 _27205_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03552_));
 sky130_fd_sc_hd__mux4_1 _27206_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03553_));
 sky130_fd_sc_hd__mux4_1 _27207_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03554_));
 sky130_fd_sc_hd__mux4_1 _27208_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03555_));
 sky130_fd_sc_hd__mux4_4 _27209_ (.A0(_03552_),
    .A1(_03553_),
    .A2(_03554_),
    .A3(_03555_),
    .S0(net598),
    .S1(net594),
    .X(_03556_));
 sky130_fd_sc_hd__mux4_1 _27210_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03557_));
 sky130_fd_sc_hd__mux4_1 _27211_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03558_));
 sky130_fd_sc_hd__mux4_1 _27212_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03559_));
 sky130_fd_sc_hd__mux4_1 _27213_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net599),
    .S1(net606),
    .X(_03560_));
 sky130_fd_sc_hd__mux4_1 _27214_ (.A0(_03557_),
    .A1(_03558_),
    .A2(_03559_),
    .A3(_03560_),
    .S0(net598),
    .S1(net594),
    .X(_03561_));
 sky130_fd_sc_hd__mux2i_4 _27215_ (.A0(_03556_),
    .A1(_03561_),
    .S(net592),
    .Y(_03562_));
 sky130_fd_sc_hd__xnor2_1 _27216_ (.A(_03551_),
    .B(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__xnor2_1 _27217_ (.A(_03411_),
    .B(_03563_),
    .Y(_12048_));
 sky130_fd_sc_hd__mux4_1 _27218_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03564_));
 sky130_fd_sc_hd__mux4_1 _27219_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03565_));
 sky130_fd_sc_hd__mux4_1 _27220_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03566_));
 sky130_fd_sc_hd__mux4_1 _27221_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03567_));
 sky130_fd_sc_hd__mux4_4 _27222_ (.A0(_03564_),
    .A1(_03565_),
    .A2(_03566_),
    .A3(_03567_),
    .S0(net670),
    .S1(net668),
    .X(_03568_));
 sky130_fd_sc_hd__mux4_1 _27223_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03569_));
 sky130_fd_sc_hd__mux4_1 _27224_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03570_));
 sky130_fd_sc_hd__mux4_1 _27225_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03571_));
 sky130_fd_sc_hd__mux4_1 _27226_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net676),
    .S1(net682),
    .X(_03572_));
 sky130_fd_sc_hd__mux4_1 _27227_ (.A0(_03569_),
    .A1(_03570_),
    .A2(_03571_),
    .A3(_03572_),
    .S0(net670),
    .S1(net668),
    .X(_03573_));
 sky130_fd_sc_hd__mux2i_4 _27228_ (.A0(_03568_),
    .A1(_03573_),
    .S(\count15_2[5] ),
    .Y(_03574_));
 sky130_fd_sc_hd__mux4_1 _27229_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03575_));
 sky130_fd_sc_hd__mux4_1 _27230_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03576_));
 sky130_fd_sc_hd__mux4_1 _27231_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03577_));
 sky130_fd_sc_hd__mux4_1 _27232_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03578_));
 sky130_fd_sc_hd__mux4_2 _27233_ (.A0(_03575_),
    .A1(_03576_),
    .A2(_03577_),
    .A3(_03578_),
    .S0(net670),
    .S1(net668),
    .X(_03579_));
 sky130_fd_sc_hd__mux4_1 _27234_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03580_));
 sky130_fd_sc_hd__mux4_1 _27235_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03581_));
 sky130_fd_sc_hd__mux4_1 _27236_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03582_));
 sky130_fd_sc_hd__mux4_1 _27237_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net675),
    .S1(net681),
    .X(_03583_));
 sky130_fd_sc_hd__mux4_1 _27238_ (.A0(_03580_),
    .A1(_03581_),
    .A2(_03582_),
    .A3(_03583_),
    .S0(net670),
    .S1(net668),
    .X(_03584_));
 sky130_fd_sc_hd__mux2i_4 _27239_ (.A0(_03579_),
    .A1(_03584_),
    .S(\count15_2[5] ),
    .Y(_03585_));
 sky130_fd_sc_hd__xnor2_2 _27240_ (.A(_03574_),
    .B(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__xnor2_2 _27241_ (.A(_03295_),
    .B(_03586_),
    .Y(_12047_));
 sky130_fd_sc_hd__mux4_1 _27242_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03587_));
 sky130_fd_sc_hd__mux4_1 _27243_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03588_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__mux4_1 _27245_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03590_));
 sky130_fd_sc_hd__mux4_1 _27246_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03591_));
 sky130_fd_sc_hd__mux4_4 _27247_ (.A0(_03587_),
    .A1(_03588_),
    .A2(_03590_),
    .A3(_03591_),
    .S0(net559),
    .S1(\count7_2[4] ),
    .X(_03592_));
 sky130_fd_sc_hd__mux4_1 _27248_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03593_));
 sky130_fd_sc_hd__mux4_1 _27249_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03594_));
 sky130_fd_sc_hd__mux4_1 _27250_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03595_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__mux4_1 _27252_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net562),
    .S1(net567),
    .X(_03597_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__mux4_1 _27254_ (.A0(_03593_),
    .A1(_03594_),
    .A2(_03595_),
    .A3(_03597_),
    .S0(net559),
    .S1(net555),
    .X(_03599_));
 sky130_fd_sc_hd__mux2i_4 _27255_ (.A0(_03592_),
    .A1(_03599_),
    .S(net553),
    .Y(_12046_));
 sky130_fd_sc_hd__mux4_1 _27256_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net635),
    .S1(net643),
    .X(_03600_));
 sky130_fd_sc_hd__mux4_1 _27257_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net635),
    .S1(net643),
    .X(_03601_));
 sky130_fd_sc_hd__mux4_1 _27258_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net635),
    .S1(net643),
    .X(_03602_));
 sky130_fd_sc_hd__mux4_1 _27259_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net635),
    .S1(net643),
    .X(_03603_));
 sky130_fd_sc_hd__mux4_4 _27260_ (.A0(_03600_),
    .A1(_03601_),
    .A2(_03602_),
    .A3(_03603_),
    .S0(net634),
    .S1(net632),
    .X(_03604_));
 sky130_fd_sc_hd__mux4_1 _27261_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net638),
    .S1(net645),
    .X(_03605_));
 sky130_fd_sc_hd__mux4_1 _27262_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net638),
    .S1(net645),
    .X(_03606_));
 sky130_fd_sc_hd__mux4_1 _27263_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net638),
    .S1(net645),
    .X(_03607_));
 sky130_fd_sc_hd__mux4_1 _27264_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net638),
    .S1(net645),
    .X(_03608_));
 sky130_fd_sc_hd__mux4_1 _27265_ (.A0(_03605_),
    .A1(_03606_),
    .A2(_03607_),
    .A3(_03608_),
    .S0(net633),
    .S1(net632),
    .X(_03609_));
 sky130_fd_sc_hd__mux2i_4 _27266_ (.A0(_03604_),
    .A1(_03609_),
    .S(net629),
    .Y(_12051_));
 sky130_fd_sc_hd__mux4_1 _27267_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net603),
    .S1(net606),
    .X(_03610_));
 sky130_fd_sc_hd__mux4_1 _27268_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net603),
    .S1(net606),
    .X(_03611_));
 sky130_fd_sc_hd__mux4_1 _27269_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net603),
    .S1(net606),
    .X(_03612_));
 sky130_fd_sc_hd__mux4_1 _27270_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net603),
    .S1(net606),
    .X(_03613_));
 sky130_fd_sc_hd__mux4_4 _27271_ (.A0(_03610_),
    .A1(_03611_),
    .A2(_03612_),
    .A3(_03613_),
    .S0(net596),
    .S1(net595),
    .X(_03614_));
 sky130_fd_sc_hd__mux4_1 _27272_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net603),
    .S1(net607),
    .X(_03615_));
 sky130_fd_sc_hd__mux4_1 _27273_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net603),
    .S1(net607),
    .X(_03616_));
 sky130_fd_sc_hd__mux4_1 _27274_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net603),
    .S1(net607),
    .X(_03617_));
 sky130_fd_sc_hd__mux4_1 _27275_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net603),
    .S1(net607),
    .X(_03618_));
 sky130_fd_sc_hd__mux4_1 _27276_ (.A0(_03615_),
    .A1(_03616_),
    .A2(_03617_),
    .A3(_03618_),
    .S0(net598),
    .S1(net595),
    .X(_03619_));
 sky130_fd_sc_hd__mux2i_4 _27277_ (.A0(_03614_),
    .A1(_03619_),
    .S(net592),
    .Y(_03620_));
 sky130_fd_sc_hd__xnor2_1 _27278_ (.A(_03492_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__xnor2_1 _27279_ (.A(_02959_),
    .B(_03621_),
    .Y(_12056_));
 sky130_fd_sc_hd__mux4_1 _27280_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net672),
    .S1(net679),
    .X(_03622_));
 sky130_fd_sc_hd__mux4_1 _27281_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net672),
    .S1(net679),
    .X(_03623_));
 sky130_fd_sc_hd__mux4_1 _27282_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net672),
    .S1(net679),
    .X(_03624_));
 sky130_fd_sc_hd__mux4_1 _27283_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net672),
    .S1(net679),
    .X(_03625_));
 sky130_fd_sc_hd__mux4_4 _27284_ (.A0(_03622_),
    .A1(_03623_),
    .A2(_03624_),
    .A3(_03625_),
    .S0(net669),
    .S1(net667),
    .X(_03626_));
 sky130_fd_sc_hd__mux4_1 _27285_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net677),
    .S1(net681),
    .X(_03627_));
 sky130_fd_sc_hd__mux4_1 _27286_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net677),
    .S1(net681),
    .X(_03628_));
 sky130_fd_sc_hd__mux4_1 _27287_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net677),
    .S1(net681),
    .X(_03629_));
 sky130_fd_sc_hd__mux4_1 _27288_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net677),
    .S1(net681),
    .X(_03630_));
 sky130_fd_sc_hd__mux4_1 _27289_ (.A0(_03627_),
    .A1(_03628_),
    .A2(_03629_),
    .A3(_03630_),
    .S0(net671),
    .S1(net668),
    .X(_03631_));
 sky130_fd_sc_hd__mux2i_4 _27290_ (.A0(_03626_),
    .A1(_03631_),
    .S(net665),
    .Y(_03632_));
 sky130_fd_sc_hd__mux4_1 _27291_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03633_));
 sky130_fd_sc_hd__mux4_1 _27292_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03634_));
 sky130_fd_sc_hd__mux4_1 _27293_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03635_));
 sky130_fd_sc_hd__mux4_1 _27294_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03636_));
 sky130_fd_sc_hd__mux4_2 _27295_ (.A0(_03633_),
    .A1(_03634_),
    .A2(_03635_),
    .A3(_03636_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03637_));
 sky130_fd_sc_hd__mux4_1 _27296_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03638_));
 sky130_fd_sc_hd__mux4_1 _27297_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(\count15_2[2] ),
    .S1(net678),
    .X(_03639_));
 sky130_fd_sc_hd__mux4_1 _27298_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03640_));
 sky130_fd_sc_hd__mux4_1 _27299_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_03641_));
 sky130_fd_sc_hd__mux4_1 _27300_ (.A0(_03638_),
    .A1(_03639_),
    .A2(_03640_),
    .A3(_03641_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03642_));
 sky130_fd_sc_hd__mux2i_4 _27301_ (.A0(_03637_),
    .A1(_03642_),
    .S(\count15_2[5] ),
    .Y(_03643_));
 sky130_fd_sc_hd__xnor2_1 _27302_ (.A(_03632_),
    .B(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__xnor2_2 _27303_ (.A(_03377_),
    .B(_03644_),
    .Y(_12055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__mux4_1 _27305_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net565),
    .S1(net570),
    .X(_03646_));
 sky130_fd_sc_hd__mux4_1 _27306_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net565),
    .S1(net570),
    .X(_03647_));
 sky130_fd_sc_hd__mux4_1 _27307_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net565),
    .S1(net570),
    .X(_03648_));
 sky130_fd_sc_hd__mux4_1 _27308_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net565),
    .S1(net570),
    .X(_03649_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__mux4_2 _27310_ (.A0(_03646_),
    .A1(_03647_),
    .A2(_03648_),
    .A3(_03649_),
    .S0(net557),
    .S1(net555),
    .X(_03651_));
 sky130_fd_sc_hd__mux4_1 _27311_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net565),
    .S1(net569),
    .X(_03652_));
 sky130_fd_sc_hd__mux4_1 _27312_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net563),
    .S1(net569),
    .X(_03653_));
 sky130_fd_sc_hd__mux4_1 _27313_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net565),
    .S1(net569),
    .X(_03654_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__mux4_1 _27315_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net563),
    .S1(net569),
    .X(_03656_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__mux4_1 _27317_ (.A0(_03652_),
    .A1(_03653_),
    .A2(_03654_),
    .A3(_03656_),
    .S0(net558),
    .S1(net556),
    .X(_03658_));
 sky130_fd_sc_hd__mux2i_4 _27318_ (.A0(_03651_),
    .A1(_03658_),
    .S(net554),
    .Y(_12054_));
 sky130_fd_sc_hd__mux4_1 _27319_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net636),
    .S1(net646),
    .X(_03659_));
 sky130_fd_sc_hd__mux4_1 _27320_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net636),
    .S1(net647),
    .X(_03660_));
 sky130_fd_sc_hd__mux4_1 _27321_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net636),
    .S1(net646),
    .X(_03661_));
 sky130_fd_sc_hd__mux4_1 _27322_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net636),
    .S1(net646),
    .X(_03662_));
 sky130_fd_sc_hd__mux4_4 _27323_ (.A0(_03659_),
    .A1(_03660_),
    .A2(_03661_),
    .A3(_03662_),
    .S0(\count16_2[3] ),
    .S1(net631),
    .X(_03663_));
 sky130_fd_sc_hd__mux4_1 _27324_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net637),
    .S1(net643),
    .X(_03664_));
 sky130_fd_sc_hd__mux4_1 _27325_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net637),
    .S1(net643),
    .X(_03665_));
 sky130_fd_sc_hd__mux4_1 _27326_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net637),
    .S1(net643),
    .X(_03666_));
 sky130_fd_sc_hd__mux4_1 _27327_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net637),
    .S1(net643),
    .X(_03667_));
 sky130_fd_sc_hd__mux4_1 _27328_ (.A0(_03664_),
    .A1(_03665_),
    .A2(_03666_),
    .A3(_03667_),
    .S0(net633),
    .S1(net631),
    .X(_03668_));
 sky130_fd_sc_hd__mux2i_4 _27329_ (.A0(_03663_),
    .A1(_03668_),
    .S(net629),
    .Y(_12059_));
 sky130_fd_sc_hd__mux4_1 _27330_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net599),
    .S1(net606),
    .X(_03669_));
 sky130_fd_sc_hd__mux4_1 _27331_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net599),
    .S1(net606),
    .X(_03670_));
 sky130_fd_sc_hd__mux4_1 _27332_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net599),
    .S1(net606),
    .X(_03671_));
 sky130_fd_sc_hd__mux4_1 _27333_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net599),
    .S1(net606),
    .X(_03672_));
 sky130_fd_sc_hd__mux4_4 _27334_ (.A0(_03669_),
    .A1(_03670_),
    .A2(_03671_),
    .A3(_03672_),
    .S0(net598),
    .S1(net595),
    .X(_03673_));
 sky130_fd_sc_hd__mux4_1 _27335_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net600),
    .S1(net607),
    .X(_03674_));
 sky130_fd_sc_hd__mux4_1 _27336_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net600),
    .S1(net607),
    .X(_03675_));
 sky130_fd_sc_hd__mux4_1 _27337_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net600),
    .S1(net607),
    .X(_03676_));
 sky130_fd_sc_hd__mux4_1 _27338_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net600),
    .S1(net607),
    .X(_03677_));
 sky130_fd_sc_hd__mux4_1 _27339_ (.A0(_03674_),
    .A1(_03675_),
    .A2(_03676_),
    .A3(_03677_),
    .S0(net598),
    .S1(net594),
    .X(_03678_));
 sky130_fd_sc_hd__mux2i_4 _27340_ (.A0(_03673_),
    .A1(_03678_),
    .S(net592),
    .Y(_03679_));
 sky130_fd_sc_hd__xnor2_1 _27341_ (.A(_03562_),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__xnor2_1 _27342_ (.A(_03135_),
    .B(_03680_),
    .Y(_12064_));
 sky130_fd_sc_hd__mux4_1 _27343_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03681_));
 sky130_fd_sc_hd__mux4_1 _27344_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03682_));
 sky130_fd_sc_hd__mux4_1 _27345_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03683_));
 sky130_fd_sc_hd__mux4_1 _27346_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03684_));
 sky130_fd_sc_hd__mux4_2 _27347_ (.A0(_03681_),
    .A1(_03682_),
    .A2(_03683_),
    .A3(_03684_),
    .S0(net669),
    .S1(net667),
    .X(_03685_));
 sky130_fd_sc_hd__mux4_1 _27348_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03686_));
 sky130_fd_sc_hd__mux4_1 _27349_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03687_));
 sky130_fd_sc_hd__mux4_1 _27350_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03688_));
 sky130_fd_sc_hd__mux4_1 _27351_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net674),
    .S1(net678),
    .X(_03689_));
 sky130_fd_sc_hd__mux4_1 _27352_ (.A0(_03686_),
    .A1(_03687_),
    .A2(_03688_),
    .A3(_03689_),
    .S0(net669),
    .S1(net667),
    .X(_03690_));
 sky130_fd_sc_hd__mux2i_4 _27353_ (.A0(_03685_),
    .A1(_03690_),
    .S(net666),
    .Y(_03691_));
 sky130_fd_sc_hd__mux4_1 _27354_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net672),
    .S1(net679),
    .X(_03692_));
 sky130_fd_sc_hd__mux4_1 _27355_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net672),
    .S1(net679),
    .X(_03693_));
 sky130_fd_sc_hd__mux4_1 _27356_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net672),
    .S1(net679),
    .X(_03694_));
 sky130_fd_sc_hd__mux4_1 _27357_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net672),
    .S1(net679),
    .X(_03695_));
 sky130_fd_sc_hd__mux4_4 _27358_ (.A0(_03692_),
    .A1(_03693_),
    .A2(_03694_),
    .A3(_03695_),
    .S0(net671),
    .S1(net667),
    .X(_03696_));
 sky130_fd_sc_hd__mux4_1 _27359_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net677),
    .S1(net682),
    .X(_03697_));
 sky130_fd_sc_hd__mux4_1 _27360_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net677),
    .S1(net682),
    .X(_03698_));
 sky130_fd_sc_hd__mux4_1 _27361_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net677),
    .S1(net682),
    .X(_03699_));
 sky130_fd_sc_hd__mux4_1 _27362_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net677),
    .S1(net682),
    .X(_03700_));
 sky130_fd_sc_hd__mux4_1 _27363_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03699_),
    .A3(_03700_),
    .S0(net671),
    .S1(net668),
    .X(_03701_));
 sky130_fd_sc_hd__mux2i_4 _27364_ (.A0(_03696_),
    .A1(_03701_),
    .S(\count15_2[5] ),
    .Y(_03702_));
 sky130_fd_sc_hd__xnor2_1 _27365_ (.A(_03691_),
    .B(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__xnor2_2 _27366_ (.A(_03447_),
    .B(_03703_),
    .Y(_12063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__mux4_1 _27368_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03705_));
 sky130_fd_sc_hd__mux4_1 _27369_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03706_));
 sky130_fd_sc_hd__mux4_1 _27370_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__mux4_1 _27372_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__mux4_4 _27374_ (.A0(_03705_),
    .A1(_03706_),
    .A2(_03707_),
    .A3(_03709_),
    .S0(net558),
    .S1(net556),
    .X(_03711_));
 sky130_fd_sc_hd__mux4_1 _27375_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03712_));
 sky130_fd_sc_hd__mux4_1 _27376_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03713_));
 sky130_fd_sc_hd__mux4_1 _27377_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03714_));
 sky130_fd_sc_hd__mux4_1 _27378_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net563),
    .S1(net568),
    .X(_03715_));
 sky130_fd_sc_hd__mux4_1 _27379_ (.A0(_03712_),
    .A1(_03713_),
    .A2(_03714_),
    .A3(_03715_),
    .S0(net558),
    .S1(net556),
    .X(_03716_));
 sky130_fd_sc_hd__mux2i_4 _27380_ (.A0(_03711_),
    .A1(_03716_),
    .S(net554),
    .Y(_12062_));
 sky130_fd_sc_hd__mux4_1 _27381_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net637),
    .S1(net643),
    .X(_03717_));
 sky130_fd_sc_hd__mux4_1 _27382_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net637),
    .S1(net643),
    .X(_03718_));
 sky130_fd_sc_hd__mux4_1 _27383_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net637),
    .S1(net643),
    .X(_03719_));
 sky130_fd_sc_hd__mux4_1 _27384_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net637),
    .S1(net643),
    .X(_03720_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__mux4_4 _27386_ (.A0(_03717_),
    .A1(_03718_),
    .A2(_03719_),
    .A3(_03720_),
    .S0(net633),
    .S1(net632),
    .X(_03722_));
 sky130_fd_sc_hd__mux4_1 _27387_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net638),
    .S1(net645),
    .X(_03723_));
 sky130_fd_sc_hd__mux4_1 _27388_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net638),
    .S1(net645),
    .X(_03724_));
 sky130_fd_sc_hd__mux4_1 _27389_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net638),
    .S1(net645),
    .X(_03725_));
 sky130_fd_sc_hd__mux4_1 _27390_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net638),
    .S1(net645),
    .X(_03726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__mux4_1 _27392_ (.A0(_03723_),
    .A1(_03724_),
    .A2(_03725_),
    .A3(_03726_),
    .S0(net633),
    .S1(net631),
    .X(_03728_));
 sky130_fd_sc_hd__mux2i_4 _27393_ (.A0(_03722_),
    .A1(_03728_),
    .S(net629),
    .Y(_12067_));
 sky130_fd_sc_hd__mux4_1 _27394_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net603),
    .S1(net607),
    .X(_03729_));
 sky130_fd_sc_hd__mux4_1 _27395_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net603),
    .S1(net607),
    .X(_03730_));
 sky130_fd_sc_hd__mux4_1 _27396_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net603),
    .S1(net607),
    .X(_03731_));
 sky130_fd_sc_hd__mux4_1 _27397_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net603),
    .S1(net607),
    .X(_03732_));
 sky130_fd_sc_hd__mux4_4 _27398_ (.A0(_03729_),
    .A1(_03730_),
    .A2(_03731_),
    .A3(_03732_),
    .S0(net596),
    .S1(net595),
    .X(_03733_));
 sky130_fd_sc_hd__mux4_1 _27399_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net603),
    .S1(net605),
    .X(_03734_));
 sky130_fd_sc_hd__mux4_1 _27400_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net603),
    .S1(net605),
    .X(_03735_));
 sky130_fd_sc_hd__mux4_1 _27401_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net603),
    .S1(net605),
    .X(_03736_));
 sky130_fd_sc_hd__mux4_1 _27402_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net603),
    .S1(net605),
    .X(_03737_));
 sky130_fd_sc_hd__mux4_1 _27403_ (.A0(_03734_),
    .A1(_03735_),
    .A2(_03736_),
    .A3(_03737_),
    .S0(net596),
    .S1(net595),
    .X(_03738_));
 sky130_fd_sc_hd__mux2i_4 _27404_ (.A0(_03733_),
    .A1(_03738_),
    .S(net593),
    .Y(_03739_));
 sky130_fd_sc_hd__xnor2_1 _27405_ (.A(_03620_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__xnor2_1 _27406_ (.A(_02910_),
    .B(_03740_),
    .Y(_12072_));
 sky130_fd_sc_hd__mux4_1 _27407_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03741_));
 sky130_fd_sc_hd__mux4_1 _27408_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03742_));
 sky130_fd_sc_hd__mux4_1 _27409_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03743_));
 sky130_fd_sc_hd__mux4_1 _27410_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03744_));
 sky130_fd_sc_hd__mux4_4 _27411_ (.A0(_03741_),
    .A1(_03742_),
    .A2(_03743_),
    .A3(_03744_),
    .S0(net670),
    .S1(net668),
    .X(_03745_));
 sky130_fd_sc_hd__mux4_1 _27412_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03746_));
 sky130_fd_sc_hd__mux4_1 _27413_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03747_));
 sky130_fd_sc_hd__mux4_1 _27414_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03748_));
 sky130_fd_sc_hd__mux4_1 _27415_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net676),
    .S1(net682),
    .X(_03749_));
 sky130_fd_sc_hd__mux4_1 _27416_ (.A0(_03746_),
    .A1(_03747_),
    .A2(_03748_),
    .A3(_03749_),
    .S0(net670),
    .S1(net668),
    .X(_03750_));
 sky130_fd_sc_hd__mux2i_4 _27417_ (.A0(_03745_),
    .A1(_03750_),
    .S(\count15_2[5] ),
    .Y(_03751_));
 sky130_fd_sc_hd__mux4_1 _27418_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03752_));
 sky130_fd_sc_hd__mux4_1 _27419_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03753_));
 sky130_fd_sc_hd__mux4_1 _27420_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03754_));
 sky130_fd_sc_hd__mux4_1 _27421_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03755_));
 sky130_fd_sc_hd__mux4_2 _27422_ (.A0(_03752_),
    .A1(_03753_),
    .A2(_03754_),
    .A3(_03755_),
    .S0(net671),
    .S1(net668),
    .X(_03756_));
 sky130_fd_sc_hd__mux4_1 _27423_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03757_));
 sky130_fd_sc_hd__mux4_1 _27424_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03758_));
 sky130_fd_sc_hd__mux4_1 _27425_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03759_));
 sky130_fd_sc_hd__mux4_1 _27426_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net672),
    .S1(net679),
    .X(_03760_));
 sky130_fd_sc_hd__mux4_1 _27427_ (.A0(_03757_),
    .A1(_03758_),
    .A2(_03759_),
    .A3(_03760_),
    .S0(net671),
    .S1(net668),
    .X(_03761_));
 sky130_fd_sc_hd__mux2i_4 _27428_ (.A0(_03756_),
    .A1(_03761_),
    .S(net665),
    .Y(_03762_));
 sky130_fd_sc_hd__xnor2_1 _27429_ (.A(_03751_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__xnor2_2 _27430_ (.A(_03505_),
    .B(_03763_),
    .Y(_12071_));
 sky130_fd_sc_hd__mux4_1 _27431_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_03764_));
 sky130_fd_sc_hd__mux4_1 _27432_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_03765_));
 sky130_fd_sc_hd__mux4_1 _27433_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_03766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__mux4_1 _27435_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(\count7_2[2] ),
    .S1(net567),
    .X(_03768_));
 sky130_fd_sc_hd__mux4_4 _27436_ (.A0(_03764_),
    .A1(_03765_),
    .A2(_03766_),
    .A3(_03768_),
    .S0(\count7_2[3] ),
    .S1(\count7_2[4] ),
    .X(_03769_));
 sky130_fd_sc_hd__mux4_1 _27437_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net566),
    .S1(net572),
    .X(_03770_));
 sky130_fd_sc_hd__mux4_1 _27438_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net566),
    .S1(net572),
    .X(_03771_));
 sky130_fd_sc_hd__mux4_1 _27439_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net562),
    .S1(net572),
    .X(_03772_));
 sky130_fd_sc_hd__mux4_1 _27440_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net566),
    .S1(net572),
    .X(_03773_));
 sky130_fd_sc_hd__mux4_1 _27441_ (.A0(_03770_),
    .A1(_03771_),
    .A2(_03772_),
    .A3(_03773_),
    .S0(net559),
    .S1(net555),
    .X(_03774_));
 sky130_fd_sc_hd__mux2i_4 _27442_ (.A0(_03769_),
    .A1(_03774_),
    .S(net553),
    .Y(_12070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__mux4_1 _27444_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net640),
    .S1(net645),
    .X(_03776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__mux4_1 _27446_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net640),
    .S1(net645),
    .X(_03778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__mux4_1 _27448_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net640),
    .S1(net645),
    .X(_03780_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__mux4_1 _27450_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net640),
    .S1(net645),
    .X(_03782_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__mux4_4 _27452_ (.A0(_03776_),
    .A1(_03778_),
    .A2(_03780_),
    .A3(_03782_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_03784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__mux4_1 _27454_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net640),
    .S1(net642),
    .X(_03786_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__mux4_1 _27456_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net640),
    .S1(net642),
    .X(_03788_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__mux4_1 _27458_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net640),
    .S1(net642),
    .X(_03790_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__mux4_1 _27460_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net640),
    .S1(net642),
    .X(_03792_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__mux4_1 _27462_ (.A0(_03786_),
    .A1(_03788_),
    .A2(_03790_),
    .A3(_03792_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_03794_));
 sky130_fd_sc_hd__mux2i_4 _27463_ (.A0(_03784_),
    .A1(_03794_),
    .S(net630),
    .Y(_12075_));
 sky130_fd_sc_hd__mux4_1 _27464_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net604),
    .S1(net609),
    .X(_03795_));
 sky130_fd_sc_hd__mux4_1 _27465_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net604),
    .S1(net609),
    .X(_03796_));
 sky130_fd_sc_hd__mux4_1 _27466_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net604),
    .S1(net609),
    .X(_03797_));
 sky130_fd_sc_hd__mux4_1 _27467_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net604),
    .S1(net609),
    .X(_03798_));
 sky130_fd_sc_hd__mux4_4 _27468_ (.A0(_03795_),
    .A1(_03796_),
    .A2(_03797_),
    .A3(_03798_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03799_));
 sky130_fd_sc_hd__mux4_1 _27469_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net602),
    .S1(net609),
    .X(_03800_));
 sky130_fd_sc_hd__mux4_1 _27470_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net602),
    .S1(net605),
    .X(_03801_));
 sky130_fd_sc_hd__mux4_1 _27471_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net602),
    .S1(net605),
    .X(_03802_));
 sky130_fd_sc_hd__mux4_1 _27472_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net602),
    .S1(net605),
    .X(_03803_));
 sky130_fd_sc_hd__mux4_1 _27473_ (.A0(_03800_),
    .A1(_03801_),
    .A2(_03802_),
    .A3(_03803_),
    .S0(net596),
    .S1(\count2_2[4] ),
    .X(_03804_));
 sky130_fd_sc_hd__mux2i_4 _27474_ (.A0(_03799_),
    .A1(_03804_),
    .S(net593),
    .Y(_03805_));
 sky130_fd_sc_hd__xnor2_1 _27475_ (.A(_03679_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__xnor2_1 _27476_ (.A(_03124_),
    .B(_03806_),
    .Y(_12080_));
 sky130_fd_sc_hd__mux4_1 _27477_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net675),
    .S1(net681),
    .X(_03807_));
 sky130_fd_sc_hd__mux4_1 _27478_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net675),
    .S1(net681),
    .X(_03808_));
 sky130_fd_sc_hd__mux4_1 _27479_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net675),
    .S1(net681),
    .X(_03809_));
 sky130_fd_sc_hd__mux4_1 _27480_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net675),
    .S1(net681),
    .X(_03810_));
 sky130_fd_sc_hd__mux4_4 _27481_ (.A0(_03807_),
    .A1(_03808_),
    .A2(_03809_),
    .A3(_03810_),
    .S0(net670),
    .S1(net668),
    .X(_03811_));
 sky130_fd_sc_hd__mux4_1 _27482_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net677),
    .S1(net681),
    .X(_03812_));
 sky130_fd_sc_hd__mux4_1 _27483_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net677),
    .S1(net681),
    .X(_03813_));
 sky130_fd_sc_hd__mux4_1 _27484_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net677),
    .S1(net681),
    .X(_03814_));
 sky130_fd_sc_hd__mux4_1 _27485_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net677),
    .S1(net681),
    .X(_03815_));
 sky130_fd_sc_hd__mux4_1 _27486_ (.A0(_03812_),
    .A1(_03813_),
    .A2(_03814_),
    .A3(_03815_),
    .S0(net671),
    .S1(net668),
    .X(_03816_));
 sky130_fd_sc_hd__mux2i_4 _27487_ (.A0(_03811_),
    .A1(_03816_),
    .S(net665),
    .Y(_03817_));
 sky130_fd_sc_hd__mux4_1 _27488_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03818_));
 sky130_fd_sc_hd__mux4_1 _27489_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03819_));
 sky130_fd_sc_hd__mux4_1 _27490_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03820_));
 sky130_fd_sc_hd__mux4_1 _27491_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03821_));
 sky130_fd_sc_hd__mux4_4 _27492_ (.A0(_03818_),
    .A1(_03819_),
    .A2(_03820_),
    .A3(_03821_),
    .S0(net670),
    .S1(net668),
    .X(_03822_));
 sky130_fd_sc_hd__mux4_1 _27493_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03823_));
 sky130_fd_sc_hd__mux4_1 _27494_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03824_));
 sky130_fd_sc_hd__mux4_1 _27495_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03825_));
 sky130_fd_sc_hd__mux4_1 _27496_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net676),
    .S1(net682),
    .X(_03826_));
 sky130_fd_sc_hd__mux4_1 _27497_ (.A0(_03823_),
    .A1(_03824_),
    .A2(_03825_),
    .A3(_03826_),
    .S0(net670),
    .S1(net668),
    .X(_03827_));
 sky130_fd_sc_hd__mux2i_4 _27498_ (.A0(_03822_),
    .A1(_03827_),
    .S(\count15_2[5] ),
    .Y(_03828_));
 sky130_fd_sc_hd__xnor2_1 _27499_ (.A(_03817_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__xnor2_2 _27500_ (.A(_03585_),
    .B(_03829_),
    .Y(_12079_));
 sky130_fd_sc_hd__mux4_1 _27501_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net564),
    .S1(net568),
    .X(_03830_));
 sky130_fd_sc_hd__mux4_1 _27502_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net564),
    .S1(net568),
    .X(_03831_));
 sky130_fd_sc_hd__mux4_1 _27503_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net564),
    .S1(net568),
    .X(_03832_));
 sky130_fd_sc_hd__mux4_1 _27504_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net564),
    .S1(net568),
    .X(_03833_));
 sky130_fd_sc_hd__mux4_4 _27505_ (.A0(_03830_),
    .A1(_03831_),
    .A2(_03832_),
    .A3(_03833_),
    .S0(net558),
    .S1(net556),
    .X(_03834_));
 sky130_fd_sc_hd__mux4_1 _27506_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net565),
    .S1(net571),
    .X(_03835_));
 sky130_fd_sc_hd__mux4_1 _27507_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net565),
    .S1(net571),
    .X(_03836_));
 sky130_fd_sc_hd__mux4_1 _27508_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net565),
    .S1(net571),
    .X(_03837_));
 sky130_fd_sc_hd__mux4_1 _27509_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net565),
    .S1(net571),
    .X(_03838_));
 sky130_fd_sc_hd__mux4_1 _27510_ (.A0(_03835_),
    .A1(_03836_),
    .A2(_03837_),
    .A3(_03838_),
    .S0(net558),
    .S1(net556),
    .X(_03839_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__mux2i_4 _27512_ (.A0(_03834_),
    .A1(_03839_),
    .S(net554),
    .Y(_12078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__mux4_1 _27514_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03842_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__mux4_1 _27516_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03844_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__mux4_1 _27518_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03846_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__mux4_1 _27520_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03848_));
 sky130_fd_sc_hd__mux4_4 _27521_ (.A0(_03842_),
    .A1(_03844_),
    .A2(_03846_),
    .A3(_03848_),
    .S0(net634),
    .S1(\count16_2[4] ),
    .X(_03849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__mux4_1 _27523_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__mux4_1 _27525_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net640),
    .S1(net645),
    .X(_03853_));
 sky130_fd_sc_hd__fa_1 _27526_ (.A(_11750_),
    .B(_11751_),
    .CIN(_11752_),
    .COUT(_11753_),
    .SUM(_11754_));
 sky130_fd_sc_hd__fa_1 _27527_ (.A(_11755_),
    .B(_11756_),
    .CIN(_11757_),
    .COUT(_11758_),
    .SUM(_11759_));
 sky130_fd_sc_hd__fa_1 _27528_ (.A(_11760_),
    .B(_11753_),
    .CIN(_11759_),
    .COUT(_11761_),
    .SUM(_11762_));
 sky130_fd_sc_hd__fa_1 _27529_ (.A(_11763_),
    .B(_11764_),
    .CIN(_11765_),
    .COUT(_11766_),
    .SUM(_11767_));
 sky130_fd_sc_hd__fa_1 _27530_ (.A(_11768_),
    .B(_11758_),
    .CIN(_11767_),
    .COUT(_11769_),
    .SUM(_11770_));
 sky130_fd_sc_hd__fa_4 _27531_ (.A(_11771_),
    .B(_11761_),
    .CIN(_11770_),
    .COUT(_11772_),
    .SUM(_11773_));
 sky130_fd_sc_hd__fa_1 _27532_ (.A(_11774_),
    .B(_11775_),
    .CIN(_11776_),
    .COUT(_11777_),
    .SUM(_11778_));
 sky130_fd_sc_hd__fa_1 _27533_ (.A(_11779_),
    .B(_11766_),
    .CIN(_11778_),
    .COUT(_11780_),
    .SUM(_11781_));
 sky130_fd_sc_hd__fa_1 _27534_ (.A(_11782_),
    .B(_11783_),
    .CIN(_11784_),
    .COUT(_11785_),
    .SUM(_11786_));
 sky130_fd_sc_hd__fa_1 _27535_ (.A(_11787_),
    .B(_11777_),
    .CIN(_11786_),
    .COUT(_11788_),
    .SUM(_11789_));
 sky130_fd_sc_hd__fa_1 _27536_ (.A(_11790_),
    .B(_11791_),
    .CIN(_11792_),
    .COUT(_11793_),
    .SUM(_11794_));
 sky130_fd_sc_hd__fa_1 _27537_ (.A(_11795_),
    .B(_11785_),
    .CIN(_11794_),
    .COUT(_11796_),
    .SUM(_11797_));
 sky130_fd_sc_hd__fa_2 _27538_ (.A(_11798_),
    .B(_11799_),
    .CIN(_11800_),
    .COUT(_11801_),
    .SUM(_11802_));
 sky130_fd_sc_hd__fa_1 _27539_ (.A(_11803_),
    .B(_11793_),
    .CIN(_11802_),
    .COUT(_11804_),
    .SUM(_11805_));
 sky130_fd_sc_hd__fa_1 _27540_ (.A(_11806_),
    .B(_11807_),
    .CIN(_11808_),
    .COUT(_11809_),
    .SUM(_11810_));
 sky130_fd_sc_hd__fa_1 _27541_ (.A(_11811_),
    .B(_11801_),
    .CIN(_11810_),
    .COUT(_11812_),
    .SUM(_11813_));
 sky130_fd_sc_hd__fa_1 _27542_ (.A(_11814_),
    .B(_11815_),
    .CIN(_11816_),
    .COUT(_11817_),
    .SUM(_11818_));
 sky130_fd_sc_hd__fa_1 _27543_ (.A(_11819_),
    .B(_11809_),
    .CIN(_11818_),
    .COUT(_11820_),
    .SUM(_11821_));
 sky130_fd_sc_hd__fa_1 _27544_ (.A(_11822_),
    .B(_11823_),
    .CIN(_11824_),
    .COUT(_11825_),
    .SUM(_11826_));
 sky130_fd_sc_hd__fa_1 _27545_ (.A(_11827_),
    .B(_11817_),
    .CIN(_11826_),
    .COUT(_11828_),
    .SUM(_11829_));
 sky130_fd_sc_hd__fa_1 _27546_ (.A(_11830_),
    .B(_11831_),
    .CIN(_11832_),
    .COUT(_11833_),
    .SUM(_11834_));
 sky130_fd_sc_hd__fa_1 _27547_ (.A(_11835_),
    .B(_11825_),
    .CIN(_11834_),
    .COUT(_11836_),
    .SUM(_11837_));
 sky130_fd_sc_hd__fa_1 _27548_ (.A(_11838_),
    .B(_11839_),
    .CIN(_11840_),
    .COUT(_11841_),
    .SUM(_11842_));
 sky130_fd_sc_hd__fa_1 _27549_ (.A(_11843_),
    .B(_11833_),
    .CIN(_11842_),
    .COUT(_11844_),
    .SUM(_11845_));
 sky130_fd_sc_hd__fa_1 _27550_ (.A(_11846_),
    .B(_11847_),
    .CIN(_11848_),
    .COUT(_11849_),
    .SUM(_11850_));
 sky130_fd_sc_hd__fa_1 _27551_ (.A(_11851_),
    .B(_11841_),
    .CIN(_11850_),
    .COUT(_11852_),
    .SUM(_11853_));
 sky130_fd_sc_hd__fa_1 _27552_ (.A(_11854_),
    .B(_11855_),
    .CIN(_11856_),
    .COUT(_11857_),
    .SUM(_11858_));
 sky130_fd_sc_hd__fa_1 _27553_ (.A(_11859_),
    .B(_11849_),
    .CIN(_11858_),
    .COUT(_11860_),
    .SUM(_11861_));
 sky130_fd_sc_hd__fa_1 _27554_ (.A(_11862_),
    .B(_11863_),
    .CIN(_11864_),
    .COUT(_11865_),
    .SUM(_11866_));
 sky130_fd_sc_hd__fa_1 _27555_ (.A(_11867_),
    .B(_11857_),
    .CIN(_11866_),
    .COUT(_11868_),
    .SUM(_11869_));
 sky130_fd_sc_hd__fa_1 _27556_ (.A(_11870_),
    .B(_11871_),
    .CIN(_11872_),
    .COUT(_11873_),
    .SUM(_11874_));
 sky130_fd_sc_hd__fa_1 _27557_ (.A(_11875_),
    .B(_11865_),
    .CIN(_11874_),
    .COUT(_11876_),
    .SUM(_11877_));
 sky130_fd_sc_hd__fa_1 _27558_ (.A(_11878_),
    .B(_11879_),
    .CIN(_11880_),
    .COUT(_11881_),
    .SUM(_11882_));
 sky130_fd_sc_hd__fa_1 _27559_ (.A(_11883_),
    .B(_11873_),
    .CIN(_11882_),
    .COUT(_11884_),
    .SUM(_11885_));
 sky130_fd_sc_hd__fa_1 _27560_ (.A(_11886_),
    .B(_11887_),
    .CIN(_11888_),
    .COUT(_11889_),
    .SUM(_11890_));
 sky130_fd_sc_hd__fa_1 _27561_ (.A(_11891_),
    .B(_11881_),
    .CIN(_11890_),
    .COUT(_11892_),
    .SUM(_11893_));
 sky130_fd_sc_hd__fa_1 _27562_ (.A(_11894_),
    .B(_11895_),
    .CIN(_11896_),
    .COUT(_11897_),
    .SUM(_11898_));
 sky130_fd_sc_hd__fa_1 _27563_ (.A(_11899_),
    .B(_11889_),
    .CIN(_11898_),
    .COUT(_11900_),
    .SUM(_11901_));
 sky130_fd_sc_hd__fa_1 _27564_ (.A(_11902_),
    .B(_11903_),
    .CIN(_11904_),
    .COUT(_11905_),
    .SUM(_11906_));
 sky130_fd_sc_hd__fa_1 _27565_ (.A(_11907_),
    .B(_11897_),
    .CIN(_11906_),
    .COUT(_11908_),
    .SUM(_11909_));
 sky130_fd_sc_hd__fa_1 _27566_ (.A(_11910_),
    .B(_11911_),
    .CIN(_11912_),
    .COUT(_11913_),
    .SUM(_11914_));
 sky130_fd_sc_hd__fa_1 _27567_ (.A(_11915_),
    .B(_11905_),
    .CIN(_11914_),
    .COUT(_11916_),
    .SUM(_11917_));
 sky130_fd_sc_hd__fa_1 _27568_ (.A(_11918_),
    .B(_11919_),
    .CIN(_11920_),
    .COUT(_11921_),
    .SUM(_11922_));
 sky130_fd_sc_hd__fa_1 _27569_ (.A(_11923_),
    .B(_11913_),
    .CIN(_11922_),
    .COUT(_11924_),
    .SUM(_11925_));
 sky130_fd_sc_hd__fa_1 _27570_ (.A(_11926_),
    .B(_11927_),
    .CIN(_11928_),
    .COUT(_11929_),
    .SUM(_11930_));
 sky130_fd_sc_hd__fa_1 _27571_ (.A(_11931_),
    .B(_11921_),
    .CIN(_11930_),
    .COUT(_11932_),
    .SUM(_11933_));
 sky130_fd_sc_hd__fa_1 _27572_ (.A(_11934_),
    .B(_11935_),
    .CIN(_11936_),
    .COUT(_11937_),
    .SUM(_11938_));
 sky130_fd_sc_hd__fa_1 _27573_ (.A(_11939_),
    .B(_11929_),
    .CIN(_11938_),
    .COUT(_11940_),
    .SUM(_11941_));
 sky130_fd_sc_hd__fa_1 _27574_ (.A(_11942_),
    .B(_11943_),
    .CIN(_11944_),
    .COUT(_11945_),
    .SUM(_11946_));
 sky130_fd_sc_hd__fa_1 _27575_ (.A(_11947_),
    .B(_11937_),
    .CIN(_11946_),
    .COUT(_11948_),
    .SUM(_11949_));
 sky130_fd_sc_hd__fa_1 _27576_ (.A(_11950_),
    .B(_11951_),
    .CIN(_11952_),
    .COUT(_11953_),
    .SUM(_11954_));
 sky130_fd_sc_hd__fa_1 _27577_ (.A(_11955_),
    .B(_11945_),
    .CIN(_11954_),
    .COUT(_11956_),
    .SUM(_11957_));
 sky130_fd_sc_hd__fa_1 _27578_ (.A(_11958_),
    .B(_11959_),
    .CIN(_11960_),
    .COUT(_11961_),
    .SUM(_11962_));
 sky130_fd_sc_hd__fa_1 _27579_ (.A(_11963_),
    .B(_11953_),
    .CIN(_11962_),
    .COUT(_11964_),
    .SUM(_11965_));
 sky130_fd_sc_hd__fa_1 _27580_ (.A(_11966_),
    .B(_11967_),
    .CIN(_11968_),
    .COUT(_11969_),
    .SUM(_11970_));
 sky130_fd_sc_hd__fa_1 _27581_ (.A(_11971_),
    .B(_11961_),
    .CIN(_11970_),
    .COUT(_11972_),
    .SUM(_11973_));
 sky130_fd_sc_hd__fa_1 _27582_ (.A(_11974_),
    .B(_11975_),
    .CIN(_11976_),
    .COUT(_11977_),
    .SUM(_11978_));
 sky130_fd_sc_hd__fa_1 _27583_ (.A(_11979_),
    .B(_11969_),
    .CIN(_11978_),
    .COUT(_11980_),
    .SUM(_11981_));
 sky130_fd_sc_hd__fa_1 _27584_ (.A(_11982_),
    .B(_11983_),
    .CIN(_11984_),
    .COUT(_11985_),
    .SUM(_11986_));
 sky130_fd_sc_hd__fa_1 _27585_ (.A(_11987_),
    .B(_11977_),
    .CIN(_11986_),
    .COUT(_11988_),
    .SUM(_11989_));
 sky130_fd_sc_hd__fa_1 _27586_ (.A(_11990_),
    .B(_11991_),
    .CIN(_11992_),
    .COUT(_11993_),
    .SUM(_11994_));
 sky130_fd_sc_hd__fa_1 _27587_ (.A(_11995_),
    .B(_11985_),
    .CIN(_11994_),
    .COUT(_11996_),
    .SUM(_11997_));
 sky130_fd_sc_hd__fa_2 _27588_ (.A(_11998_),
    .B(_11999_),
    .CIN(_12000_),
    .COUT(_12001_),
    .SUM(_12002_));
 sky130_fd_sc_hd__fa_1 _27589_ (.A(_12003_),
    .B(_12004_),
    .CIN(_12005_),
    .COUT(_12006_),
    .SUM(_12007_));
 sky130_fd_sc_hd__fa_1 _27590_ (.A(_12008_),
    .B(_12001_),
    .CIN(_12007_),
    .COUT(_12009_),
    .SUM(_12010_));
 sky130_fd_sc_hd__fa_1 _27591_ (.A(_12011_),
    .B(_12012_),
    .CIN(_12013_),
    .COUT(_12014_),
    .SUM(_12015_));
 sky130_fd_sc_hd__fa_1 _27592_ (.A(_12016_),
    .B(_12006_),
    .CIN(_12015_),
    .COUT(_12017_),
    .SUM(_12018_));
 sky130_fd_sc_hd__fa_4 _27593_ (.A(_12019_),
    .B(_12009_),
    .CIN(_12018_),
    .COUT(_12020_),
    .SUM(_12021_));
 sky130_fd_sc_hd__fa_1 _27594_ (.A(_12022_),
    .B(_12023_),
    .CIN(_12024_),
    .COUT(_12025_),
    .SUM(_12026_));
 sky130_fd_sc_hd__fa_1 _27595_ (.A(_12027_),
    .B(_12014_),
    .CIN(_12026_),
    .COUT(_12028_),
    .SUM(_12029_));
 sky130_fd_sc_hd__fa_1 _27596_ (.A(_12030_),
    .B(_12031_),
    .CIN(_12032_),
    .COUT(_12033_),
    .SUM(_12034_));
 sky130_fd_sc_hd__fa_1 _27597_ (.A(_12035_),
    .B(_12025_),
    .CIN(_12034_),
    .COUT(_12036_),
    .SUM(_12037_));
 sky130_fd_sc_hd__fa_1 _27598_ (.A(_12038_),
    .B(_12039_),
    .CIN(_12040_),
    .COUT(_12041_),
    .SUM(_12042_));
 sky130_fd_sc_hd__fa_1 _27599_ (.A(_12043_),
    .B(_12033_),
    .CIN(_12042_),
    .COUT(_12044_),
    .SUM(_12045_));
 sky130_fd_sc_hd__fa_1 _27600_ (.A(_12046_),
    .B(_12047_),
    .CIN(_12048_),
    .COUT(_12049_),
    .SUM(_12050_));
 sky130_fd_sc_hd__fa_1 _27601_ (.A(_12051_),
    .B(_12041_),
    .CIN(_12050_),
    .COUT(_12052_),
    .SUM(_12053_));
 sky130_fd_sc_hd__fa_1 _27602_ (.A(_12054_),
    .B(_12055_),
    .CIN(_12056_),
    .COUT(_12057_),
    .SUM(_12058_));
 sky130_fd_sc_hd__fa_1 _27603_ (.A(_12059_),
    .B(_12049_),
    .CIN(_12058_),
    .COUT(_12060_),
    .SUM(_12061_));
 sky130_fd_sc_hd__fa_1 _27604_ (.A(_12062_),
    .B(_12063_),
    .CIN(_12064_),
    .COUT(_12065_),
    .SUM(_12066_));
 sky130_fd_sc_hd__fa_1 _27605_ (.A(_12067_),
    .B(_12057_),
    .CIN(_12066_),
    .COUT(_12068_),
    .SUM(_12069_));
 sky130_fd_sc_hd__fa_1 _27606_ (.A(_12070_),
    .B(_12071_),
    .CIN(_12072_),
    .COUT(_12073_),
    .SUM(_12074_));
 sky130_fd_sc_hd__fa_1 _27607_ (.A(_12075_),
    .B(_12065_),
    .CIN(_12074_),
    .COUT(_12076_),
    .SUM(_12077_));
 sky130_fd_sc_hd__fa_1 _27608_ (.A(_12078_),
    .B(_12079_),
    .CIN(_12080_),
    .COUT(_12081_),
    .SUM(_12082_));
 sky130_fd_sc_hd__fa_1 _27609_ (.A(_12083_),
    .B(_12073_),
    .CIN(_12082_),
    .COUT(_12084_),
    .SUM(_12085_));
 sky130_fd_sc_hd__fa_2 _27610_ (.A(_12086_),
    .B(_12087_),
    .CIN(_12088_),
    .COUT(_12089_),
    .SUM(_12090_));
 sky130_fd_sc_hd__fa_1 _27611_ (.A(_12091_),
    .B(_12081_),
    .CIN(_12090_),
    .COUT(_12092_),
    .SUM(_12093_));
 sky130_fd_sc_hd__fa_1 _27612_ (.A(_12094_),
    .B(_12095_),
    .CIN(_12096_),
    .COUT(_12097_),
    .SUM(_12098_));
 sky130_fd_sc_hd__fa_1 _27613_ (.A(_12099_),
    .B(_12089_),
    .CIN(_12098_),
    .COUT(_12100_),
    .SUM(_12101_));
 sky130_fd_sc_hd__fa_1 _27614_ (.A(_12102_),
    .B(_12103_),
    .CIN(_12104_),
    .COUT(_12105_),
    .SUM(_12106_));
 sky130_fd_sc_hd__fa_1 _27615_ (.A(_12107_),
    .B(_12097_),
    .CIN(_12106_),
    .COUT(_12108_),
    .SUM(_12109_));
 sky130_fd_sc_hd__fa_1 _27616_ (.A(_12110_),
    .B(_12111_),
    .CIN(_12112_),
    .COUT(_12113_),
    .SUM(_12114_));
 sky130_fd_sc_hd__fa_1 _27617_ (.A(_12115_),
    .B(_12105_),
    .CIN(_12114_),
    .COUT(_12116_),
    .SUM(_12117_));
 sky130_fd_sc_hd__fa_1 _27618_ (.A(_12118_),
    .B(_12119_),
    .CIN(_12120_),
    .COUT(_12121_),
    .SUM(_12122_));
 sky130_fd_sc_hd__fa_1 _27619_ (.A(_12123_),
    .B(_12113_),
    .CIN(_12122_),
    .COUT(_12124_),
    .SUM(_12125_));
 sky130_fd_sc_hd__fa_1 _27620_ (.A(_12126_),
    .B(_12127_),
    .CIN(_12128_),
    .COUT(_12129_),
    .SUM(_12130_));
 sky130_fd_sc_hd__fa_1 _27621_ (.A(_12131_),
    .B(_12121_),
    .CIN(_12130_),
    .COUT(_12132_),
    .SUM(_12133_));
 sky130_fd_sc_hd__fa_1 _27622_ (.A(_12134_),
    .B(_12135_),
    .CIN(_12136_),
    .COUT(_12137_),
    .SUM(_12138_));
 sky130_fd_sc_hd__fa_1 _27623_ (.A(_12139_),
    .B(_12129_),
    .CIN(_12138_),
    .COUT(_12140_),
    .SUM(_12141_));
 sky130_fd_sc_hd__fa_1 _27624_ (.A(_12142_),
    .B(_12143_),
    .CIN(_12144_),
    .COUT(_12145_),
    .SUM(_12146_));
 sky130_fd_sc_hd__fa_1 _27625_ (.A(_12147_),
    .B(_12137_),
    .CIN(_12146_),
    .COUT(_12148_),
    .SUM(_12149_));
 sky130_fd_sc_hd__fa_1 _27626_ (.A(_12150_),
    .B(_12151_),
    .CIN(_12152_),
    .COUT(_12153_),
    .SUM(_12154_));
 sky130_fd_sc_hd__fa_1 _27627_ (.A(_12155_),
    .B(_12145_),
    .CIN(_12154_),
    .COUT(_12156_),
    .SUM(_12157_));
 sky130_fd_sc_hd__fa_1 _27628_ (.A(_12158_),
    .B(_12159_),
    .CIN(_12160_),
    .COUT(_12161_),
    .SUM(_12162_));
 sky130_fd_sc_hd__fa_1 _27629_ (.A(_12163_),
    .B(_12153_),
    .CIN(_12162_),
    .COUT(_12164_),
    .SUM(_12165_));
 sky130_fd_sc_hd__fa_1 _27630_ (.A(_12166_),
    .B(_12167_),
    .CIN(_12168_),
    .COUT(_12169_),
    .SUM(_12170_));
 sky130_fd_sc_hd__fa_1 _27631_ (.A(_12171_),
    .B(_12161_),
    .CIN(_12170_),
    .COUT(_12172_),
    .SUM(_12173_));
 sky130_fd_sc_hd__fa_1 _27632_ (.A(_12174_),
    .B(_12175_),
    .CIN(_12176_),
    .COUT(_12177_),
    .SUM(_12178_));
 sky130_fd_sc_hd__fa_1 _27633_ (.A(_12179_),
    .B(_12169_),
    .CIN(_12178_),
    .COUT(_12180_),
    .SUM(_12181_));
 sky130_fd_sc_hd__fa_1 _27634_ (.A(_12182_),
    .B(_12183_),
    .CIN(_12184_),
    .COUT(_12185_),
    .SUM(_12186_));
 sky130_fd_sc_hd__fa_1 _27635_ (.A(_12187_),
    .B(_12177_),
    .CIN(_12186_),
    .COUT(_12188_),
    .SUM(_12189_));
 sky130_fd_sc_hd__fa_2 _27636_ (.A(_12190_),
    .B(_12191_),
    .CIN(_12192_),
    .COUT(_12193_),
    .SUM(_12194_));
 sky130_fd_sc_hd__fa_1 _27637_ (.A(_12195_),
    .B(_12185_),
    .CIN(_12194_),
    .COUT(_12196_),
    .SUM(_12197_));
 sky130_fd_sc_hd__fa_1 _27638_ (.A(_12198_),
    .B(_12199_),
    .CIN(_12200_),
    .COUT(_12201_),
    .SUM(_12202_));
 sky130_fd_sc_hd__fa_1 _27639_ (.A(_12203_),
    .B(_12193_),
    .CIN(_12202_),
    .COUT(_12204_),
    .SUM(_12205_));
 sky130_fd_sc_hd__fa_1 _27640_ (.A(_12206_),
    .B(_12207_),
    .CIN(_12208_),
    .COUT(_12209_),
    .SUM(_12210_));
 sky130_fd_sc_hd__fa_1 _27641_ (.A(_12211_),
    .B(_12201_),
    .CIN(_12210_),
    .COUT(_12212_),
    .SUM(_12213_));
 sky130_fd_sc_hd__fa_1 _27642_ (.A(_12214_),
    .B(_12215_),
    .CIN(_12216_),
    .COUT(_12217_),
    .SUM(_12218_));
 sky130_fd_sc_hd__fa_1 _27643_ (.A(_12219_),
    .B(_12209_),
    .CIN(_12218_),
    .COUT(_12220_),
    .SUM(_12221_));
 sky130_fd_sc_hd__fa_1 _27644_ (.A(_12222_),
    .B(_12223_),
    .CIN(_12224_),
    .COUT(_12225_),
    .SUM(_12226_));
 sky130_fd_sc_hd__fa_1 _27645_ (.A(_12227_),
    .B(_12217_),
    .CIN(_12226_),
    .COUT(_12228_),
    .SUM(_12229_));
 sky130_fd_sc_hd__fa_1 _27646_ (.A(_12230_),
    .B(_12231_),
    .CIN(_12232_),
    .COUT(_12233_),
    .SUM(_12234_));
 sky130_fd_sc_hd__fa_1 _27647_ (.A(_12235_),
    .B(_12225_),
    .CIN(_12234_),
    .COUT(_12236_),
    .SUM(_12237_));
 sky130_fd_sc_hd__fa_1 _27648_ (.A(_12238_),
    .B(_12239_),
    .CIN(_12240_),
    .COUT(_12241_),
    .SUM(_12242_));
 sky130_fd_sc_hd__fa_1 _27649_ (.A(_12243_),
    .B(_12233_),
    .CIN(_12242_),
    .COUT(_12244_),
    .SUM(_12245_));
 sky130_fd_sc_hd__fa_1 _27650_ (.A(_12246_),
    .B(_12247_),
    .CIN(_12248_),
    .COUT(_12249_),
    .SUM(_12250_));
 sky130_fd_sc_hd__fa_4 _27651_ (.A(\hash.CA2.p1[1] ),
    .B(\hash.CA2.p3[1] ),
    .CIN(_12251_),
    .COUT(_12252_),
    .SUM(_12253_));
 sky130_fd_sc_hd__fa_2 _27652_ (.A(_12256_),
    .B(_12255_),
    .CIN(_12254_),
    .COUT(_12257_),
    .SUM(_12258_));
 sky130_fd_sc_hd__fa_1 _27653_ (.A(_12259_),
    .B(_12260_),
    .CIN(_12261_),
    .COUT(_12262_),
    .SUM(_12263_));
 sky130_fd_sc_hd__fa_1 _27654_ (.A(\hash.CA2.p4[1] ),
    .B(_12264_),
    .CIN(_12265_),
    .COUT(_12266_),
    .SUM(_12267_));
 sky130_fd_sc_hd__fa_1 _27655_ (.A(_12268_),
    .B(_12269_),
    .CIN(_12270_),
    .COUT(_12271_),
    .SUM(_12272_));
 sky130_fd_sc_hd__fa_1 _27656_ (.A(\hash.CA2.p4[2] ),
    .B(_12273_),
    .CIN(_12274_),
    .COUT(_12275_),
    .SUM(_12276_));
 sky130_fd_sc_hd__fa_4 _27657_ (.A(_12277_),
    .B(_12278_),
    .CIN(_12279_),
    .COUT(_12280_),
    .SUM(_12281_));
 sky130_fd_sc_hd__fa_1 _27658_ (.A(_12282_),
    .B(_12283_),
    .CIN(_12284_),
    .COUT(_12285_),
    .SUM(_12286_));
 sky130_fd_sc_hd__fa_1 _27659_ (.A(\hash.CA2.p4[3] ),
    .B(_12287_),
    .CIN(_12288_),
    .COUT(_12289_),
    .SUM(_12290_));
 sky130_fd_sc_hd__fa_1 _27660_ (.A(_12291_),
    .B(_12292_),
    .CIN(_12293_),
    .COUT(_12294_),
    .SUM(_12295_));
 sky130_fd_sc_hd__fa_1 _27661_ (.A(\hash.CA2.p4[4] ),
    .B(_12296_),
    .CIN(_12297_),
    .COUT(_12298_),
    .SUM(_12299_));
 sky130_fd_sc_hd__fa_1 _27662_ (.A(_12300_),
    .B(_12301_),
    .CIN(_12302_),
    .COUT(_12303_),
    .SUM(_12304_));
 sky130_fd_sc_hd__fa_1 _27663_ (.A(\hash.CA2.p4[5] ),
    .B(_12305_),
    .CIN(_12306_),
    .COUT(_12307_),
    .SUM(_12308_));
 sky130_fd_sc_hd__fa_1 _27664_ (.A(_12309_),
    .B(_12310_),
    .CIN(_12311_),
    .COUT(_12312_),
    .SUM(_12313_));
 sky130_fd_sc_hd__fa_1 _27665_ (.A(\hash.CA2.p4[6] ),
    .B(_12314_),
    .CIN(_12315_),
    .COUT(_12316_),
    .SUM(_12317_));
 sky130_fd_sc_hd__fa_1 _27666_ (.A(_12318_),
    .B(_12319_),
    .CIN(_12320_),
    .COUT(_12321_),
    .SUM(_12322_));
 sky130_fd_sc_hd__fa_1 _27667_ (.A(\hash.CA2.p4[7] ),
    .B(_12323_),
    .CIN(_12324_),
    .COUT(_12325_),
    .SUM(_12326_));
 sky130_fd_sc_hd__fa_1 _27668_ (.A(_12327_),
    .B(_12328_),
    .CIN(_12329_),
    .COUT(_12330_),
    .SUM(_12331_));
 sky130_fd_sc_hd__fa_1 _27669_ (.A(\hash.CA2.p4[8] ),
    .B(_12332_),
    .CIN(_12333_),
    .COUT(_12334_),
    .SUM(_12335_));
 sky130_fd_sc_hd__fa_1 _27670_ (.A(_12336_),
    .B(_12337_),
    .CIN(_12338_),
    .COUT(_12339_),
    .SUM(_12340_));
 sky130_fd_sc_hd__fa_1 _27671_ (.A(\hash.CA2.p4[9] ),
    .B(_12341_),
    .CIN(_12342_),
    .COUT(_12343_),
    .SUM(_12344_));
 sky130_fd_sc_hd__fa_1 _27672_ (.A(_12345_),
    .B(_12346_),
    .CIN(_12347_),
    .COUT(_12348_),
    .SUM(_12349_));
 sky130_fd_sc_hd__fa_1 _27673_ (.A(\hash.CA2.p4[10] ),
    .B(_12350_),
    .CIN(_12351_),
    .COUT(_12352_),
    .SUM(_12353_));
 sky130_fd_sc_hd__fa_1 _27674_ (.A(_12354_),
    .B(_12355_),
    .CIN(_12356_),
    .COUT(_12357_),
    .SUM(_12358_));
 sky130_fd_sc_hd__fa_1 _27675_ (.A(\hash.CA2.p4[11] ),
    .B(_12359_),
    .CIN(_12360_),
    .COUT(_12361_),
    .SUM(_12362_));
 sky130_fd_sc_hd__fa_1 _27676_ (.A(_12363_),
    .B(_12364_),
    .CIN(_12365_),
    .COUT(_12366_),
    .SUM(_12367_));
 sky130_fd_sc_hd__fa_1 _27677_ (.A(\hash.CA2.p4[12] ),
    .B(_12368_),
    .CIN(_12369_),
    .COUT(_12370_),
    .SUM(_12371_));
 sky130_fd_sc_hd__fa_1 _27678_ (.A(_12372_),
    .B(_12373_),
    .CIN(_12374_),
    .COUT(_12375_),
    .SUM(_12376_));
 sky130_fd_sc_hd__fa_1 _27679_ (.A(\hash.CA2.p4[13] ),
    .B(_12378_),
    .CIN(_12377_),
    .COUT(_12379_),
    .SUM(_12380_));
 sky130_fd_sc_hd__fa_1 _27680_ (.A(_12381_),
    .B(_12382_),
    .CIN(_12383_),
    .COUT(_12384_),
    .SUM(_12385_));
 sky130_fd_sc_hd__fa_1 _27681_ (.A(\hash.CA2.p4[14] ),
    .B(_12386_),
    .CIN(_12387_),
    .COUT(_12388_),
    .SUM(_12389_));
 sky130_fd_sc_hd__fa_1 _27682_ (.A(_12390_),
    .B(_12391_),
    .CIN(_12392_),
    .COUT(_12393_),
    .SUM(_12394_));
 sky130_fd_sc_hd__fa_1 _27683_ (.A(\hash.CA2.p4[15] ),
    .B(_12395_),
    .CIN(_12396_),
    .COUT(_12397_),
    .SUM(_12398_));
 sky130_fd_sc_hd__fa_1 _27684_ (.A(_12399_),
    .B(_12400_),
    .CIN(_12401_),
    .COUT(_12402_),
    .SUM(_12403_));
 sky130_fd_sc_hd__fa_1 _27685_ (.A(\hash.CA2.p4[16] ),
    .B(_12404_),
    .CIN(_12405_),
    .COUT(_12406_),
    .SUM(_12407_));
 sky130_fd_sc_hd__fa_1 _27686_ (.A(_12408_),
    .B(_12409_),
    .CIN(_12410_),
    .COUT(_12411_),
    .SUM(_12412_));
 sky130_fd_sc_hd__fa_1 _27687_ (.A(\hash.CA2.p4[17] ),
    .B(_12413_),
    .CIN(_12414_),
    .COUT(_12415_),
    .SUM(_12416_));
 sky130_fd_sc_hd__fa_1 _27688_ (.A(_12417_),
    .B(_12418_),
    .CIN(_12419_),
    .COUT(_12420_),
    .SUM(_12421_));
 sky130_fd_sc_hd__fa_1 _27689_ (.A(\hash.CA2.p4[18] ),
    .B(_12422_),
    .CIN(_12423_),
    .COUT(_12424_),
    .SUM(_12425_));
 sky130_fd_sc_hd__fa_1 _27690_ (.A(_12426_),
    .B(_12427_),
    .CIN(_12428_),
    .COUT(_12429_),
    .SUM(_12430_));
 sky130_fd_sc_hd__fa_1 _27691_ (.A(\hash.CA2.p4[19] ),
    .B(_12431_),
    .CIN(_12432_),
    .COUT(_12433_),
    .SUM(_12434_));
 sky130_fd_sc_hd__fa_1 _27692_ (.A(_12435_),
    .B(_12436_),
    .CIN(_12437_),
    .COUT(_12438_),
    .SUM(_12439_));
 sky130_fd_sc_hd__fa_1 _27693_ (.A(\hash.CA2.p4[20] ),
    .B(_12440_),
    .CIN(_12441_),
    .COUT(_12442_),
    .SUM(_12443_));
 sky130_fd_sc_hd__fa_1 _27694_ (.A(_12444_),
    .B(_12445_),
    .CIN(_12446_),
    .COUT(_12447_),
    .SUM(_12448_));
 sky130_fd_sc_hd__fa_1 _27695_ (.A(\hash.CA2.p4[21] ),
    .B(_12449_),
    .CIN(_12450_),
    .COUT(_12451_),
    .SUM(_12452_));
 sky130_fd_sc_hd__fa_1 _27696_ (.A(_12453_),
    .B(_12454_),
    .CIN(_12455_),
    .COUT(_12456_),
    .SUM(_12457_));
 sky130_fd_sc_hd__fa_1 _27697_ (.A(\hash.CA2.p4[22] ),
    .B(_12458_),
    .CIN(_12459_),
    .COUT(_12460_),
    .SUM(_12461_));
 sky130_fd_sc_hd__fa_1 _27698_ (.A(_12462_),
    .B(_12463_),
    .CIN(_12464_),
    .COUT(_12465_),
    .SUM(_12466_));
 sky130_fd_sc_hd__fa_1 _27699_ (.A(\hash.CA2.p4[23] ),
    .B(_12467_),
    .CIN(_12468_),
    .COUT(_12469_),
    .SUM(_12470_));
 sky130_fd_sc_hd__fa_1 _27700_ (.A(_12471_),
    .B(_12472_),
    .CIN(_12473_),
    .COUT(_12474_),
    .SUM(_12475_));
 sky130_fd_sc_hd__fa_1 _27701_ (.A(\hash.CA2.p4[24] ),
    .B(_12476_),
    .CIN(_12477_),
    .COUT(_12478_),
    .SUM(_12479_));
 sky130_fd_sc_hd__fa_1 _27702_ (.A(_12480_),
    .B(_12481_),
    .CIN(_12482_),
    .COUT(_12483_),
    .SUM(_12484_));
 sky130_fd_sc_hd__fa_1 _27703_ (.A(\hash.CA2.p4[25] ),
    .B(_12485_),
    .CIN(_12486_),
    .COUT(_12487_),
    .SUM(_12488_));
 sky130_fd_sc_hd__fa_1 _27704_ (.A(_12489_),
    .B(_12490_),
    .CIN(_12491_),
    .COUT(_12492_),
    .SUM(_12493_));
 sky130_fd_sc_hd__fa_1 _27705_ (.A(\hash.CA2.p4[26] ),
    .B(_12494_),
    .CIN(_12495_),
    .COUT(_12496_),
    .SUM(_12497_));
 sky130_fd_sc_hd__fa_1 _27706_ (.A(_12498_),
    .B(_12499_),
    .CIN(_12500_),
    .COUT(_12501_),
    .SUM(_12502_));
 sky130_fd_sc_hd__fa_1 _27707_ (.A(\hash.CA2.p4[27] ),
    .B(_12503_),
    .CIN(_12504_),
    .COUT(_12505_),
    .SUM(_12506_));
 sky130_fd_sc_hd__fa_1 _27708_ (.A(_12507_),
    .B(_12508_),
    .CIN(_12509_),
    .COUT(_12510_),
    .SUM(_12511_));
 sky130_fd_sc_hd__fa_1 _27709_ (.A(\hash.CA2.p4[28] ),
    .B(_12512_),
    .CIN(_12513_),
    .COUT(_12514_),
    .SUM(_12515_));
 sky130_fd_sc_hd__fa_1 _27710_ (.A(_12516_),
    .B(_12517_),
    .CIN(_12518_),
    .COUT(_12519_),
    .SUM(_12520_));
 sky130_fd_sc_hd__fa_1 _27711_ (.A(\hash.CA2.p4[29] ),
    .B(_12521_),
    .CIN(_12522_),
    .COUT(_12523_),
    .SUM(_12524_));
 sky130_fd_sc_hd__fa_1 _27712_ (.A(_12525_),
    .B(_12526_),
    .CIN(_12527_),
    .COUT(_12528_),
    .SUM(_12529_));
 sky130_fd_sc_hd__fa_1 _27713_ (.A(\hash.CA2.p4[30] ),
    .B(_12530_),
    .CIN(_12531_),
    .COUT(_12532_),
    .SUM(_12533_));
 sky130_fd_sc_hd__fa_4 _27714_ (.A(\hash.CA2.p5[1] ),
    .B(_12534_),
    .CIN(_12258_),
    .COUT(_12535_),
    .SUM(_12536_));
 sky130_fd_sc_hd__fa_1 _27715_ (.A(_12537_),
    .B(_12538_),
    .CIN(_12539_),
    .COUT(_12540_),
    .SUM(_12541_));
 sky130_fd_sc_hd__fa_4 _27716_ (.A(_12542_),
    .B(_12543_),
    .CIN(_00843_),
    .COUT(_12544_),
    .SUM(_12545_));
 sky130_fd_sc_hd__fa_1 _27717_ (.A(\hash.CA1.k_i2[2] ),
    .B(\hash.CA1.w_i2[2] ),
    .CIN(_12546_),
    .COUT(_12547_),
    .SUM(_12548_));
 sky130_fd_sc_hd__fa_4 _27718_ (.A(_12549_),
    .B(_12550_),
    .CIN(_12548_),
    .COUT(_12551_),
    .SUM(\hash.CA1.p4[2] ));
 sky130_fd_sc_hd__fa_1 _27719_ (.A(_12552_),
    .B(_12553_),
    .CIN(_12554_),
    .COUT(_12555_),
    .SUM(_12556_));
 sky130_fd_sc_hd__fa_1 _27720_ (.A(\hash.CA1.k_i2[4] ),
    .B(\hash.CA1.w_i2[4] ),
    .CIN(_12557_),
    .COUT(_12558_),
    .SUM(_12559_));
 sky130_fd_sc_hd__fa_1 _27721_ (.A(_12560_),
    .B(_12561_),
    .CIN(_12562_),
    .COUT(_12563_),
    .SUM(_12564_));
 sky130_fd_sc_hd__fa_1 _27722_ (.A(\hash.CA1.k_i2[6] ),
    .B(\hash.CA1.w_i2[6] ),
    .CIN(_12565_),
    .COUT(_12566_),
    .SUM(_12567_));
 sky130_fd_sc_hd__fa_1 _27723_ (.A(_12568_),
    .B(_12569_),
    .CIN(_12570_),
    .COUT(_12571_),
    .SUM(_12572_));
 sky130_fd_sc_hd__fa_1 _27724_ (.A(_12573_),
    .B(_12574_),
    .CIN(_12575_),
    .COUT(_12576_),
    .SUM(_12577_));
 sky130_fd_sc_hd__fa_1 _27725_ (.A(\hash.CA1.k_i2[9] ),
    .B(\hash.CA1.w_i2[9] ),
    .CIN(_12578_),
    .COUT(_12579_),
    .SUM(_12580_));
 sky130_fd_sc_hd__fa_1 _27726_ (.A(\hash.CA1.k_i2[10] ),
    .B(\hash.CA1.w_i2[10] ),
    .CIN(_12581_),
    .COUT(_12582_),
    .SUM(_12583_));
 sky130_fd_sc_hd__fa_1 _27727_ (.A(_12584_),
    .B(_12585_),
    .CIN(_12586_),
    .COUT(_12587_),
    .SUM(_12588_));
 sky130_fd_sc_hd__fa_1 _27728_ (.A(_12589_),
    .B(_12590_),
    .CIN(_12591_),
    .COUT(_12592_),
    .SUM(_12593_));
 sky130_fd_sc_hd__fa_1 _27729_ (.A(\hash.CA1.k_i2[13] ),
    .B(\hash.CA1.w_i2[13] ),
    .CIN(_12594_),
    .COUT(_12595_),
    .SUM(_12596_));
 sky130_fd_sc_hd__fa_1 _27730_ (.A(_12597_),
    .B(_12598_),
    .CIN(_12599_),
    .COUT(_12600_),
    .SUM(_12601_));
 sky130_fd_sc_hd__fa_1 _27731_ (.A(_12602_),
    .B(_12603_),
    .CIN(_12604_),
    .COUT(_12605_),
    .SUM(_12606_));
 sky130_fd_sc_hd__fa_1 _27732_ (.A(_12607_),
    .B(_12608_),
    .CIN(_12609_),
    .COUT(_12610_),
    .SUM(_12611_));
 sky130_fd_sc_hd__fa_1 _27733_ (.A(_12612_),
    .B(_12613_),
    .CIN(_12614_),
    .COUT(_12615_),
    .SUM(_12616_));
 sky130_fd_sc_hd__fa_1 _27734_ (.A(\hash.CA1.k_i2[18] ),
    .B(\hash.CA1.w_i2[18] ),
    .CIN(_12617_),
    .COUT(_12618_),
    .SUM(_12619_));
 sky130_fd_sc_hd__fa_1 _27735_ (.A(\hash.CA1.k_i2[19] ),
    .B(\hash.CA1.w_i2[19] ),
    .CIN(_12620_),
    .COUT(_12621_),
    .SUM(_12622_));
 sky130_fd_sc_hd__fa_1 _27736_ (.A(\hash.CA1.k_i2[20] ),
    .B(\hash.CA1.w_i2[20] ),
    .CIN(_12623_),
    .COUT(_12624_),
    .SUM(_12625_));
 sky130_fd_sc_hd__fa_1 _27737_ (.A(\hash.CA1.k_i2[21] ),
    .B(\hash.CA1.w_i2[21] ),
    .CIN(_12626_),
    .COUT(_12627_),
    .SUM(_12628_));
 sky130_fd_sc_hd__fa_1 _27738_ (.A(\hash.CA1.k_i2[22] ),
    .B(\hash.CA1.w_i2[22] ),
    .CIN(_12629_),
    .COUT(_12630_),
    .SUM(_12631_));
 sky130_fd_sc_hd__fa_1 _27739_ (.A(_12632_),
    .B(_12633_),
    .CIN(_12634_),
    .COUT(_12635_),
    .SUM(_12636_));
 sky130_fd_sc_hd__fa_1 _27740_ (.A(_12637_),
    .B(_12638_),
    .CIN(_12639_),
    .COUT(_12640_),
    .SUM(_12641_));
 sky130_fd_sc_hd__fa_1 _27741_ (.A(_12642_),
    .B(_12643_),
    .CIN(_12644_),
    .COUT(_12645_),
    .SUM(_12646_));
 sky130_fd_sc_hd__fa_1 _27742_ (.A(_12647_),
    .B(_12648_),
    .CIN(_12649_),
    .COUT(_12650_),
    .SUM(_12651_));
 sky130_fd_sc_hd__fa_1 _27743_ (.A(_12652_),
    .B(_12653_),
    .CIN(_12654_),
    .COUT(_12655_),
    .SUM(_12656_));
 sky130_fd_sc_hd__fa_1 _27744_ (.A(_12657_),
    .B(_12658_),
    .CIN(_12659_),
    .COUT(_12660_),
    .SUM(_12661_));
 sky130_fd_sc_hd__fa_1 _27745_ (.A(\hash.CA1.k_i2[29] ),
    .B(\hash.CA1.w_i2[29] ),
    .CIN(_12662_),
    .COUT(_12663_),
    .SUM(_12664_));
 sky130_fd_sc_hd__fa_1 _27746_ (.A(\hash.CA1.k_i2[30] ),
    .B(\hash.CA1.w_i2[30] ),
    .CIN(_12665_),
    .COUT(_12666_),
    .SUM(_12667_));
 sky130_fd_sc_hd__fa_1 _27747_ (.A(\hash.CA1.k_i1[1] ),
    .B(\hash.CA1.w_i1[1] ),
    .CIN(_12668_),
    .COUT(_12669_),
    .SUM(_12670_));
 sky130_fd_sc_hd__fa_2 _27748_ (.A(_12673_),
    .B(_12672_),
    .CIN(_12671_),
    .COUT(_12674_),
    .SUM(_12675_));
 sky130_fd_sc_hd__fa_1 _27749_ (.A(_12675_),
    .B(_12670_),
    .CIN(_12676_),
    .COUT(_12677_),
    .SUM(_12678_));
 sky130_fd_sc_hd__fa_1 _27750_ (.A(_12679_),
    .B(_12680_),
    .CIN(_12681_),
    .COUT(_12682_),
    .SUM(_12683_));
 sky130_fd_sc_hd__fa_1 _27751_ (.A(_12684_),
    .B(_12685_),
    .CIN(_12686_),
    .COUT(_12687_),
    .SUM(_12688_));
 sky130_fd_sc_hd__fa_1 _27752_ (.A(_12689_),
    .B(_12690_),
    .CIN(_12691_),
    .COUT(_12692_),
    .SUM(_12693_));
 sky130_fd_sc_hd__fa_1 _27753_ (.A(_12694_),
    .B(_12695_),
    .CIN(_12696_),
    .COUT(_12697_),
    .SUM(_12698_));
 sky130_fd_sc_hd__fa_1 _27754_ (.A(_12699_),
    .B(_12700_),
    .CIN(_12701_),
    .COUT(_12702_),
    .SUM(_12703_));
 sky130_fd_sc_hd__fa_1 _27755_ (.A(_12704_),
    .B(_12705_),
    .CIN(_12706_),
    .COUT(_12707_),
    .SUM(_12708_));
 sky130_fd_sc_hd__fa_1 _27756_ (.A(_12709_),
    .B(_12710_),
    .CIN(_12711_),
    .COUT(_12712_),
    .SUM(_12713_));
 sky130_fd_sc_hd__fa_1 _27757_ (.A(_12714_),
    .B(_12715_),
    .CIN(_12716_),
    .COUT(_12717_),
    .SUM(_12718_));
 sky130_fd_sc_hd__fa_1 _27758_ (.A(_12719_),
    .B(_12720_),
    .CIN(_12721_),
    .COUT(_12722_),
    .SUM(_12723_));
 sky130_fd_sc_hd__fa_1 _27759_ (.A(_12724_),
    .B(_12725_),
    .CIN(_12726_),
    .COUT(_12727_),
    .SUM(_12728_));
 sky130_fd_sc_hd__fa_1 _27760_ (.A(_12729_),
    .B(_12730_),
    .CIN(_12731_),
    .COUT(_12732_),
    .SUM(_12733_));
 sky130_fd_sc_hd__fa_1 _27761_ (.A(_12734_),
    .B(_12735_),
    .CIN(_12736_),
    .COUT(_12737_),
    .SUM(_12738_));
 sky130_fd_sc_hd__fa_1 _27762_ (.A(_12740_),
    .B(_12739_),
    .CIN(_12741_),
    .COUT(_12742_),
    .SUM(_12743_));
 sky130_fd_sc_hd__fa_1 _27763_ (.A(_12744_),
    .B(_12745_),
    .CIN(_12746_),
    .COUT(_12747_),
    .SUM(_12748_));
 sky130_fd_sc_hd__fa_1 _27764_ (.A(_12749_),
    .B(_12750_),
    .CIN(_12751_),
    .COUT(_12752_),
    .SUM(_12753_));
 sky130_fd_sc_hd__fa_1 _27765_ (.A(_12756_),
    .B(_12755_),
    .CIN(_12754_),
    .COUT(_12757_),
    .SUM(_12758_));
 sky130_fd_sc_hd__fa_1 _27766_ (.A(_12761_),
    .B(_12760_),
    .CIN(_12759_),
    .COUT(_12762_),
    .SUM(_12763_));
 sky130_fd_sc_hd__fa_1 _27767_ (.A(_12764_),
    .B(_12765_),
    .CIN(_12766_),
    .COUT(_12767_),
    .SUM(_12768_));
 sky130_fd_sc_hd__fa_1 _27768_ (.A(_12769_),
    .B(_12770_),
    .CIN(_12771_),
    .COUT(_12772_),
    .SUM(_12773_));
 sky130_fd_sc_hd__fa_1 _27769_ (.A(_12775_),
    .B(_12774_),
    .CIN(_12776_),
    .COUT(_12777_),
    .SUM(_12778_));
 sky130_fd_sc_hd__fa_1 _27770_ (.A(_12779_),
    .B(_12780_),
    .CIN(_12781_),
    .COUT(_12782_),
    .SUM(_12783_));
 sky130_fd_sc_hd__fa_1 _27771_ (.A(_12786_),
    .B(_12785_),
    .CIN(_12784_),
    .COUT(_12787_),
    .SUM(_12788_));
 sky130_fd_sc_hd__fa_1 _27772_ (.A(_12789_),
    .B(_12790_),
    .CIN(_12791_),
    .COUT(_12792_),
    .SUM(_12793_));
 sky130_fd_sc_hd__fa_1 _27773_ (.A(_12794_),
    .B(_12795_),
    .CIN(_12796_),
    .COUT(_12797_),
    .SUM(_12798_));
 sky130_fd_sc_hd__fa_1 _27774_ (.A(_12799_),
    .B(_12800_),
    .CIN(_12801_),
    .COUT(_12802_),
    .SUM(_12803_));
 sky130_fd_sc_hd__fa_1 _27775_ (.A(_12804_),
    .B(_12805_),
    .CIN(_12806_),
    .COUT(_12807_),
    .SUM(_12808_));
 sky130_fd_sc_hd__fa_1 _27776_ (.A(_12809_),
    .B(_12810_),
    .CIN(_12811_),
    .COUT(_12812_),
    .SUM(_12813_));
 sky130_fd_sc_hd__fa_1 _27777_ (.A(_12814_),
    .B(_12815_),
    .CIN(_12816_),
    .COUT(_12817_),
    .SUM(_12818_));
 sky130_fd_sc_hd__fa_1 _27778_ (.A(_12819_),
    .B(_12820_),
    .CIN(_12821_),
    .COUT(_12822_),
    .SUM(_12823_));
 sky130_fd_sc_hd__fa_1 _27779_ (.A(\hash.CA1.d[0] ),
    .B(_12824_),
    .CIN(_12825_),
    .COUT(_12826_),
    .SUM(_12827_));
 sky130_fd_sc_hd__fa_1 _27780_ (.A(_12828_),
    .B(_12670_),
    .CIN(_12676_),
    .COUT(_12829_),
    .SUM(_12830_));
 sky130_fd_sc_hd__fa_1 _27781_ (.A(_12831_),
    .B(_12832_),
    .CIN(_12833_),
    .COUT(_12834_),
    .SUM(_12835_));
 sky130_fd_sc_hd__fa_1 _27782_ (.A(_12836_),
    .B(_12837_),
    .CIN(_12838_),
    .COUT(_12839_),
    .SUM(_12840_));
 sky130_fd_sc_hd__fa_1 _27783_ (.A(_12841_),
    .B(_12840_),
    .CIN(_12842_),
    .COUT(_12843_),
    .SUM(_12844_));
 sky130_fd_sc_hd__fa_1 _27784_ (.A(_12685_),
    .B(_12845_),
    .CIN(_12686_),
    .COUT(_12846_),
    .SUM(_12847_));
 sky130_fd_sc_hd__fa_1 _27785_ (.A(_12839_),
    .B(_12847_),
    .CIN(_12684_),
    .COUT(_12848_),
    .SUM(_12849_));
 sky130_fd_sc_hd__fa_1 _27786_ (.A(_12690_),
    .B(_12850_),
    .CIN(_12691_),
    .COUT(_12851_),
    .SUM(_12852_));
 sky130_fd_sc_hd__fa_1 _27787_ (.A(_12846_),
    .B(_12852_),
    .CIN(_12689_),
    .COUT(_12853_),
    .SUM(_12854_));
 sky130_fd_sc_hd__fa_1 _27788_ (.A(_12695_),
    .B(_12855_),
    .CIN(_12696_),
    .COUT(_12856_),
    .SUM(_12857_));
 sky130_fd_sc_hd__fa_1 _27789_ (.A(_12851_),
    .B(_12858_),
    .CIN(_12859_),
    .COUT(_12860_),
    .SUM(_12861_));
 sky130_fd_sc_hd__fa_1 _27790_ (.A(_12862_),
    .B(_12863_),
    .CIN(_12864_),
    .COUT(_12865_),
    .SUM(_12866_));
 sky130_fd_sc_hd__fa_1 _27791_ (.A(_12867_),
    .B(_12866_),
    .CIN(_12868_),
    .COUT(_12869_),
    .SUM(_12870_));
 sky130_fd_sc_hd__fa_1 _27792_ (.A(_12871_),
    .B(_12872_),
    .CIN(_12873_),
    .COUT(_12874_),
    .SUM(_12875_));
 sky130_fd_sc_hd__fa_1 _27793_ (.A(_12865_),
    .B(_12875_),
    .CIN(_12876_),
    .COUT(_12877_),
    .SUM(_12878_));
 sky130_fd_sc_hd__fa_1 _27794_ (.A(_12710_),
    .B(_12879_),
    .CIN(_12711_),
    .COUT(_12880_),
    .SUM(_12881_));
 sky130_fd_sc_hd__fa_1 _27795_ (.A(_12874_),
    .B(_12881_),
    .CIN(_12709_),
    .COUT(_12882_),
    .SUM(_12883_));
 sky130_fd_sc_hd__fa_1 _27796_ (.A(_12884_),
    .B(_12885_),
    .CIN(_12886_),
    .COUT(_12887_),
    .SUM(_12888_));
 sky130_fd_sc_hd__fa_1 _27797_ (.A(_12889_),
    .B(_12890_),
    .CIN(_12891_),
    .COUT(_12892_),
    .SUM(_12893_));
 sky130_fd_sc_hd__fa_1 _27798_ (.A(_12720_),
    .B(_12894_),
    .CIN(_12721_),
    .COUT(_12895_),
    .SUM(_12896_));
 sky130_fd_sc_hd__fa_1 _27799_ (.A(_12897_),
    .B(_12899_),
    .CIN(_12898_),
    .COUT(_12900_),
    .SUM(_12901_));
 sky130_fd_sc_hd__fa_1 _27800_ (.A(_12902_),
    .B(_12903_),
    .CIN(_12904_),
    .COUT(_12905_),
    .SUM(_12906_));
 sky130_fd_sc_hd__fa_1 _27801_ (.A(_12907_),
    .B(_12906_),
    .CIN(_12908_),
    .COUT(_12909_),
    .SUM(_12910_));
 sky130_fd_sc_hd__fa_1 _27802_ (.A(_12730_),
    .B(_12911_),
    .CIN(_12731_),
    .COUT(_12912_),
    .SUM(_12913_));
 sky130_fd_sc_hd__fa_1 _27803_ (.A(_12905_),
    .B(_12914_),
    .CIN(_12913_),
    .COUT(_12915_),
    .SUM(_12916_));
 sky130_fd_sc_hd__fa_1 _27804_ (.A(_12735_),
    .B(_12917_),
    .CIN(_12736_),
    .COUT(_12918_),
    .SUM(_12919_));
 sky130_fd_sc_hd__fa_1 _27805_ (.A(_12912_),
    .B(_12919_),
    .CIN(_12920_),
    .COUT(_12921_),
    .SUM(_12922_));
 sky130_fd_sc_hd__fa_1 _27806_ (.A(_12740_),
    .B(_12923_),
    .CIN(_12741_),
    .COUT(_12924_),
    .SUM(_12925_));
 sky130_fd_sc_hd__fa_1 _27807_ (.A(_12918_),
    .B(_12926_),
    .CIN(_12927_),
    .COUT(_12928_),
    .SUM(_12929_));
 sky130_fd_sc_hd__fa_1 _27808_ (.A(_12745_),
    .B(_12930_),
    .CIN(_12746_),
    .COUT(_12931_),
    .SUM(_12932_));
 sky130_fd_sc_hd__fa_1 _27809_ (.A(_12933_),
    .B(_12934_),
    .CIN(_12935_),
    .COUT(_12936_),
    .SUM(_12937_));
 sky130_fd_sc_hd__fa_1 _27810_ (.A(_12750_),
    .B(_12938_),
    .CIN(_12751_),
    .COUT(_12939_),
    .SUM(_12940_));
 sky130_fd_sc_hd__fa_1 _27811_ (.A(_12941_),
    .B(_12940_),
    .CIN(_12942_),
    .COUT(_12943_),
    .SUM(_12944_));
 sky130_fd_sc_hd__fa_1 _27812_ (.A(_12755_),
    .B(_12945_),
    .CIN(_12756_),
    .COUT(_12946_),
    .SUM(_12947_));
 sky130_fd_sc_hd__fa_1 _27813_ (.A(_12939_),
    .B(_12947_),
    .CIN(_12948_),
    .COUT(_12949_),
    .SUM(_12950_));
 sky130_fd_sc_hd__fa_1 _27814_ (.A(_12760_),
    .B(_12951_),
    .CIN(_12761_),
    .COUT(_12952_),
    .SUM(_12953_));
 sky130_fd_sc_hd__fa_1 _27815_ (.A(_12946_),
    .B(_12953_),
    .CIN(_12954_),
    .COUT(_12955_),
    .SUM(_12956_));
 sky130_fd_sc_hd__fa_1 _27816_ (.A(_12765_),
    .B(_12957_),
    .CIN(_12766_),
    .COUT(_12958_),
    .SUM(_12959_));
 sky130_fd_sc_hd__fa_1 _27817_ (.A(_12952_),
    .B(_12959_),
    .CIN(_12960_),
    .COUT(_12961_),
    .SUM(_12962_));
 sky130_fd_sc_hd__fa_1 _27818_ (.A(_12963_),
    .B(_12964_),
    .CIN(_12965_),
    .COUT(_12966_),
    .SUM(_12967_));
 sky130_fd_sc_hd__fa_1 _27819_ (.A(_12958_),
    .B(_12968_),
    .CIN(_12969_),
    .COUT(_12970_),
    .SUM(_12971_));
 sky130_fd_sc_hd__fa_1 _27820_ (.A(_12972_),
    .B(_12973_),
    .CIN(_12974_),
    .COUT(_12975_),
    .SUM(_12976_));
 sky130_fd_sc_hd__fa_1 _27821_ (.A(_12977_),
    .B(_12976_),
    .CIN(_12978_),
    .COUT(_12979_),
    .SUM(_12980_));
 sky130_fd_sc_hd__fa_1 _27822_ (.A(_12780_),
    .B(_12981_),
    .CIN(_12781_),
    .COUT(_12982_),
    .SUM(_12983_));
 sky130_fd_sc_hd__fa_1 _27823_ (.A(_12975_),
    .B(_12984_),
    .CIN(_12985_),
    .COUT(_12986_),
    .SUM(_12987_));
 sky130_fd_sc_hd__fa_1 _27824_ (.A(_12988_),
    .B(_12989_),
    .CIN(_12990_),
    .COUT(_12991_),
    .SUM(_12992_));
 sky130_fd_sc_hd__fa_1 _27825_ (.A(_12993_),
    .B(_12992_),
    .CIN(_12994_),
    .COUT(_12995_),
    .SUM(_12996_));
 sky130_fd_sc_hd__fa_1 _27826_ (.A(_12790_),
    .B(_12997_),
    .CIN(_12791_),
    .COUT(_12998_),
    .SUM(_12999_));
 sky130_fd_sc_hd__fa_1 _27827_ (.A(_12991_),
    .B(_13000_),
    .CIN(_13001_),
    .COUT(_13002_),
    .SUM(_13003_));
 sky130_fd_sc_hd__fa_1 _27828_ (.A(_13004_),
    .B(_13005_),
    .CIN(_13006_),
    .COUT(_13007_),
    .SUM(_13008_));
 sky130_fd_sc_hd__fa_1 _27829_ (.A(_13009_),
    .B(_13008_),
    .CIN(_13010_),
    .COUT(_13011_),
    .SUM(_13012_));
 sky130_fd_sc_hd__fa_1 _27830_ (.A(_12800_),
    .B(_13013_),
    .CIN(_12801_),
    .COUT(_13014_),
    .SUM(_13015_));
 sky130_fd_sc_hd__fa_1 _27831_ (.A(_13007_),
    .B(_13015_),
    .CIN(_13016_),
    .COUT(_13017_),
    .SUM(_13018_));
 sky130_fd_sc_hd__fa_1 _27832_ (.A(_13019_),
    .B(_13020_),
    .CIN(_13021_),
    .COUT(_13022_),
    .SUM(_13023_));
 sky130_fd_sc_hd__fa_1 _27833_ (.A(_13014_),
    .B(_13023_),
    .CIN(_13024_),
    .COUT(_13025_),
    .SUM(_13026_));
 sky130_fd_sc_hd__fa_1 _27834_ (.A(_13027_),
    .B(_13028_),
    .CIN(_13029_),
    .COUT(_13030_),
    .SUM(_13031_));
 sky130_fd_sc_hd__fa_1 _27835_ (.A(_13022_),
    .B(_13031_),
    .CIN(_13032_),
    .COUT(_13033_),
    .SUM(_13034_));
 sky130_fd_sc_hd__fa_1 _27836_ (.A(_12815_),
    .B(_13035_),
    .CIN(_12816_),
    .COUT(_13036_),
    .SUM(_13037_));
 sky130_fd_sc_hd__fa_1 _27837_ (.A(_13030_),
    .B(_13037_),
    .CIN(_13038_),
    .COUT(_13039_),
    .SUM(_13040_));
 sky130_fd_sc_hd__fa_1 _27838_ (.A(_13041_),
    .B(_13042_),
    .CIN(_13043_),
    .COUT(_13044_),
    .SUM(_13045_));
 sky130_fd_sc_hd__fa_1 _27839_ (.A(_13046_),
    .B(_13047_),
    .CIN(_12819_),
    .COUT(_13048_),
    .SUM(_13049_));
 sky130_fd_sc_hd__fa_1 _27840_ (.A(_13050_),
    .B(_13051_),
    .CIN(_13052_),
    .COUT(_13053_),
    .SUM(\hash.CA1.p1[1] ));
 sky130_fd_sc_hd__fa_1 _27841_ (.A(_13054_),
    .B(_12834_),
    .CIN(_12844_),
    .COUT(_13055_),
    .SUM(\hash.CA1.p2[2] ));
 sky130_fd_sc_hd__fa_1 _27842_ (.A(_12824_),
    .B(_13056_),
    .CIN(_12825_),
    .COUT(_13057_),
    .SUM(_13058_));
 sky130_fd_sc_hd__fa_1 _27843_ (.A(_13059_),
    .B(_13060_),
    .CIN(_13061_),
    .COUT(_13062_),
    .SUM(\hash.CA1.p3[2] ));
 sky130_fd_sc_hd__fa_1 _27844_ (.A(_00721_),
    .B(_13063_),
    .CIN(_13064_),
    .COUT(_13065_),
    .SUM(\hash.CA1.p5[1] ));
 sky130_fd_sc_hd__ha_4 _27845_ (.A(_00656_),
    .B(_13068_),
    .COUT(_13069_),
    .SUM(_00657_));
 sky130_fd_sc_hd__ha_4 _27846_ (.A(_00656_),
    .B(\count_hash2[2] ),
    .COUT(_13070_),
    .SUM(_13071_));
 sky130_fd_sc_hd__ha_4 _27847_ (.A(\count_hash2[1] ),
    .B(_13068_),
    .COUT(_13072_),
    .SUM(_13073_));
 sky130_fd_sc_hd__ha_4 _27848_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_13074_),
    .SUM(_13075_));
 sky130_fd_sc_hd__ha_4 _27849_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_13076_),
    .SUM(_13077_));
 sky130_fd_sc_hd__ha_4 _27850_ (.A(_00642_),
    .B(_13078_),
    .COUT(_13079_),
    .SUM(_00655_));
 sky130_fd_sc_hd__ha_4 _27851_ (.A(_00642_),
    .B(\count_hash1[2] ),
    .COUT(_13080_),
    .SUM(_13081_));
 sky130_fd_sc_hd__ha_1 _27852_ (.A(_00642_),
    .B(\count_hash1[2] ),
    .COUT(_13082_),
    .SUM(_13083_));
 sky130_fd_sc_hd__ha_4 _27853_ (.A(\count_hash1[1] ),
    .B(_13078_),
    .COUT(_13084_),
    .SUM(_13085_));
 sky130_fd_sc_hd__ha_4 _27854_ (.A(\count_hash1[1] ),
    .B(\count_hash1[2] ),
    .COUT(_13086_),
    .SUM(_13087_));
 sky130_fd_sc_hd__ha_4 _27855_ (.A(\count_hash1[1] ),
    .B(\count_hash1[2] ),
    .COUT(_13088_),
    .SUM(_13089_));
 sky130_fd_sc_hd__ha_4 _27856_ (.A(\hash.CA2.p1[0] ),
    .B(\hash.CA2.p3[0] ),
    .COUT(_12251_),
    .SUM(_13090_));
 sky130_fd_sc_hd__ha_4 _27857_ (.A(\hash.CA2.p1[2] ),
    .B(\hash.CA2.p3[2] ),
    .COUT(_13091_),
    .SUM(_13092_));
 sky130_fd_sc_hd__ha_1 _27858_ (.A(\hash.CA2.p1[1] ),
    .B(\hash.CA2.p3[1] ),
    .COUT(_13093_),
    .SUM(_13094_));
 sky130_fd_sc_hd__ha_2 _27859_ (.A(\hash.CA2.p1[7] ),
    .B(\hash.CA2.p3[7] ),
    .COUT(_13095_),
    .SUM(_13096_));
 sky130_fd_sc_hd__ha_2 _27860_ (.A(\hash.CA2.p1[6] ),
    .B(\hash.CA2.p3[6] ),
    .COUT(_13097_),
    .SUM(_13098_));
 sky130_fd_sc_hd__ha_2 _27861_ (.A(\hash.CA2.p1[5] ),
    .B(\hash.CA2.p3[5] ),
    .COUT(_13099_),
    .SUM(_13100_));
 sky130_fd_sc_hd__ha_2 _27862_ (.A(\hash.CA2.p1[4] ),
    .B(\hash.CA2.p3[4] ),
    .COUT(_13101_),
    .SUM(_13102_));
 sky130_fd_sc_hd__ha_2 _27863_ (.A(\hash.CA2.p1[3] ),
    .B(\hash.CA2.p3[3] ),
    .COUT(_13103_),
    .SUM(_13104_));
 sky130_fd_sc_hd__ha_2 _27864_ (.A(\hash.CA2.p1[9] ),
    .B(\hash.CA2.p3[9] ),
    .COUT(_13105_),
    .SUM(_13106_));
 sky130_fd_sc_hd__ha_4 _27865_ (.A(\hash.CA2.p1[8] ),
    .B(\hash.CA2.p3[8] ),
    .COUT(_13107_),
    .SUM(_13108_));
 sky130_fd_sc_hd__ha_2 _27866_ (.A(\hash.CA2.p1[10] ),
    .B(\hash.CA2.p3[10] ),
    .COUT(_13109_),
    .SUM(_13110_));
 sky130_fd_sc_hd__ha_2 _27867_ (.A(\hash.CA2.p1[11] ),
    .B(\hash.CA2.p3[11] ),
    .COUT(_13111_),
    .SUM(_13112_));
 sky130_fd_sc_hd__ha_4 _27868_ (.A(\hash.CA2.p1[13] ),
    .B(\hash.CA2.p3[13] ),
    .COUT(_13113_),
    .SUM(_13114_));
 sky130_fd_sc_hd__ha_2 _27869_ (.A(\hash.CA2.p1[12] ),
    .B(\hash.CA2.p3[12] ),
    .COUT(_13115_),
    .SUM(_13116_));
 sky130_fd_sc_hd__ha_2 _27870_ (.A(\hash.CA2.p1[15] ),
    .B(\hash.CA2.p3[15] ),
    .COUT(_13117_),
    .SUM(_13118_));
 sky130_fd_sc_hd__ha_2 _27871_ (.A(\hash.CA2.p1[14] ),
    .B(\hash.CA2.p3[14] ),
    .COUT(_13119_),
    .SUM(_13120_));
 sky130_fd_sc_hd__ha_2 _27872_ (.A(\hash.CA2.p1[16] ),
    .B(\hash.CA2.p3[16] ),
    .COUT(_13121_),
    .SUM(_13122_));
 sky130_fd_sc_hd__ha_4 _27873_ (.A(\hash.CA2.p1[17] ),
    .B(\hash.CA2.p3[17] ),
    .COUT(_13123_),
    .SUM(_13124_));
 sky130_fd_sc_hd__ha_2 _27874_ (.A(\hash.CA2.p1[18] ),
    .B(\hash.CA2.p3[18] ),
    .COUT(_13125_),
    .SUM(_13126_));
 sky130_fd_sc_hd__ha_2 _27875_ (.A(\hash.CA2.p1[21] ),
    .B(\hash.CA2.p3[21] ),
    .COUT(_13127_),
    .SUM(_13128_));
 sky130_fd_sc_hd__ha_1 _27876_ (.A(\hash.CA2.p1[20] ),
    .B(\hash.CA2.p3[20] ),
    .COUT(_13129_),
    .SUM(_13130_));
 sky130_fd_sc_hd__ha_4 _27877_ (.A(\hash.CA2.p1[19] ),
    .B(\hash.CA2.p3[19] ),
    .COUT(_13131_),
    .SUM(_13132_));
 sky130_fd_sc_hd__ha_4 _27878_ (.A(\hash.CA2.p1[22] ),
    .B(\hash.CA2.p3[22] ),
    .COUT(_13133_),
    .SUM(_13134_));
 sky130_fd_sc_hd__ha_2 _27879_ (.A(\hash.CA2.p1[24] ),
    .B(\hash.CA2.p3[24] ),
    .COUT(_13135_),
    .SUM(_13136_));
 sky130_fd_sc_hd__ha_2 _27880_ (.A(\hash.CA2.p1[23] ),
    .B(\hash.CA2.p3[23] ),
    .COUT(_13137_),
    .SUM(_13138_));
 sky130_fd_sc_hd__ha_2 _27881_ (.A(\hash.CA2.p1[25] ),
    .B(\hash.CA2.p3[25] ),
    .COUT(_13139_),
    .SUM(_13140_));
 sky130_fd_sc_hd__ha_2 _27882_ (.A(\hash.CA2.p1[27] ),
    .B(\hash.CA2.p3[27] ),
    .COUT(_13141_),
    .SUM(_13142_));
 sky130_fd_sc_hd__ha_2 _27883_ (.A(\hash.CA2.p1[26] ),
    .B(\hash.CA2.p3[26] ),
    .COUT(_13143_),
    .SUM(_13144_));
 sky130_fd_sc_hd__ha_2 _27884_ (.A(\hash.CA2.p1[28] ),
    .B(\hash.CA2.p3[28] ),
    .COUT(_13145_),
    .SUM(_13146_));
 sky130_fd_sc_hd__ha_2 _27885_ (.A(\hash.CA2.p1[29] ),
    .B(\hash.CA2.p3[29] ),
    .COUT(_13147_),
    .SUM(_13148_));
 sky130_fd_sc_hd__ha_1 _27886_ (.A(\hash.CA2.p1[30] ),
    .B(\hash.CA2.p3[30] ),
    .COUT(_13149_),
    .SUM(_13150_));
 sky130_fd_sc_hd__ha_1 _27887_ (.A(_13151_),
    .B(_13152_),
    .COUT(_13153_),
    .SUM(_13154_));
 sky130_fd_sc_hd__ha_1 _27888_ (.A(_13153_),
    .B(_13155_),
    .COUT(_13156_),
    .SUM(_13157_));
 sky130_fd_sc_hd__ha_1 _27889_ (.A(_13158_),
    .B(_13159_),
    .COUT(_13160_),
    .SUM(_13161_));
 sky130_fd_sc_hd__ha_1 _27890_ (.A(_13162_),
    .B(_13163_),
    .COUT(_13164_),
    .SUM(_13165_));
 sky130_fd_sc_hd__ha_1 _27891_ (.A(_13166_),
    .B(_13167_),
    .COUT(_13168_),
    .SUM(_13169_));
 sky130_fd_sc_hd__ha_1 _27892_ (.A(_13170_),
    .B(_13171_),
    .COUT(_13172_),
    .SUM(_13173_));
 sky130_fd_sc_hd__ha_1 _27893_ (.A(_13174_),
    .B(_13175_),
    .COUT(_13176_),
    .SUM(_13177_));
 sky130_fd_sc_hd__ha_4 _27894_ (.A(_13178_),
    .B(_13179_),
    .COUT(_13180_),
    .SUM(_13181_));
 sky130_fd_sc_hd__ha_1 _27895_ (.A(_13182_),
    .B(_13183_),
    .COUT(_13184_),
    .SUM(_13185_));
 sky130_fd_sc_hd__ha_2 _27896_ (.A(_13186_),
    .B(_13187_),
    .COUT(_13188_),
    .SUM(_13189_));
 sky130_fd_sc_hd__ha_2 _27897_ (.A(_13190_),
    .B(_13191_),
    .COUT(_13192_),
    .SUM(_13193_));
 sky130_fd_sc_hd__ha_1 _27898_ (.A(_13194_),
    .B(_13195_),
    .COUT(_13196_),
    .SUM(_13197_));
 sky130_fd_sc_hd__ha_1 _27899_ (.A(_13198_),
    .B(_13199_),
    .COUT(_13200_),
    .SUM(_13201_));
 sky130_fd_sc_hd__ha_1 _27900_ (.A(_13202_),
    .B(_13203_),
    .COUT(_13204_),
    .SUM(_13205_));
 sky130_fd_sc_hd__ha_1 _27901_ (.A(_13206_),
    .B(_13207_),
    .COUT(_13208_),
    .SUM(_13209_));
 sky130_fd_sc_hd__ha_2 _27902_ (.A(_13210_),
    .B(_13211_),
    .COUT(_13212_),
    .SUM(_13213_));
 sky130_fd_sc_hd__ha_2 _27903_ (.A(_13214_),
    .B(_13215_),
    .COUT(_13216_),
    .SUM(_13217_));
 sky130_fd_sc_hd__ha_2 _27904_ (.A(_13218_),
    .B(_13219_),
    .COUT(_13220_),
    .SUM(_13221_));
 sky130_fd_sc_hd__ha_1 _27905_ (.A(_13222_),
    .B(_13223_),
    .COUT(_13224_),
    .SUM(_13225_));
 sky130_fd_sc_hd__ha_2 _27906_ (.A(_13226_),
    .B(_13227_),
    .COUT(_13228_),
    .SUM(_13229_));
 sky130_fd_sc_hd__ha_2 _27907_ (.A(_13230_),
    .B(_13231_),
    .COUT(_13232_),
    .SUM(_13233_));
 sky130_fd_sc_hd__ha_1 _27908_ (.A(_13234_),
    .B(_13235_),
    .COUT(_13236_),
    .SUM(_13237_));
 sky130_fd_sc_hd__ha_1 _27909_ (.A(_13238_),
    .B(_13239_),
    .COUT(_13240_),
    .SUM(_13241_));
 sky130_fd_sc_hd__ha_1 _27910_ (.A(_13242_),
    .B(_13243_),
    .COUT(_13244_),
    .SUM(_13245_));
 sky130_fd_sc_hd__ha_1 _27911_ (.A(_13246_),
    .B(_13247_),
    .COUT(_13248_),
    .SUM(_13249_));
 sky130_fd_sc_hd__ha_1 _27912_ (.A(_13250_),
    .B(_13251_),
    .COUT(_13252_),
    .SUM(_13253_));
 sky130_fd_sc_hd__ha_1 _27913_ (.A(_13254_),
    .B(_13255_),
    .COUT(_13256_),
    .SUM(_13257_));
 sky130_fd_sc_hd__ha_1 _27914_ (.A(_13258_),
    .B(_13259_),
    .COUT(_13260_),
    .SUM(_13261_));
 sky130_fd_sc_hd__ha_2 _27915_ (.A(_13262_),
    .B(_13263_),
    .COUT(_13264_),
    .SUM(_13265_));
 sky130_fd_sc_hd__ha_1 _27916_ (.A(_13266_),
    .B(_13267_),
    .COUT(_13268_),
    .SUM(_13269_));
 sky130_fd_sc_hd__ha_2 _27917_ (.A(_13270_),
    .B(_13271_),
    .COUT(_13272_),
    .SUM(_13273_));
 sky130_fd_sc_hd__ha_1 _27918_ (.A(_13274_),
    .B(_13275_),
    .COUT(_13276_),
    .SUM(_13277_));
 sky130_fd_sc_hd__ha_1 _27919_ (.A(_13276_),
    .B(_13278_),
    .COUT(_13279_),
    .SUM(_13280_));
 sky130_fd_sc_hd__ha_1 _27920_ (.A(_13281_),
    .B(_13282_),
    .COUT(_13283_),
    .SUM(_13284_));
 sky130_fd_sc_hd__ha_1 _27921_ (.A(_13285_),
    .B(_13286_),
    .COUT(_13287_),
    .SUM(_13288_));
 sky130_fd_sc_hd__ha_1 _27922_ (.A(_13289_),
    .B(_13290_),
    .COUT(_13291_),
    .SUM(_13292_));
 sky130_fd_sc_hd__ha_1 _27923_ (.A(_13293_),
    .B(_13294_),
    .COUT(_13295_),
    .SUM(_13296_));
 sky130_fd_sc_hd__ha_1 _27924_ (.A(_13297_),
    .B(_13298_),
    .COUT(_13299_),
    .SUM(_13300_));
 sky130_fd_sc_hd__ha_2 _27925_ (.A(_13301_),
    .B(_13302_),
    .COUT(_13303_),
    .SUM(_13304_));
 sky130_fd_sc_hd__ha_1 _27926_ (.A(_13305_),
    .B(_13306_),
    .COUT(_13307_),
    .SUM(_13308_));
 sky130_fd_sc_hd__ha_1 _27927_ (.A(_13309_),
    .B(_13310_),
    .COUT(_13311_),
    .SUM(_13312_));
 sky130_fd_sc_hd__ha_1 _27928_ (.A(_13313_),
    .B(_13314_),
    .COUT(_13315_),
    .SUM(_13316_));
 sky130_fd_sc_hd__ha_1 _27929_ (.A(_13317_),
    .B(_13318_),
    .COUT(_13319_),
    .SUM(_13320_));
 sky130_fd_sc_hd__ha_1 _27930_ (.A(_13321_),
    .B(_13322_),
    .COUT(_13323_),
    .SUM(_13324_));
 sky130_fd_sc_hd__ha_1 _27931_ (.A(_13325_),
    .B(_13326_),
    .COUT(_13327_),
    .SUM(_13328_));
 sky130_fd_sc_hd__ha_1 _27932_ (.A(_13329_),
    .B(_13330_),
    .COUT(_13331_),
    .SUM(_13332_));
 sky130_fd_sc_hd__ha_1 _27933_ (.A(_13333_),
    .B(_13334_),
    .COUT(_13335_),
    .SUM(_13336_));
 sky130_fd_sc_hd__ha_1 _27934_ (.A(_13337_),
    .B(_13338_),
    .COUT(_13339_),
    .SUM(_13340_));
 sky130_fd_sc_hd__ha_2 _27935_ (.A(_13341_),
    .B(_13342_),
    .COUT(_13343_),
    .SUM(_13344_));
 sky130_fd_sc_hd__ha_1 _27936_ (.A(_13345_),
    .B(_13346_),
    .COUT(_13347_),
    .SUM(_13348_));
 sky130_fd_sc_hd__ha_1 _27937_ (.A(_13349_),
    .B(_13350_),
    .COUT(_13351_),
    .SUM(_13352_));
 sky130_fd_sc_hd__ha_2 _27938_ (.A(_13353_),
    .B(_13354_),
    .COUT(_13355_),
    .SUM(_13356_));
 sky130_fd_sc_hd__ha_1 _27939_ (.A(_13357_),
    .B(_13358_),
    .COUT(_13359_),
    .SUM(_13360_));
 sky130_fd_sc_hd__ha_2 _27940_ (.A(_13361_),
    .B(_13362_),
    .COUT(_13363_),
    .SUM(_13364_));
 sky130_fd_sc_hd__ha_1 _27941_ (.A(_13365_),
    .B(_13366_),
    .COUT(_13367_),
    .SUM(_13368_));
 sky130_fd_sc_hd__ha_2 _27942_ (.A(_13369_),
    .B(_13370_),
    .COUT(_13371_),
    .SUM(_13372_));
 sky130_fd_sc_hd__ha_1 _27943_ (.A(_13373_),
    .B(_13374_),
    .COUT(_13375_),
    .SUM(_13376_));
 sky130_fd_sc_hd__ha_2 _27944_ (.A(_13377_),
    .B(_13378_),
    .COUT(_13379_),
    .SUM(_13380_));
 sky130_fd_sc_hd__ha_1 _27945_ (.A(_13381_),
    .B(_13382_),
    .COUT(_13383_),
    .SUM(_13384_));
 sky130_fd_sc_hd__ha_1 _27946_ (.A(_13385_),
    .B(_13386_),
    .COUT(_13387_),
    .SUM(_13388_));
 sky130_fd_sc_hd__ha_2 _27947_ (.A(_13389_),
    .B(_13390_),
    .COUT(_13391_),
    .SUM(_13392_));
 sky130_fd_sc_hd__ha_1 _27948_ (.A(_13393_),
    .B(_13394_),
    .COUT(_13395_),
    .SUM(_13396_));
 sky130_fd_sc_hd__ha_2 _27949_ (.A(_13397_),
    .B(_13398_),
    .COUT(_13399_),
    .SUM(_13400_));
 sky130_fd_sc_hd__ha_4 _27950_ (.A(\hash.CA2.p4[0] ),
    .B(_13401_),
    .COUT(_13402_),
    .SUM(_13403_));
 sky130_fd_sc_hd__ha_1 _27951_ (.A(_13404_),
    .B(_13405_),
    .COUT(_13406_),
    .SUM(_13407_));
 sky130_fd_sc_hd__ha_4 _27952_ (.A(_13402_),
    .B(_12267_),
    .COUT(_13408_),
    .SUM(_13409_));
 sky130_fd_sc_hd__ha_1 _27953_ (.A(_13410_),
    .B(_13411_),
    .COUT(_13412_),
    .SUM(_13413_));
 sky130_fd_sc_hd__ha_1 _27954_ (.A(_12266_),
    .B(_12276_),
    .COUT(_13415_),
    .SUM(_13416_));
 sky130_fd_sc_hd__ha_1 _27955_ (.A(_13417_),
    .B(_13418_),
    .COUT(_13419_),
    .SUM(_13420_));
 sky130_fd_sc_hd__ha_2 _27956_ (.A(_12275_),
    .B(_12290_),
    .COUT(_13422_),
    .SUM(_13423_));
 sky130_fd_sc_hd__ha_1 _27957_ (.A(_13424_),
    .B(_13425_),
    .COUT(_13426_),
    .SUM(_13427_));
 sky130_fd_sc_hd__ha_2 _27958_ (.A(_12289_),
    .B(_12299_),
    .COUT(_13429_),
    .SUM(_13430_));
 sky130_fd_sc_hd__ha_1 _27959_ (.A(_13431_),
    .B(_13432_),
    .COUT(_13433_),
    .SUM(_13434_));
 sky130_fd_sc_hd__ha_1 _27960_ (.A(_12298_),
    .B(_12308_),
    .COUT(_13436_),
    .SUM(_13437_));
 sky130_fd_sc_hd__ha_1 _27961_ (.A(_13438_),
    .B(_13439_),
    .COUT(_13440_),
    .SUM(_13441_));
 sky130_fd_sc_hd__ha_4 _27962_ (.A(_12307_),
    .B(_12317_),
    .COUT(_13443_),
    .SUM(_13444_));
 sky130_fd_sc_hd__ha_1 _27963_ (.A(_13445_),
    .B(_13446_),
    .COUT(_13447_),
    .SUM(_13448_));
 sky130_fd_sc_hd__ha_1 _27964_ (.A(_12316_),
    .B(_12326_),
    .COUT(_13450_),
    .SUM(_13451_));
 sky130_fd_sc_hd__ha_1 _27965_ (.A(_13452_),
    .B(_13453_),
    .COUT(_13454_),
    .SUM(_13455_));
 sky130_fd_sc_hd__ha_4 _27966_ (.A(_12325_),
    .B(_12335_),
    .COUT(_13457_),
    .SUM(_13458_));
 sky130_fd_sc_hd__ha_1 _27967_ (.A(_13459_),
    .B(_13460_),
    .COUT(_13461_),
    .SUM(_13462_));
 sky130_fd_sc_hd__ha_2 _27968_ (.A(_12334_),
    .B(_12344_),
    .COUT(_13464_),
    .SUM(_13465_));
 sky130_fd_sc_hd__ha_1 _27969_ (.A(_13466_),
    .B(_13467_),
    .COUT(_13468_),
    .SUM(_13469_));
 sky130_fd_sc_hd__ha_2 _27970_ (.A(_12343_),
    .B(_12353_),
    .COUT(_13471_),
    .SUM(_13472_));
 sky130_fd_sc_hd__ha_2 _27971_ (.A(_13473_),
    .B(_13474_),
    .COUT(_13475_),
    .SUM(_13476_));
 sky130_fd_sc_hd__ha_2 _27972_ (.A(_12352_),
    .B(_12362_),
    .COUT(_13478_),
    .SUM(_13479_));
 sky130_fd_sc_hd__ha_1 _27973_ (.A(_13480_),
    .B(_13481_),
    .COUT(_13482_),
    .SUM(_13483_));
 sky130_fd_sc_hd__ha_2 _27974_ (.A(_12361_),
    .B(_12371_),
    .COUT(_13485_),
    .SUM(_13486_));
 sky130_fd_sc_hd__ha_1 _27975_ (.A(_13487_),
    .B(_13488_),
    .COUT(_13489_),
    .SUM(_13490_));
 sky130_fd_sc_hd__ha_4 _27976_ (.A(_12380_),
    .B(_12370_),
    .COUT(_13492_),
    .SUM(_13493_));
 sky130_fd_sc_hd__ha_2 _27977_ (.A(_13495_),
    .B(_13494_),
    .COUT(_13496_),
    .SUM(_13497_));
 sky130_fd_sc_hd__ha_2 _27978_ (.A(_12379_),
    .B(_12389_),
    .COUT(_13499_),
    .SUM(_13500_));
 sky130_fd_sc_hd__ha_1 _27979_ (.A(_13501_),
    .B(_13502_),
    .COUT(_13503_),
    .SUM(_13504_));
 sky130_fd_sc_hd__ha_1 _27980_ (.A(_12388_),
    .B(_12398_),
    .COUT(_13506_),
    .SUM(_13507_));
 sky130_fd_sc_hd__ha_1 _27981_ (.A(_13508_),
    .B(_13509_),
    .COUT(_13510_),
    .SUM(_13511_));
 sky130_fd_sc_hd__ha_1 _27982_ (.A(_12397_),
    .B(_12407_),
    .COUT(_13513_),
    .SUM(_13514_));
 sky130_fd_sc_hd__ha_1 _27983_ (.A(_13515_),
    .B(_13516_),
    .COUT(_13517_),
    .SUM(_13518_));
 sky130_fd_sc_hd__ha_1 _27984_ (.A(_12406_),
    .B(_12416_),
    .COUT(_13520_),
    .SUM(_13521_));
 sky130_fd_sc_hd__ha_1 _27985_ (.A(_13522_),
    .B(_13523_),
    .COUT(_13524_),
    .SUM(_13525_));
 sky130_fd_sc_hd__ha_1 _27986_ (.A(_12415_),
    .B(_12425_),
    .COUT(_13527_),
    .SUM(_13528_));
 sky130_fd_sc_hd__ha_1 _27987_ (.A(_13529_),
    .B(_13530_),
    .COUT(_13531_),
    .SUM(_13532_));
 sky130_fd_sc_hd__ha_1 _27988_ (.A(_12424_),
    .B(_12434_),
    .COUT(_13534_),
    .SUM(_13535_));
 sky130_fd_sc_hd__ha_1 _27989_ (.A(_13536_),
    .B(_13537_),
    .COUT(_13538_),
    .SUM(_13539_));
 sky130_fd_sc_hd__ha_1 _27990_ (.A(_12433_),
    .B(_12443_),
    .COUT(_13541_),
    .SUM(_13542_));
 sky130_fd_sc_hd__ha_1 _27991_ (.A(_13543_),
    .B(_13544_),
    .COUT(_13545_),
    .SUM(_13546_));
 sky130_fd_sc_hd__ha_2 _27992_ (.A(_12442_),
    .B(_12452_),
    .COUT(_13548_),
    .SUM(_13549_));
 sky130_fd_sc_hd__ha_2 _27993_ (.A(_13550_),
    .B(_13551_),
    .COUT(_13552_),
    .SUM(_13553_));
 sky130_fd_sc_hd__ha_1 _27994_ (.A(_12451_),
    .B(_12461_),
    .COUT(_13555_),
    .SUM(_13556_));
 sky130_fd_sc_hd__ha_1 _27995_ (.A(_13557_),
    .B(_13558_),
    .COUT(_13559_),
    .SUM(_13560_));
 sky130_fd_sc_hd__ha_2 _27996_ (.A(_12460_),
    .B(_12470_),
    .COUT(_13562_),
    .SUM(_13563_));
 sky130_fd_sc_hd__ha_1 _27997_ (.A(_13564_),
    .B(_13565_),
    .COUT(_13566_),
    .SUM(_13567_));
 sky130_fd_sc_hd__ha_1 _27998_ (.A(_12469_),
    .B(_12479_),
    .COUT(_13569_),
    .SUM(_13570_));
 sky130_fd_sc_hd__ha_1 _27999_ (.A(_13571_),
    .B(_13572_),
    .COUT(_13573_),
    .SUM(_13574_));
 sky130_fd_sc_hd__ha_2 _28000_ (.A(_12478_),
    .B(_12488_),
    .COUT(_13576_),
    .SUM(_13577_));
 sky130_fd_sc_hd__ha_1 _28001_ (.A(_13578_),
    .B(_13579_),
    .COUT(_13580_),
    .SUM(_13581_));
 sky130_fd_sc_hd__ha_1 _28002_ (.A(_12487_),
    .B(_12497_),
    .COUT(_13583_),
    .SUM(_13584_));
 sky130_fd_sc_hd__ha_1 _28003_ (.A(_13585_),
    .B(_13586_),
    .COUT(_13587_),
    .SUM(_13588_));
 sky130_fd_sc_hd__ha_1 _28004_ (.A(_12496_),
    .B(_12506_),
    .COUT(_13590_),
    .SUM(_13591_));
 sky130_fd_sc_hd__ha_1 _28005_ (.A(_13592_),
    .B(_13593_),
    .COUT(_13594_),
    .SUM(_13595_));
 sky130_fd_sc_hd__ha_2 _28006_ (.A(_12505_),
    .B(_12515_),
    .COUT(_13597_),
    .SUM(_13598_));
 sky130_fd_sc_hd__ha_1 _28007_ (.A(_13599_),
    .B(_13600_),
    .COUT(_13601_),
    .SUM(_13602_));
 sky130_fd_sc_hd__ha_2 _28008_ (.A(_12514_),
    .B(_12524_),
    .COUT(_13604_),
    .SUM(_13605_));
 sky130_fd_sc_hd__ha_1 _28009_ (.A(_13606_),
    .B(_13607_),
    .COUT(_13608_),
    .SUM(_13609_));
 sky130_fd_sc_hd__ha_1 _28010_ (.A(_12523_),
    .B(_12533_),
    .COUT(_13611_),
    .SUM(_13612_));
 sky130_fd_sc_hd__ha_4 _28011_ (.A(\hash.CA2.p5[0] ),
    .B(_13400_),
    .COUT(_12534_),
    .SUM(_13613_));
 sky130_fd_sc_hd__ha_1 _28012_ (.A(\hash.CA2.p5[1] ),
    .B(_12258_),
    .COUT(_13614_),
    .SUM(_13615_));
 sky130_fd_sc_hd__ha_2 _28013_ (.A(\hash.CA2.p5[2] ),
    .B(_13414_),
    .COUT(_13616_),
    .SUM(_13617_));
 sky130_fd_sc_hd__ha_2 _28014_ (.A(\hash.CA2.p5[3] ),
    .B(_13421_),
    .COUT(_13618_),
    .SUM(_13619_));
 sky130_fd_sc_hd__ha_2 _28015_ (.A(\hash.CA2.p5[4] ),
    .B(_13428_),
    .COUT(_13620_),
    .SUM(_13621_));
 sky130_fd_sc_hd__ha_2 _28016_ (.A(\hash.CA2.p5[5] ),
    .B(_13435_),
    .COUT(_13622_),
    .SUM(_13623_));
 sky130_fd_sc_hd__ha_1 _28017_ (.A(\hash.CA2.p5[6] ),
    .B(_13442_),
    .COUT(_13624_),
    .SUM(_13625_));
 sky130_fd_sc_hd__ha_1 _28018_ (.A(\hash.CA2.p5[7] ),
    .B(_13449_),
    .COUT(_13626_),
    .SUM(_13627_));
 sky130_fd_sc_hd__ha_1 _28019_ (.A(\hash.CA2.p5[8] ),
    .B(_13456_),
    .COUT(_13628_),
    .SUM(_13629_));
 sky130_fd_sc_hd__ha_2 _28020_ (.A(\hash.CA2.p5[9] ),
    .B(_13463_),
    .COUT(_13630_),
    .SUM(_13631_));
 sky130_fd_sc_hd__ha_2 _28021_ (.A(\hash.CA2.p5[10] ),
    .B(_13470_),
    .COUT(_13632_),
    .SUM(_13633_));
 sky130_fd_sc_hd__ha_2 _28022_ (.A(\hash.CA2.p5[11] ),
    .B(_13477_),
    .COUT(_13634_),
    .SUM(_13635_));
 sky130_fd_sc_hd__ha_1 _28023_ (.A(\hash.CA2.p5[12] ),
    .B(_13484_),
    .COUT(_13636_),
    .SUM(_13637_));
 sky130_fd_sc_hd__ha_2 _28024_ (.A(\hash.CA2.p5[13] ),
    .B(_13491_),
    .COUT(_13638_),
    .SUM(_13639_));
 sky130_fd_sc_hd__ha_2 _28025_ (.A(\hash.CA2.p5[14] ),
    .B(_13498_),
    .COUT(_13640_),
    .SUM(_13641_));
 sky130_fd_sc_hd__ha_2 _28026_ (.A(\hash.CA2.p5[15] ),
    .B(_13505_),
    .COUT(_13642_),
    .SUM(_13643_));
 sky130_fd_sc_hd__ha_1 _28027_ (.A(\hash.CA2.p5[16] ),
    .B(_13512_),
    .COUT(_13644_),
    .SUM(_13645_));
 sky130_fd_sc_hd__ha_1 _28028_ (.A(\hash.CA2.p5[17] ),
    .B(_13519_),
    .COUT(_13646_),
    .SUM(_13647_));
 sky130_fd_sc_hd__ha_1 _28029_ (.A(\hash.CA2.p5[16] ),
    .B(_13512_),
    .COUT(_13648_),
    .SUM(_13649_));
 sky130_fd_sc_hd__ha_2 _28030_ (.A(\hash.CA2.p5[18] ),
    .B(_13526_),
    .COUT(_13650_),
    .SUM(_13651_));
 sky130_fd_sc_hd__ha_1 _28031_ (.A(\hash.CA2.p5[19] ),
    .B(_13533_),
    .COUT(_13652_),
    .SUM(_13653_));
 sky130_fd_sc_hd__ha_4 _28032_ (.A(_13540_),
    .B(\hash.CA2.p5[20] ),
    .COUT(_13654_),
    .SUM(_13655_));
 sky130_fd_sc_hd__ha_1 _28033_ (.A(\hash.CA2.p5[21] ),
    .B(_13547_),
    .COUT(_13656_),
    .SUM(_13657_));
 sky130_fd_sc_hd__ha_4 _28034_ (.A(\hash.CA2.p5[20] ),
    .B(_13540_),
    .COUT(_13658_),
    .SUM(_13659_));
 sky130_fd_sc_hd__ha_1 _28035_ (.A(_13554_),
    .B(\hash.CA2.p5[22] ),
    .COUT(_13660_),
    .SUM(_13661_));
 sky130_fd_sc_hd__ha_4 _28036_ (.A(\hash.CA2.p5[21] ),
    .B(_13547_),
    .COUT(_13662_),
    .SUM(_13663_));
 sky130_fd_sc_hd__ha_1 _28037_ (.A(\hash.CA2.p5[23] ),
    .B(_13561_),
    .COUT(_13664_),
    .SUM(_13665_));
 sky130_fd_sc_hd__ha_1 _28038_ (.A(\hash.CA2.p5[22] ),
    .B(_13554_),
    .COUT(_13666_),
    .SUM(_13667_));
 sky130_fd_sc_hd__ha_1 _28039_ (.A(\hash.CA2.p5[24] ),
    .B(_13568_),
    .COUT(_13668_),
    .SUM(_13669_));
 sky130_fd_sc_hd__ha_1 _28040_ (.A(\hash.CA2.p5[23] ),
    .B(_13561_),
    .COUT(_13670_),
    .SUM(_13671_));
 sky130_fd_sc_hd__ha_1 _28041_ (.A(\hash.CA2.p5[25] ),
    .B(_13575_),
    .COUT(_13672_),
    .SUM(_13673_));
 sky130_fd_sc_hd__ha_2 _28042_ (.A(\hash.CA2.p5[26] ),
    .B(_13582_),
    .COUT(_13674_),
    .SUM(_13675_));
 sky130_fd_sc_hd__ha_1 _28043_ (.A(\hash.CA2.p5[25] ),
    .B(_13575_),
    .COUT(_13676_),
    .SUM(_13677_));
 sky130_fd_sc_hd__ha_2 _28044_ (.A(\hash.CA2.p5[27] ),
    .B(_13589_),
    .COUT(_13678_),
    .SUM(_13679_));
 sky130_fd_sc_hd__ha_1 _28045_ (.A(\hash.CA2.p5[26] ),
    .B(_13582_),
    .COUT(_13680_),
    .SUM(_13681_));
 sky130_fd_sc_hd__ha_2 _28046_ (.A(\hash.CA2.p5[28] ),
    .B(_13596_),
    .COUT(_13682_),
    .SUM(_13683_));
 sky130_fd_sc_hd__ha_1 _28047_ (.A(\hash.CA2.p5[29] ),
    .B(_13603_),
    .COUT(_13684_),
    .SUM(_13685_));
 sky130_fd_sc_hd__ha_1 _28048_ (.A(\hash.CA2.p5[30] ),
    .B(_13610_),
    .COUT(_13686_),
    .SUM(_13687_));
 sky130_fd_sc_hd__ha_1 _28049_ (.A(net590),
    .B(\count7_1[2] ),
    .COUT(_13688_),
    .SUM(_00644_));
 sky130_fd_sc_hd__ha_1 _28050_ (.A(net701),
    .B(\count15_1[2] ),
    .COUT(_13689_),
    .SUM(_00645_));
 sky130_fd_sc_hd__ha_1 _28051_ (.A(\count16_1[1] ),
    .B(\count16_1[2] ),
    .COUT(_13690_),
    .SUM(_00646_));
 sky130_fd_sc_hd__ha_1 _28052_ (.A(\count2_2[1] ),
    .B(\count2_2[2] ),
    .COUT(_13691_),
    .SUM(_00647_));
 sky130_fd_sc_hd__ha_1 _28053_ (.A(net572),
    .B(\count7_2[2] ),
    .COUT(_13692_),
    .SUM(_00648_));
 sky130_fd_sc_hd__ha_1 _28054_ (.A(\count15_2[1] ),
    .B(\count15_2[2] ),
    .COUT(_13693_),
    .SUM(_00649_));
 sky130_fd_sc_hd__ha_1 _28055_ (.A(net642),
    .B(net641),
    .COUT(_13694_),
    .SUM(_00650_));
 sky130_fd_sc_hd__ha_4 _28056_ (.A(_00651_),
    .B(_13695_),
    .COUT(_13696_),
    .SUM(_00652_));
 sky130_fd_sc_hd__ha_4 _28057_ (.A(_00651_),
    .B(\count_1[2] ),
    .COUT(_13697_),
    .SUM(_13698_));
 sky130_fd_sc_hd__ha_4 _28058_ (.A(\count_1[1] ),
    .B(_13695_),
    .COUT(_13699_),
    .SUM(_13700_));
 sky130_fd_sc_hd__ha_4 _28059_ (.A(\count_1[1] ),
    .B(\count_1[2] ),
    .COUT(_13701_),
    .SUM(_13702_));
 sky130_fd_sc_hd__ha_4 _28060_ (.A(_00653_),
    .B(_13703_),
    .COUT(_13704_),
    .SUM(_00654_));
 sky130_fd_sc_hd__ha_4 _28061_ (.A(_00653_),
    .B(\count_2[2] ),
    .COUT(_13705_),
    .SUM(_13706_));
 sky130_fd_sc_hd__ha_4 _28062_ (.A(\count_2[1] ),
    .B(_13703_),
    .COUT(_13707_),
    .SUM(_13708_));
 sky130_fd_sc_hd__ha_4 _28063_ (.A(\count_2[1] ),
    .B(\count_2[2] ),
    .COUT(_13709_),
    .SUM(_13710_));
 sky130_fd_sc_hd__ha_1 _28064_ (.A(_00658_),
    .B(_13711_),
    .COUT(_13712_),
    .SUM(_13713_));
 sky130_fd_sc_hd__ha_1 _28065_ (.A(\count2_1[1] ),
    .B(\count2_1[2] ),
    .COUT(_13714_),
    .SUM(_00643_));
 sky130_fd_sc_hd__ha_1 _28066_ (.A(_13715_),
    .B(_13716_),
    .COUT(_13717_),
    .SUM(_13718_));
 sky130_fd_sc_hd__ha_1 _28067_ (.A(_13719_),
    .B(_13720_),
    .COUT(_13721_),
    .SUM(_13722_));
 sky130_fd_sc_hd__ha_4 _28068_ (.A(_13723_),
    .B(_13724_),
    .COUT(_13725_),
    .SUM(_13726_));
 sky130_fd_sc_hd__ha_1 _28069_ (.A(_13727_),
    .B(_13728_),
    .COUT(_13729_),
    .SUM(_13730_));
 sky130_fd_sc_hd__ha_4 _28070_ (.A(_13732_),
    .B(_13731_),
    .COUT(_13733_),
    .SUM(_13734_));
 sky130_fd_sc_hd__ha_1 _28071_ (.A(_13735_),
    .B(_13736_),
    .COUT(_13737_),
    .SUM(_13738_));
 sky130_fd_sc_hd__ha_1 _28072_ (.A(_13739_),
    .B(_13740_),
    .COUT(_13741_),
    .SUM(_13742_));
 sky130_fd_sc_hd__ha_1 _28073_ (.A(_13743_),
    .B(_13744_),
    .COUT(_13745_),
    .SUM(_13746_));
 sky130_fd_sc_hd__ha_2 _28074_ (.A(_13747_),
    .B(_13748_),
    .COUT(_13749_),
    .SUM(_13750_));
 sky130_fd_sc_hd__ha_2 _28075_ (.A(_13751_),
    .B(_13752_),
    .COUT(_13753_),
    .SUM(_13754_));
 sky130_fd_sc_hd__ha_2 _28076_ (.A(_13755_),
    .B(_13756_),
    .COUT(_13757_),
    .SUM(_13758_));
 sky130_fd_sc_hd__ha_1 _28077_ (.A(_13759_),
    .B(_13760_),
    .COUT(_13761_),
    .SUM(_13762_));
 sky130_fd_sc_hd__ha_1 _28078_ (.A(_13763_),
    .B(_13764_),
    .COUT(_13765_),
    .SUM(_13766_));
 sky130_fd_sc_hd__ha_4 _28079_ (.A(_13768_),
    .B(_13767_),
    .COUT(_13769_),
    .SUM(_13770_));
 sky130_fd_sc_hd__ha_1 _28080_ (.A(_13771_),
    .B(_13772_),
    .COUT(_13773_),
    .SUM(_13774_));
 sky130_fd_sc_hd__ha_1 _28081_ (.A(_13775_),
    .B(_13776_),
    .COUT(_13777_),
    .SUM(_13778_));
 sky130_fd_sc_hd__ha_1 _28082_ (.A(_13779_),
    .B(_13780_),
    .COUT(_13781_),
    .SUM(_13782_));
 sky130_fd_sc_hd__ha_1 _28083_ (.A(_13783_),
    .B(_13784_),
    .COUT(_13785_),
    .SUM(_13786_));
 sky130_fd_sc_hd__ha_2 _28084_ (.A(_13787_),
    .B(_13788_),
    .COUT(_13789_),
    .SUM(_13790_));
 sky130_fd_sc_hd__ha_1 _28085_ (.A(_13791_),
    .B(_13792_),
    .COUT(_13793_),
    .SUM(_13794_));
 sky130_fd_sc_hd__ha_1 _28086_ (.A(_13795_),
    .B(_13796_),
    .COUT(_13797_),
    .SUM(_13798_));
 sky130_fd_sc_hd__ha_1 _28087_ (.A(_13799_),
    .B(_13800_),
    .COUT(_13801_),
    .SUM(_13802_));
 sky130_fd_sc_hd__ha_1 _28088_ (.A(_13803_),
    .B(_13804_),
    .COUT(_13805_),
    .SUM(_13806_));
 sky130_fd_sc_hd__ha_1 _28089_ (.A(_13807_),
    .B(_13808_),
    .COUT(_13809_),
    .SUM(_13810_));
 sky130_fd_sc_hd__ha_1 _28090_ (.A(_13811_),
    .B(_13812_),
    .COUT(_13813_),
    .SUM(_13814_));
 sky130_fd_sc_hd__ha_1 _28091_ (.A(_13815_),
    .B(_13816_),
    .COUT(_13817_),
    .SUM(_13818_));
 sky130_fd_sc_hd__ha_1 _28092_ (.A(_13819_),
    .B(_13820_),
    .COUT(_13821_),
    .SUM(_13822_));
 sky130_fd_sc_hd__ha_1 _28093_ (.A(_13823_),
    .B(_13824_),
    .COUT(_13825_),
    .SUM(_13826_));
 sky130_fd_sc_hd__ha_1 _28094_ (.A(_13827_),
    .B(_13828_),
    .COUT(_13829_),
    .SUM(_13830_));
 sky130_fd_sc_hd__ha_1 _28095_ (.A(_13831_),
    .B(_13832_),
    .COUT(_13833_),
    .SUM(_13834_));
 sky130_fd_sc_hd__ha_2 _28096_ (.A(_13835_),
    .B(_13836_),
    .COUT(_12549_),
    .SUM(\hash.CA1.p4[1] ));
 sky130_fd_sc_hd__ha_1 _28097_ (.A(_13067_),
    .B(\hash.CA1.p4[1] ),
    .COUT(_13837_),
    .SUM(_13838_));
 sky130_fd_sc_hd__ha_1 _28098_ (.A(_12550_),
    .B(_12548_),
    .COUT(_13839_),
    .SUM(_13840_));
 sky130_fd_sc_hd__ha_1 _28099_ (.A(\hash.CA1.p4[2] ),
    .B(_13841_),
    .COUT(_13842_),
    .SUM(_13843_));
 sky130_fd_sc_hd__ha_2 _28100_ (.A(_12547_),
    .B(_13844_),
    .COUT(_13845_),
    .SUM(_13846_));
 sky130_fd_sc_hd__ha_1 _28101_ (.A(\hash.CA1.p4[3] ),
    .B(_13847_),
    .COUT(_13848_),
    .SUM(_13849_));
 sky130_fd_sc_hd__ha_2 _28102_ (.A(_13850_),
    .B(_12559_),
    .COUT(_13851_),
    .SUM(_13852_));
 sky130_fd_sc_hd__ha_1 _28103_ (.A(\hash.CA1.p4[4] ),
    .B(_13853_),
    .COUT(_13854_),
    .SUM(_13855_));
 sky130_fd_sc_hd__ha_2 _28104_ (.A(_12558_),
    .B(_13856_),
    .COUT(_13857_),
    .SUM(_13858_));
 sky130_fd_sc_hd__ha_1 _28105_ (.A(\hash.CA1.p4[5] ),
    .B(_13859_),
    .COUT(_13860_),
    .SUM(_13861_));
 sky130_fd_sc_hd__ha_2 _28106_ (.A(_13862_),
    .B(_12567_),
    .COUT(_13863_),
    .SUM(_13864_));
 sky130_fd_sc_hd__ha_1 _28107_ (.A(\hash.CA1.p4[6] ),
    .B(_13865_),
    .COUT(_13866_),
    .SUM(_13867_));
 sky130_fd_sc_hd__ha_1 _28108_ (.A(_12566_),
    .B(_13868_),
    .COUT(_13869_),
    .SUM(_13870_));
 sky130_fd_sc_hd__ha_1 _28109_ (.A(\hash.CA1.p4[7] ),
    .B(_13871_),
    .COUT(_13872_),
    .SUM(_13873_));
 sky130_fd_sc_hd__ha_1 _28110_ (.A(_13874_),
    .B(_13875_),
    .COUT(_13876_),
    .SUM(_13877_));
 sky130_fd_sc_hd__ha_1 _28111_ (.A(\hash.CA1.p4[8] ),
    .B(_13878_),
    .COUT(_13879_),
    .SUM(_13880_));
 sky130_fd_sc_hd__ha_2 _28112_ (.A(_13881_),
    .B(_12580_),
    .COUT(_13882_),
    .SUM(_13883_));
 sky130_fd_sc_hd__ha_1 _28113_ (.A(\hash.CA1.p4[9] ),
    .B(_13884_),
    .COUT(_13885_),
    .SUM(_13886_));
 sky130_fd_sc_hd__ha_2 _28114_ (.A(_12579_),
    .B(_12583_),
    .COUT(_13887_),
    .SUM(_13888_));
 sky130_fd_sc_hd__ha_1 _28115_ (.A(\hash.CA1.p4[10] ),
    .B(_13889_),
    .COUT(_13890_),
    .SUM(_13891_));
 sky130_fd_sc_hd__ha_2 _28116_ (.A(_12582_),
    .B(_13892_),
    .COUT(_13893_),
    .SUM(_13894_));
 sky130_fd_sc_hd__ha_1 _28117_ (.A(\hash.CA1.p4[11] ),
    .B(_13895_),
    .COUT(_13896_),
    .SUM(_13897_));
 sky130_fd_sc_hd__ha_1 _28118_ (.A(_13898_),
    .B(_13899_),
    .COUT(_13900_),
    .SUM(_13901_));
 sky130_fd_sc_hd__ha_1 _28119_ (.A(\hash.CA1.p4[12] ),
    .B(_13902_),
    .COUT(_13903_),
    .SUM(_13904_));
 sky130_fd_sc_hd__ha_2 _28120_ (.A(_13905_),
    .B(_12596_),
    .COUT(_13906_),
    .SUM(_13907_));
 sky130_fd_sc_hd__ha_1 _28121_ (.A(\hash.CA1.p4[13] ),
    .B(_13908_),
    .COUT(_13909_),
    .SUM(_13910_));
 sky130_fd_sc_hd__ha_2 _28122_ (.A(_12595_),
    .B(_13911_),
    .COUT(_13912_),
    .SUM(_13913_));
 sky130_fd_sc_hd__ha_1 _28123_ (.A(\hash.CA1.p4[14] ),
    .B(_13914_),
    .COUT(_13915_),
    .SUM(_13916_));
 sky130_fd_sc_hd__ha_2 _28124_ (.A(_13917_),
    .B(_13918_),
    .COUT(_13919_),
    .SUM(_13920_));
 sky130_fd_sc_hd__ha_1 _28125_ (.A(\hash.CA1.p4[15] ),
    .B(_13921_),
    .COUT(_13922_),
    .SUM(_13923_));
 sky130_fd_sc_hd__ha_2 _28126_ (.A(_13924_),
    .B(_13925_),
    .COUT(_13926_),
    .SUM(_13927_));
 sky130_fd_sc_hd__ha_1 _28127_ (.A(\hash.CA1.p4[16] ),
    .B(_13928_),
    .COUT(_13929_),
    .SUM(_13930_));
 sky130_fd_sc_hd__ha_2 _28128_ (.A(_13931_),
    .B(_13932_),
    .COUT(_13933_),
    .SUM(_13934_));
 sky130_fd_sc_hd__ha_1 _28129_ (.A(\hash.CA1.p4[17] ),
    .B(_13935_),
    .COUT(_13936_),
    .SUM(_13937_));
 sky130_fd_sc_hd__ha_2 _28130_ (.A(_13938_),
    .B(_12619_),
    .COUT(_13939_),
    .SUM(_13940_));
 sky130_fd_sc_hd__ha_2 _28131_ (.A(\hash.CA1.p4[18] ),
    .B(_13941_),
    .COUT(_13942_),
    .SUM(_13943_));
 sky130_fd_sc_hd__ha_2 _28132_ (.A(_12618_),
    .B(_12622_),
    .COUT(_13944_),
    .SUM(_13945_));
 sky130_fd_sc_hd__ha_2 _28133_ (.A(\hash.CA1.p4[19] ),
    .B(_13946_),
    .COUT(_13947_),
    .SUM(_13948_));
 sky130_fd_sc_hd__ha_2 _28134_ (.A(_12621_),
    .B(_12625_),
    .COUT(_13949_),
    .SUM(_13950_));
 sky130_fd_sc_hd__ha_2 _28135_ (.A(\hash.CA1.p4[20] ),
    .B(_13951_),
    .COUT(_13952_),
    .SUM(_13953_));
 sky130_fd_sc_hd__ha_2 _28136_ (.A(_12624_),
    .B(_12628_),
    .COUT(_13954_),
    .SUM(_13955_));
 sky130_fd_sc_hd__ha_1 _28137_ (.A(\hash.CA1.p4[21] ),
    .B(_13956_),
    .COUT(_13957_),
    .SUM(_13958_));
 sky130_fd_sc_hd__ha_2 _28138_ (.A(_12627_),
    .B(_12631_),
    .COUT(_13959_),
    .SUM(_13960_));
 sky130_fd_sc_hd__ha_1 _28139_ (.A(\hash.CA1.p4[22] ),
    .B(_13961_),
    .COUT(_13962_),
    .SUM(_13963_));
 sky130_fd_sc_hd__ha_2 _28140_ (.A(_12630_),
    .B(_13964_),
    .COUT(_13965_),
    .SUM(_13966_));
 sky130_fd_sc_hd__ha_2 _28141_ (.A(\hash.CA1.p4[23] ),
    .B(_13967_),
    .COUT(_13968_),
    .SUM(_13969_));
 sky130_fd_sc_hd__ha_2 _28142_ (.A(_13970_),
    .B(_13971_),
    .COUT(_13972_),
    .SUM(_13973_));
 sky130_fd_sc_hd__ha_2 _28143_ (.A(\hash.CA1.p4[24] ),
    .B(_13974_),
    .COUT(_13975_),
    .SUM(_13976_));
 sky130_fd_sc_hd__ha_2 _28144_ (.A(_13977_),
    .B(_13978_),
    .COUT(_13979_),
    .SUM(_13980_));
 sky130_fd_sc_hd__ha_2 _28145_ (.A(\hash.CA1.p4[25] ),
    .B(_13981_),
    .COUT(_13982_),
    .SUM(_13983_));
 sky130_fd_sc_hd__ha_2 _28146_ (.A(_13984_),
    .B(_13985_),
    .COUT(_13986_),
    .SUM(_13987_));
 sky130_fd_sc_hd__ha_1 _28147_ (.A(\hash.CA1.p4[26] ),
    .B(_06480_),
    .COUT(_13989_),
    .SUM(_13990_));
 sky130_fd_sc_hd__ha_2 _28148_ (.A(_13991_),
    .B(_13992_),
    .COUT(_13993_),
    .SUM(_13994_));
 sky130_fd_sc_hd__ha_1 _28149_ (.A(\hash.CA1.p4[27] ),
    .B(_13995_),
    .COUT(_13996_),
    .SUM(_13997_));
 sky130_fd_sc_hd__ha_2 _28150_ (.A(_13998_),
    .B(_13999_),
    .COUT(_14000_),
    .SUM(_14001_));
 sky130_fd_sc_hd__ha_1 _28151_ (.A(\hash.CA1.p4[28] ),
    .B(_14002_),
    .COUT(_14003_),
    .SUM(_14004_));
 sky130_fd_sc_hd__ha_2 _28152_ (.A(_14005_),
    .B(_12664_),
    .COUT(_14006_),
    .SUM(_14007_));
 sky130_fd_sc_hd__ha_1 _28153_ (.A(\hash.CA1.p4[29] ),
    .B(_14008_),
    .COUT(_14009_),
    .SUM(_14010_));
 sky130_fd_sc_hd__ha_2 _28154_ (.A(_12663_),
    .B(_12667_),
    .COUT(_14011_),
    .SUM(_14012_));
 sky130_fd_sc_hd__ha_1 _28155_ (.A(\hash.CA1.p4[30] ),
    .B(_14013_),
    .COUT(_14014_),
    .SUM(_14015_));
 sky130_fd_sc_hd__ha_1 _28156_ (.A(_12824_),
    .B(_12676_),
    .COUT(_14016_),
    .SUM(_11749_));
 sky130_fd_sc_hd__ha_1 _28157_ (.A(_00843_),
    .B(_12539_),
    .COUT(_14017_),
    .SUM(_14018_));
 sky130_fd_sc_hd__ha_1 _28158_ (.A(_00813_),
    .B(_14019_),
    .COUT(_14020_),
    .SUM(_14021_));
 sky130_fd_sc_hd__ha_1 _28159_ (.A(_14022_),
    .B(_00781_),
    .COUT(_14023_),
    .SUM(_14024_));
 sky130_fd_sc_hd__ha_1 _28160_ (.A(_12828_),
    .B(_14025_),
    .COUT(_14026_),
    .SUM(_11748_));
 sky130_fd_sc_hd__ha_1 _28161_ (.A(_13067_),
    .B(_13841_),
    .COUT(_14027_),
    .SUM(_11747_));
 sky130_fd_sc_hd__ha_1 _28162_ (.A(\hash.CA1.b[1] ),
    .B(\hash.CA1.b[0] ),
    .COUT(_14028_),
    .SUM(_11746_));
 sky130_fd_sc_hd__ha_1 _28163_ (.A(\hash.CA1.k_i1[0] ),
    .B(\hash.CA1.w_i1[0] ),
    .COUT(_12668_),
    .SUM(_12825_));
 sky130_fd_sc_hd__ha_4 _28164_ (.A(_14030_),
    .B(_14029_),
    .COUT(_14031_),
    .SUM(_13056_));
 sky130_fd_sc_hd__ha_1 _28165_ (.A(\hash.CA1.k_i1[1] ),
    .B(\hash.CA1.w_i1[1] ),
    .COUT(_14032_),
    .SUM(_14033_));
 sky130_fd_sc_hd__ha_1 _28166_ (.A(_14034_),
    .B(_14035_),
    .COUT(_14036_),
    .SUM(_14037_));
 sky130_fd_sc_hd__ha_1 _28167_ (.A(\hash.CA1.k_i1[2] ),
    .B(\hash.CA1.w_i1[2] ),
    .COUT(_14038_),
    .SUM(_14039_));
 sky130_fd_sc_hd__ha_4 _28168_ (.A(_14040_),
    .B(_14041_),
    .COUT(_14042_),
    .SUM(_14043_));
 sky130_fd_sc_hd__ha_1 _28169_ (.A(_12677_),
    .B(_12683_),
    .COUT(_14044_),
    .SUM(_14045_));
 sky130_fd_sc_hd__ha_2 _28170_ (.A(\hash.CA1.k_i1[3] ),
    .B(\hash.CA1.w_i1[3] ),
    .COUT(_14046_),
    .SUM(_14047_));
 sky130_fd_sc_hd__ha_1 _28171_ (.A(_14048_),
    .B(_14049_),
    .COUT(_14050_),
    .SUM(_14051_));
 sky130_fd_sc_hd__ha_1 _28172_ (.A(_12682_),
    .B(_14052_),
    .COUT(_14053_),
    .SUM(_14054_));
 sky130_fd_sc_hd__ha_1 _28173_ (.A(\hash.CA1.k_i1[4] ),
    .B(\hash.CA1.w_i1[4] ),
    .COUT(_14055_),
    .SUM(_14056_));
 sky130_fd_sc_hd__ha_4 _28174_ (.A(_14057_),
    .B(_14058_),
    .COUT(_14059_),
    .SUM(_14060_));
 sky130_fd_sc_hd__ha_1 _28175_ (.A(_14061_),
    .B(_14062_),
    .COUT(_14063_),
    .SUM(_14064_));
 sky130_fd_sc_hd__ha_2 _28176_ (.A(\hash.CA1.k_i1[5] ),
    .B(\hash.CA1.w_i1[5] ),
    .COUT(_14065_),
    .SUM(_14066_));
 sky130_fd_sc_hd__ha_4 _28177_ (.A(_14067_),
    .B(_14068_),
    .COUT(_14069_),
    .SUM(_14070_));
 sky130_fd_sc_hd__ha_2 _28178_ (.A(_14071_),
    .B(_12698_),
    .COUT(_14072_),
    .SUM(_14073_));
 sky130_fd_sc_hd__ha_2 _28179_ (.A(\hash.CA1.k_i1[6] ),
    .B(\hash.CA1.w_i1[6] ),
    .COUT(_14074_),
    .SUM(_14075_));
 sky130_fd_sc_hd__ha_4 _28180_ (.A(_14076_),
    .B(_14077_),
    .COUT(_14078_),
    .SUM(_14079_));
 sky130_fd_sc_hd__ha_2 _28181_ (.A(_12697_),
    .B(_12703_),
    .COUT(_14080_),
    .SUM(_14081_));
 sky130_fd_sc_hd__ha_2 _28182_ (.A(\hash.CA1.k_i1[7] ),
    .B(\hash.CA1.w_i1[7] ),
    .COUT(_14082_),
    .SUM(_14083_));
 sky130_fd_sc_hd__ha_1 _28183_ (.A(_14084_),
    .B(_14085_),
    .COUT(_14086_),
    .SUM(_14087_));
 sky130_fd_sc_hd__ha_2 _28184_ (.A(_12702_),
    .B(_12708_),
    .COUT(_14088_),
    .SUM(_14089_));
 sky130_fd_sc_hd__ha_2 _28185_ (.A(\hash.CA1.k_i1[8] ),
    .B(\hash.CA1.w_i1[8] ),
    .COUT(_14090_),
    .SUM(_14091_));
 sky130_fd_sc_hd__ha_1 _28186_ (.A(_14092_),
    .B(_14093_),
    .COUT(_14094_),
    .SUM(_14095_));
 sky130_fd_sc_hd__ha_2 _28187_ (.A(_12707_),
    .B(_14096_),
    .COUT(_14097_),
    .SUM(_14098_));
 sky130_fd_sc_hd__ha_2 _28188_ (.A(\hash.CA1.k_i1[9] ),
    .B(\hash.CA1.w_i1[9] ),
    .COUT(_14099_),
    .SUM(_14100_));
 sky130_fd_sc_hd__ha_1 _28189_ (.A(_14101_),
    .B(_14102_),
    .COUT(_14103_),
    .SUM(_14104_));
 sky130_fd_sc_hd__ha_2 _28190_ (.A(_14105_),
    .B(_12718_),
    .COUT(_14106_),
    .SUM(_14107_));
 sky130_fd_sc_hd__ha_2 _28191_ (.A(\hash.CA1.k_i1[10] ),
    .B(\hash.CA1.w_i1[10] ),
    .COUT(_14108_),
    .SUM(_14109_));
 sky130_fd_sc_hd__ha_2 _28192_ (.A(_14110_),
    .B(_14111_),
    .COUT(_14112_),
    .SUM(_14113_));
 sky130_fd_sc_hd__ha_4 _28193_ (.A(_12717_),
    .B(_14114_),
    .COUT(_14115_),
    .SUM(_14116_));
 sky130_fd_sc_hd__ha_2 _28194_ (.A(\hash.CA1.k_i1[11] ),
    .B(\hash.CA1.w_i1[11] ),
    .COUT(_14117_),
    .SUM(_14118_));
 sky130_fd_sc_hd__ha_2 _28195_ (.A(_14119_),
    .B(_14120_),
    .COUT(_14121_),
    .SUM(_14122_));
 sky130_fd_sc_hd__ha_2 _28196_ (.A(_14123_),
    .B(_14124_),
    .COUT(_14125_),
    .SUM(_14126_));
 sky130_fd_sc_hd__ha_2 _28197_ (.A(\hash.CA1.k_i1[12] ),
    .B(\hash.CA1.w_i1[12] ),
    .COUT(_14127_),
    .SUM(_14128_));
 sky130_fd_sc_hd__ha_1 _28198_ (.A(_14129_),
    .B(_14130_),
    .COUT(_14131_),
    .SUM(_14132_));
 sky130_fd_sc_hd__ha_1 _28199_ (.A(_14133_),
    .B(_12733_),
    .COUT(_14134_),
    .SUM(_14135_));
 sky130_fd_sc_hd__ha_2 _28200_ (.A(\hash.CA1.k_i1[13] ),
    .B(\hash.CA1.w_i1[13] ),
    .COUT(_14136_),
    .SUM(_14137_));
 sky130_fd_sc_hd__ha_2 _28201_ (.A(_14138_),
    .B(_14139_),
    .COUT(_14140_),
    .SUM(_14141_));
 sky130_fd_sc_hd__ha_1 _28202_ (.A(_12732_),
    .B(_12738_),
    .COUT(_14142_),
    .SUM(_14143_));
 sky130_fd_sc_hd__ha_2 _28203_ (.A(\hash.CA1.k_i1[14] ),
    .B(\hash.CA1.w_i1[14] ),
    .COUT(_14144_),
    .SUM(_14145_));
 sky130_fd_sc_hd__ha_1 _28204_ (.A(_14146_),
    .B(_14147_),
    .COUT(_14148_),
    .SUM(_14149_));
 sky130_fd_sc_hd__ha_4 _28205_ (.A(_12737_),
    .B(_14150_),
    .COUT(_14151_),
    .SUM(_14152_));
 sky130_fd_sc_hd__ha_2 _28206_ (.A(\hash.CA1.k_i1[15] ),
    .B(\hash.CA1.w_i1[15] ),
    .COUT(_14153_),
    .SUM(_14154_));
 sky130_fd_sc_hd__ha_1 _28207_ (.A(_14155_),
    .B(_14156_),
    .COUT(_14157_),
    .SUM(_14158_));
 sky130_fd_sc_hd__ha_2 _28208_ (.A(_14159_),
    .B(_14160_),
    .COUT(_14161_),
    .SUM(_14162_));
 sky130_fd_sc_hd__ha_2 _28209_ (.A(\hash.CA1.k_i1[16] ),
    .B(\hash.CA1.w_i1[16] ),
    .COUT(_14163_),
    .SUM(_14164_));
 sky130_fd_sc_hd__ha_2 _28210_ (.A(_14165_),
    .B(_14166_),
    .COUT(_14167_),
    .SUM(_14168_));
 sky130_fd_sc_hd__ha_2 _28211_ (.A(_14169_),
    .B(_12753_),
    .COUT(_14170_),
    .SUM(_14171_));
 sky130_fd_sc_hd__ha_2 _28212_ (.A(\hash.CA1.k_i1[17] ),
    .B(\hash.CA1.w_i1[17] ),
    .COUT(_14172_),
    .SUM(_14173_));
 sky130_fd_sc_hd__ha_2 _28213_ (.A(_14174_),
    .B(_14175_),
    .COUT(_14176_),
    .SUM(_14177_));
 sky130_fd_sc_hd__ha_4 _28214_ (.A(_12752_),
    .B(_12758_),
    .COUT(_14178_),
    .SUM(_14179_));
 sky130_fd_sc_hd__ha_2 _28215_ (.A(\hash.CA1.k_i1[18] ),
    .B(\hash.CA1.w_i1[18] ),
    .COUT(_14180_),
    .SUM(_14181_));
 sky130_fd_sc_hd__ha_2 _28216_ (.A(_14182_),
    .B(_14183_),
    .COUT(_14184_),
    .SUM(_14185_));
 sky130_fd_sc_hd__ha_4 _28217_ (.A(_12757_),
    .B(_12763_),
    .COUT(_14186_),
    .SUM(_14187_));
 sky130_fd_sc_hd__ha_4 _28218_ (.A(\hash.CA1.k_i1[19] ),
    .B(\hash.CA1.w_i1[19] ),
    .COUT(_14188_),
    .SUM(_14189_));
 sky130_fd_sc_hd__ha_2 _28219_ (.A(_14190_),
    .B(_14191_),
    .COUT(_14192_),
    .SUM(_14193_));
 sky130_fd_sc_hd__ha_4 _28220_ (.A(_12762_),
    .B(_12768_),
    .COUT(_14194_),
    .SUM(_14195_));
 sky130_fd_sc_hd__ha_2 _28221_ (.A(\hash.CA1.k_i1[20] ),
    .B(\hash.CA1.w_i1[20] ),
    .COUT(_14196_),
    .SUM(_14197_));
 sky130_fd_sc_hd__ha_2 _28222_ (.A(_14198_),
    .B(_14199_),
    .COUT(_14200_),
    .SUM(_14201_));
 sky130_fd_sc_hd__ha_1 _28223_ (.A(_12767_),
    .B(_12773_),
    .COUT(_14202_),
    .SUM(_14203_));
 sky130_fd_sc_hd__ha_2 _28224_ (.A(\hash.CA1.k_i1[21] ),
    .B(\hash.CA1.w_i1[21] ),
    .COUT(_14204_),
    .SUM(_14205_));
 sky130_fd_sc_hd__ha_1 _28225_ (.A(_14206_),
    .B(_14207_),
    .COUT(_14208_),
    .SUM(_14209_));
 sky130_fd_sc_hd__ha_4 _28226_ (.A(_14210_),
    .B(_12772_),
    .COUT(_14211_),
    .SUM(_14212_));
 sky130_fd_sc_hd__ha_2 _28227_ (.A(\hash.CA1.k_i1[22] ),
    .B(\hash.CA1.w_i1[22] ),
    .COUT(_14213_),
    .SUM(_14214_));
 sky130_fd_sc_hd__ha_1 _28228_ (.A(_14215_),
    .B(_14216_),
    .COUT(_14217_),
    .SUM(_14218_));
 sky130_fd_sc_hd__ha_1 _28229_ (.A(_14219_),
    .B(_14220_),
    .COUT(_14221_),
    .SUM(_14222_));
 sky130_fd_sc_hd__ha_2 _28230_ (.A(\hash.CA1.k_i1[23] ),
    .B(\hash.CA1.w_i1[23] ),
    .COUT(_14223_),
    .SUM(_14224_));
 sky130_fd_sc_hd__ha_1 _28231_ (.A(_14225_),
    .B(_14226_),
    .COUT(_14227_),
    .SUM(_14228_));
 sky130_fd_sc_hd__ha_4 _28232_ (.A(_14230_),
    .B(_14229_),
    .COUT(_14231_),
    .SUM(_14232_));
 sky130_fd_sc_hd__ha_2 _28233_ (.A(\hash.CA1.k_i1[24] ),
    .B(\hash.CA1.w_i1[24] ),
    .COUT(_14233_),
    .SUM(_14234_));
 sky130_fd_sc_hd__ha_1 _28234_ (.A(_14235_),
    .B(_14236_),
    .COUT(_14237_),
    .SUM(_14238_));
 sky130_fd_sc_hd__ha_1 _28235_ (.A(_14239_),
    .B(_14240_),
    .COUT(_14241_),
    .SUM(_14242_));
 sky130_fd_sc_hd__ha_2 _28236_ (.A(\hash.CA1.k_i1[25] ),
    .B(\hash.CA1.w_i1[25] ),
    .COUT(_14243_),
    .SUM(_14244_));
 sky130_fd_sc_hd__ha_1 _28237_ (.A(_14245_),
    .B(_14246_),
    .COUT(_14247_),
    .SUM(_14248_));
 sky130_fd_sc_hd__ha_1 _28238_ (.A(_14249_),
    .B(_14250_),
    .COUT(_14251_),
    .SUM(_14252_));
 sky130_fd_sc_hd__ha_1 _28239_ (.A(\hash.CA1.k_i1[26] ),
    .B(\hash.CA1.w_i1[26] ),
    .COUT(_14253_),
    .SUM(_14254_));
 sky130_fd_sc_hd__ha_2 _28240_ (.A(_14255_),
    .B(_14256_),
    .COUT(_14257_),
    .SUM(_14258_));
 sky130_fd_sc_hd__ha_1 _28241_ (.A(_14259_),
    .B(_12803_),
    .COUT(_14260_),
    .SUM(_14261_));
 sky130_fd_sc_hd__ha_2 _28242_ (.A(\hash.CA1.k_i1[27] ),
    .B(\hash.CA1.w_i1[27] ),
    .COUT(_14262_),
    .SUM(_14263_));
 sky130_fd_sc_hd__ha_1 _28243_ (.A(_14264_),
    .B(_14265_),
    .COUT(_14266_),
    .SUM(_14267_));
 sky130_fd_sc_hd__ha_1 _28244_ (.A(_12802_),
    .B(_14268_),
    .COUT(_14269_),
    .SUM(_14270_));
 sky130_fd_sc_hd__ha_4 _28245_ (.A(\hash.CA1.k_i1[28] ),
    .B(\hash.CA1.w_i1[28] ),
    .COUT(_14271_),
    .SUM(_14272_));
 sky130_fd_sc_hd__ha_2 _28246_ (.A(_14273_),
    .B(_14274_),
    .COUT(_14275_),
    .SUM(_14276_));
 sky130_fd_sc_hd__ha_1 _28247_ (.A(_14277_),
    .B(_14278_),
    .COUT(_14279_),
    .SUM(_14280_));
 sky130_fd_sc_hd__ha_2 _28248_ (.A(\hash.CA1.k_i1[29] ),
    .B(\hash.CA1.w_i1[29] ),
    .COUT(_14281_),
    .SUM(_14282_));
 sky130_fd_sc_hd__ha_1 _28249_ (.A(_14283_),
    .B(_14284_),
    .COUT(_14285_),
    .SUM(_14286_));
 sky130_fd_sc_hd__ha_1 _28250_ (.A(_14287_),
    .B(_12818_),
    .COUT(_14288_),
    .SUM(_14289_));
 sky130_fd_sc_hd__ha_4 _28251_ (.A(\hash.CA1.k_i1[30] ),
    .B(\hash.CA1.w_i1[30] ),
    .COUT(_14290_),
    .SUM(_14291_));
 sky130_fd_sc_hd__ha_1 _28252_ (.A(_14292_),
    .B(_14293_),
    .COUT(_14294_),
    .SUM(_14295_));
 sky130_fd_sc_hd__ha_1 _28253_ (.A(_12817_),
    .B(_14296_),
    .COUT(_14297_),
    .SUM(_14298_));
 sky130_fd_sc_hd__ha_1 _28254_ (.A(_14299_),
    .B(_14300_),
    .COUT(_14301_),
    .SUM(_14302_));
 sky130_fd_sc_hd__ha_1 _28255_ (.A(_14303_),
    .B(_14304_),
    .COUT(_14305_),
    .SUM(_14306_));
 sky130_fd_sc_hd__ha_1 _28256_ (.A(_14307_),
    .B(_14308_),
    .COUT(_14309_),
    .SUM(_14310_));
 sky130_fd_sc_hd__ha_1 _28257_ (.A(_14311_),
    .B(_14312_),
    .COUT(_14313_),
    .SUM(_14314_));
 sky130_fd_sc_hd__ha_1 _28258_ (.A(_14315_),
    .B(_14316_),
    .COUT(_14317_),
    .SUM(_14318_));
 sky130_fd_sc_hd__ha_1 _28259_ (.A(_14319_),
    .B(_14320_),
    .COUT(_14321_),
    .SUM(_14322_));
 sky130_fd_sc_hd__ha_1 _28260_ (.A(_14323_),
    .B(_14324_),
    .COUT(_14325_),
    .SUM(_14326_));
 sky130_fd_sc_hd__ha_1 _28261_ (.A(_14327_),
    .B(_12893_),
    .COUT(_14328_),
    .SUM(_14329_));
 sky130_fd_sc_hd__ha_4 _28262_ (.A(_12901_),
    .B(_12892_),
    .COUT(_14330_),
    .SUM(_14331_));
 sky130_fd_sc_hd__ha_1 _28263_ (.A(_12900_),
    .B(_12910_),
    .COUT(_14332_),
    .SUM(_14333_));
 sky130_fd_sc_hd__ha_4 _28264_ (.A(_12909_),
    .B(_12916_),
    .COUT(_14334_),
    .SUM(_14335_));
 sky130_fd_sc_hd__ha_1 _28265_ (.A(_12915_),
    .B(_12922_),
    .COUT(_14336_),
    .SUM(_14337_));
 sky130_fd_sc_hd__ha_1 _28266_ (.A(_12921_),
    .B(_12929_),
    .COUT(_14338_),
    .SUM(_14339_));
 sky130_fd_sc_hd__ha_1 _28267_ (.A(_12928_),
    .B(_12937_),
    .COUT(_14340_),
    .SUM(_14341_));
 sky130_fd_sc_hd__ha_4 _28268_ (.A(_12936_),
    .B(_12944_),
    .COUT(_14342_),
    .SUM(_14343_));
 sky130_fd_sc_hd__ha_4 _28269_ (.A(_12943_),
    .B(_12950_),
    .COUT(_14344_),
    .SUM(_14345_));
 sky130_fd_sc_hd__ha_4 _28270_ (.A(_12949_),
    .B(_12956_),
    .COUT(_14346_),
    .SUM(_14347_));
 sky130_fd_sc_hd__ha_4 _28271_ (.A(_12955_),
    .B(_12962_),
    .COUT(_14348_),
    .SUM(_14349_));
 sky130_fd_sc_hd__ha_1 _28272_ (.A(_12961_),
    .B(_12971_),
    .COUT(_14350_),
    .SUM(_14351_));
 sky130_fd_sc_hd__ha_1 _28273_ (.A(_12970_),
    .B(_12980_),
    .COUT(_14352_),
    .SUM(_14353_));
 sky130_fd_sc_hd__ha_1 _28274_ (.A(_12979_),
    .B(_12987_),
    .COUT(_14354_),
    .SUM(_14355_));
 sky130_fd_sc_hd__ha_2 _28275_ (.A(_12986_),
    .B(_12996_),
    .COUT(_14356_),
    .SUM(_14357_));
 sky130_fd_sc_hd__ha_1 _28276_ (.A(_12995_),
    .B(_13003_),
    .COUT(_14358_),
    .SUM(_14359_));
 sky130_fd_sc_hd__ha_2 _28277_ (.A(_13002_),
    .B(_13012_),
    .COUT(_14360_),
    .SUM(_14361_));
 sky130_fd_sc_hd__ha_2 _28278_ (.A(_13011_),
    .B(_13018_),
    .COUT(_14362_),
    .SUM(_14363_));
 sky130_fd_sc_hd__ha_2 _28279_ (.A(_13017_),
    .B(_13026_),
    .COUT(_14364_),
    .SUM(_14365_));
 sky130_fd_sc_hd__ha_1 _28280_ (.A(_13025_),
    .B(_13034_),
    .COUT(_14366_),
    .SUM(_14367_));
 sky130_fd_sc_hd__ha_1 _28281_ (.A(_13033_),
    .B(_13040_),
    .COUT(_14368_),
    .SUM(_14369_));
 sky130_fd_sc_hd__ha_1 _28282_ (.A(_13039_),
    .B(_14370_),
    .COUT(_14371_),
    .SUM(_14372_));
 sky130_fd_sc_hd__ha_1 _28283_ (.A(_14373_),
    .B(_14374_),
    .COUT(_14375_),
    .SUM(\hash.CA1.p1[0] ));
 sky130_fd_sc_hd__ha_1 _28284_ (.A(_12827_),
    .B(_13056_),
    .COUT(_14376_),
    .SUM(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__ha_1 _28285_ (.A(_14376_),
    .B(_14377_),
    .COUT(_14378_),
    .SUM(\hash.CA1.p2[1] ));
 sky130_fd_sc_hd__ha_1 _28286_ (.A(_13057_),
    .B(_12678_),
    .COUT(_14379_),
    .SUM(\hash.CA1.p3[1] ));
 sky130_fd_sc_hd__ha_1 _28287_ (.A(\hash.CA1.c[0] ),
    .B(\hash.CA1.p4[0] ),
    .COUT(_13066_),
    .SUM(\hash.CA1.p5[0] ));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[1]$_SDFF_PP0_  (.D(_00907_),
    .Q(\count15_1[1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[2]$_SDFF_PP0_  (.D(_00908_),
    .Q(\count15_1[2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[3]$_SDFF_PP0_  (.D(_00909_),
    .Q(\count15_1[3] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[4]$_SDFF_PP0_  (.D(_00910_),
    .Q(\count15_1[4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[5]$_SDFF_PP0_  (.D(_00911_),
    .Q(\count15_1[5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[1]$_SDFF_PP1_  (.D(_00912_),
    .Q(\count15_2[1] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[2]$_SDFF_PP0_  (.D(_00913_),
    .Q(\count15_2[2] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[3]$_SDFF_PP0_  (.D(_00914_),
    .Q(\count15_2[3] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[4]$_SDFF_PP0_  (.D(_00915_),
    .Q(\count15_2[4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[5]$_SDFF_PP0_  (.D(_00916_),
    .Q(\count15_2[5] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[1]$_SDFF_PP0_  (.D(_00917_),
    .Q(\count16_1[1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[2]$_SDFF_PP0_  (.D(_00918_),
    .Q(\count16_1[2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[3]$_SDFF_PP0_  (.D(_00919_),
    .Q(\count16_1[3] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[4]$_SDFF_PP0_  (.D(_00920_),
    .Q(\count16_1[4] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_1[5]$_SDFF_PP0_  (.D(_00921_),
    .Q(\count16_1[5] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[1]$_SDFF_PP0_  (.D(_00922_),
    .Q(\count16_2[1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[2]$_SDFF_PP0_  (.D(_00923_),
    .Q(\count16_2[2] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[3]$_SDFF_PP0_  (.D(_00924_),
    .Q(\count16_2[3] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[4]$_SDFF_PP0_  (.D(_00925_),
    .Q(\count16_2[4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_4 \count16_2[5]$_SDFF_PP0_  (.D(_00926_),
    .Q(\count16_2[5] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[1]$_SDFF_PP1_  (.D(_00927_),
    .Q(\count2_1[1] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[2]$_SDFF_PP1_  (.D(_00928_),
    .Q(\count2_1[2] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[3]$_SDFF_PP1_  (.D(_00929_),
    .Q(\count2_1[3] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[4]$_SDFF_PP0_  (.D(_00930_),
    .Q(\count2_1[4] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[5]$_SDFF_PP0_  (.D(_00931_),
    .Q(\count2_1[5] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[1]$_SDFF_PP1_  (.D(_00932_),
    .Q(\count2_2[1] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[2]$_SDFF_PP1_  (.D(_00933_),
    .Q(\count2_2[2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[3]$_SDFF_PP1_  (.D(_00934_),
    .Q(\count2_2[3] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[4]$_SDFF_PP0_  (.D(_00935_),
    .Q(\count2_2[4] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 \count2_2[5]$_SDFF_PP0_  (.D(_00936_),
    .Q(\count2_2[5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[1]$_SDFF_PP0_  (.D(_00937_),
    .Q(\count7_1[1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[2]$_SDFF_PP0_  (.D(_00938_),
    .Q(\count7_1[2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[3]$_SDFF_PP1_  (.D(_00939_),
    .Q(\count7_1[3] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[4]$_SDFF_PP0_  (.D(_00940_),
    .Q(\count7_1[4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_1[5]$_SDFF_PP0_  (.D(_00941_),
    .Q(\count7_1[5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[1]$_SDFF_PP1_  (.D(_00942_),
    .Q(\count7_2[1] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[2]$_SDFF_PP0_  (.D(_00943_),
    .Q(\count7_2[2] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[3]$_SDFF_PP1_  (.D(_00944_),
    .Q(\count7_2[3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[4]$_SDFF_PP0_  (.D(_00945_),
    .Q(\count7_2[4] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_4 \count7_2[5]$_SDFF_PP0_  (.D(_00946_),
    .Q(\count7_2[5] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 \count_1[1]$_SDFFE_PP0N_  (.D(_00947_),
    .Q(\count_1[1] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 \count_1[2]$_SDFFE_PP0N_  (.D(_00948_),
    .Q(\count_1[2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_1[3]$_SDFFE_PP0N_  (.D(_00949_),
    .Q(\count_1[3] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_1[4]$_SDFFE_PP1N_  (.D(_00950_),
    .Q(\count_1[4] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_1[5]$_SDFFE_PP0N_  (.D(_00951_),
    .Q(\count_1[5] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 \count_2[1]$_SDFFE_PP0N_  (.D(_00952_),
    .Q(\count_2[1] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 \count_2[2]$_SDFFE_PP0N_  (.D(_00953_),
    .Q(\count_2[2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_2[3]$_SDFFE_PP0N_  (.D(_00954_),
    .Q(\count_2[3] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_2[4]$_SDFFE_PP1N_  (.D(_00955_),
    .Q(\count_2[4] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_2[5]$_SDFFE_PP0N_  (.D(_00956_),
    .Q(\count_2[5] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[6]$_SDFFE_PP0N_  (.D(_00957_),
    .Q(\count_2[6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash1[1]$_SDFFE_PP0N_  (.D(_00958_),
    .Q(\count_hash1[1] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash1[2]$_SDFFE_PP0N_  (.D(_00959_),
    .Q(\count_hash1[2] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash1[3]$_SDFFE_PP0N_  (.D(_00960_),
    .Q(\count_hash1[3] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash1[4]$_SDFFE_PP0N_  (.D(_00961_),
    .Q(\count_hash1[4] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash1[5]$_SDFFE_PP0N_  (.D(_00962_),
    .Q(\count_hash1[5] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 \count_hash1[6]$_SDFFE_PP0N_  (.D(_00963_),
    .Q(\count_hash1[6] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash2[1]$_SDFFE_PP0N_  (.D(_00964_),
    .Q(\count_hash2[1] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash2[2]$_SDFFE_PP0N_  (.D(_00965_),
    .Q(\count_hash2[2] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash2[3]$_SDFFE_PP0N_  (.D(_00966_),
    .Q(\count_hash2[3] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_4 \count_hash2[4]$_SDFFE_PP0N_  (.D(_00967_),
    .Q(\count_hash2[4] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 \count_hash2[5]$_SDFFE_PP0N_  (.D(_00968_),
    .Q(\count_hash2[5] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \done$_DFFE_PN_  (.D(_00128_),
    .DE(_09893_),
    .Q(done),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[0]$_DFF_P_  (.D(\hash.CA1.S0.X[0] ),
    .Q(\hash.CA2.a_dash[0] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[10]$_DFF_P_  (.D(\hash.CA1.S0.X[10] ),
    .Q(\hash.CA2.a_dash[10] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[11]$_DFF_P_  (.D(\hash.CA1.S0.X[11] ),
    .Q(\hash.CA2.a_dash[11] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[12]$_DFF_P_  (.D(\hash.CA1.S0.X[12] ),
    .Q(\hash.CA2.a_dash[12] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[13]$_DFF_P_  (.D(\hash.CA1.S0.X[13] ),
    .Q(\hash.CA2.a_dash[13] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[14]$_DFF_P_  (.D(\hash.CA1.S0.X[14] ),
    .Q(\hash.CA2.a_dash[14] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[15]$_DFF_P_  (.D(\hash.CA1.S0.X[15] ),
    .Q(\hash.CA2.a_dash[15] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[16]$_DFF_P_  (.D(\hash.CA1.S0.X[16] ),
    .Q(\hash.CA2.a_dash[16] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[17]$_DFF_P_  (.D(\hash.CA1.S0.X[17] ),
    .Q(\hash.CA2.a_dash[17] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[18]$_DFF_P_  (.D(_06312_),
    .Q(\hash.CA2.a_dash[18] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[19]$_DFF_P_  (.D(\hash.CA1.S0.X[19] ),
    .Q(\hash.CA2.a_dash[19] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[1]$_DFF_P_  (.D(\hash.CA1.S0.X[1] ),
    .Q(\hash.CA2.a_dash[1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[20]$_DFF_P_  (.D(\hash.CA1.S0.X[20] ),
    .Q(\hash.CA2.a_dash[20] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[21]$_DFF_P_  (.D(_06338_),
    .Q(\hash.CA2.a_dash[21] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[22]$_DFF_P_  (.D(\hash.CA1.S0.X[22] ),
    .Q(\hash.CA2.a_dash[22] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[23]$_DFF_P_  (.D(\hash.CA1.S0.X[23] ),
    .Q(\hash.CA2.a_dash[23] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[24]$_DFF_P_  (.D(\hash.CA1.S0.X[24] ),
    .Q(\hash.CA2.a_dash[24] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[25]$_DFF_P_  (.D(\hash.CA1.S0.X[25] ),
    .Q(\hash.CA2.a_dash[25] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[26]$_DFF_P_  (.D(\hash.CA1.S0.X[26] ),
    .Q(\hash.CA2.a_dash[26] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[27]$_DFF_P_  (.D(\hash.CA1.S0.X[27] ),
    .Q(\hash.CA2.a_dash[27] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[28]$_DFF_P_  (.D(\hash.CA1.S0.X[28] ),
    .Q(\hash.CA2.a_dash[28] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[29]$_DFF_P_  (.D(\hash.CA1.S0.X[29] ),
    .Q(\hash.CA2.a_dash[29] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[2]$_DFF_P_  (.D(\hash.CA1.S0.X[2] ),
    .Q(\hash.CA2.a_dash[2] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[30]$_DFF_P_  (.D(\hash.CA1.S0.X[30] ),
    .Q(\hash.CA2.a_dash[30] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[31]$_DFF_P_  (.D(\hash.CA1.S0.X[31] ),
    .Q(\hash.CA2.a_dash[31] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[3]$_DFF_P_  (.D(\hash.CA1.S0.X[3] ),
    .Q(\hash.CA2.a_dash[3] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[4]$_DFF_P_  (.D(\hash.CA1.S0.X[4] ),
    .Q(\hash.CA2.a_dash[4] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[5]$_DFF_P_  (.D(\hash.CA1.S0.X[5] ),
    .Q(\hash.CA2.a_dash[5] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[6]$_DFF_P_  (.D(\hash.CA1.S0.X[6] ),
    .Q(\hash.CA2.a_dash[6] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[7]$_DFF_P_  (.D(\hash.CA1.S0.X[7] ),
    .Q(\hash.CA2.a_dash[7] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[8]$_DFF_P_  (.D(\hash.CA1.S0.X[8] ),
    .Q(\hash.CA2.a_dash[8] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.a_cap[9]$_DFF_P_  (.D(\hash.CA1.S0.X[9] ),
    .Q(\hash.CA2.a_dash[9] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[0]$_DFF_P_  (.D(\hash.CA1.b[0] ),
    .Q(\hash.CA2.b_dash[0] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[10]$_DFF_P_  (.D(\hash.CA1.b[10] ),
    .Q(\hash.CA2.b_dash[10] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[11]$_DFF_P_  (.D(\hash.CA1.b[11] ),
    .Q(\hash.CA2.b_dash[11] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[12]$_DFF_P_  (.D(\hash.CA1.b[12] ),
    .Q(\hash.CA2.b_dash[12] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[13]$_DFF_P_  (.D(\hash.CA1.b[13] ),
    .Q(\hash.CA2.b_dash[13] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[14]$_DFF_P_  (.D(\hash.CA1.b[14] ),
    .Q(\hash.CA2.b_dash[14] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[15]$_DFF_P_  (.D(\hash.CA1.b[15] ),
    .Q(\hash.CA2.b_dash[15] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[16]$_DFF_P_  (.D(\hash.CA1.b[16] ),
    .Q(\hash.CA2.b_dash[16] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[17]$_DFF_P_  (.D(\hash.CA1.b[17] ),
    .Q(\hash.CA2.b_dash[17] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[18]$_DFF_P_  (.D(\hash.CA1.b[18] ),
    .Q(\hash.CA2.b_dash[18] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[19]$_DFF_P_  (.D(\hash.CA1.b[19] ),
    .Q(\hash.CA2.b_dash[19] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[1]$_DFF_P_  (.D(\hash.CA1.b[1] ),
    .Q(\hash.CA2.b_dash[1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[20]$_DFF_P_  (.D(\hash.CA1.b[20] ),
    .Q(\hash.CA2.b_dash[20] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[21]$_DFF_P_  (.D(_06478_),
    .Q(\hash.CA2.b_dash[21] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[22]$_DFF_P_  (.D(\hash.CA1.b[22] ),
    .Q(\hash.CA2.b_dash[22] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[23]$_DFF_P_  (.D(_06479_),
    .Q(\hash.CA2.b_dash[23] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[24]$_DFF_P_  (.D(\hash.CA1.b[24] ),
    .Q(\hash.CA2.b_dash[24] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[25]$_DFF_P_  (.D(\hash.CA1.b[25] ),
    .Q(\hash.CA2.b_dash[25] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[26]$_DFF_P_  (.D(\hash.CA1.b[26] ),
    .Q(\hash.CA2.b_dash[26] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[27]$_DFF_P_  (.D(_06481_),
    .Q(\hash.CA2.b_dash[27] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[28]$_DFF_P_  (.D(\hash.CA1.b[28] ),
    .Q(\hash.CA2.b_dash[28] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[29]$_DFF_P_  (.D(\hash.CA1.b[29] ),
    .Q(\hash.CA2.b_dash[29] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[2]$_DFF_P_  (.D(\hash.CA1.b[2] ),
    .Q(\hash.CA2.b_dash[2] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[30]$_DFF_P_  (.D(\hash.CA1.b[30] ),
    .Q(\hash.CA2.b_dash[30] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[31]$_DFF_P_  (.D(\hash.CA1.b[31] ),
    .Q(\hash.CA2.b_dash[31] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[3]$_DFF_P_  (.D(\hash.CA1.b[3] ),
    .Q(\hash.CA2.b_dash[3] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[4]$_DFF_P_  (.D(\hash.CA1.b[4] ),
    .Q(\hash.CA2.b_dash[4] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[5]$_DFF_P_  (.D(\hash.CA1.b[5] ),
    .Q(\hash.CA2.b_dash[5] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[6]$_DFF_P_  (.D(\hash.CA1.b[6] ),
    .Q(\hash.CA2.b_dash[6] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.b_cap[7]$_DFF_P_  (.D(\hash.CA1.b[7] ),
    .Q(\hash.CA2.b_dash[7] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[8]$_DFF_P_  (.D(\hash.CA1.b[8] ),
    .Q(\hash.CA2.b_dash[8] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[9]$_DFF_P_  (.D(\hash.CA1.b[9] ),
    .Q(\hash.CA2.b_dash[9] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[0]$_DFF_P_  (.D(\hash.CA1.S1.X[0] ),
    .Q(\hash.CA2.e_dash[0] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[10]$_DFF_P_  (.D(\hash.CA1.S1.X[10] ),
    .Q(\hash.CA2.e_dash[10] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[11]$_DFF_P_  (.D(\hash.CA1.S1.X[11] ),
    .Q(\hash.CA2.e_dash[11] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[12]$_DFF_P_  (.D(\hash.CA1.S1.X[12] ),
    .Q(\hash.CA2.e_dash[12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[13]$_DFF_P_  (.D(\hash.CA1.S1.X[13] ),
    .Q(\hash.CA2.e_dash[13] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[14]$_DFF_P_  (.D(\hash.CA1.S1.X[14] ),
    .Q(\hash.CA2.e_dash[14] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[15]$_DFF_P_  (.D(\hash.CA1.S1.X[15] ),
    .Q(\hash.CA2.e_dash[15] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[16]$_DFF_P_  (.D(_06804_),
    .Q(\hash.CA2.e_dash[16] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[17]$_DFF_P_  (.D(\hash.CA1.S1.X[17] ),
    .Q(\hash.CA2.e_dash[17] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[18]$_DFF_P_  (.D(\hash.CA1.S1.X[18] ),
    .Q(\hash.CA2.e_dash[18] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[19]$_DFF_P_  (.D(\hash.CA1.S1.X[19] ),
    .Q(\hash.CA2.e_dash[19] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[1]$_DFF_P_  (.D(\hash.CA1.S1.X[1] ),
    .Q(\hash.CA2.e_dash[1] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[20]$_DFF_P_  (.D(\hash.CA1.S1.X[20] ),
    .Q(\hash.CA2.e_dash[20] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[21]$_DFF_P_  (.D(\hash.CA1.S1.X[21] ),
    .Q(\hash.CA2.e_dash[21] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[22]$_DFF_P_  (.D(_06854_),
    .Q(\hash.CA2.e_dash[22] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[23]$_DFF_P_  (.D(\hash.CA1.S1.X[23] ),
    .Q(\hash.CA2.e_dash[23] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[24]$_DFF_P_  (.D(\hash.CA1.S1.X[24] ),
    .Q(\hash.CA2.e_dash[24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[25]$_DFF_P_  (.D(net1020),
    .Q(\hash.CA2.e_dash[25] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[26]$_DFF_P_  (.D(\hash.CA1.S1.X[26] ),
    .Q(\hash.CA2.e_dash[26] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[27]$_DFF_P_  (.D(\hash.CA1.S1.X[27] ),
    .Q(\hash.CA2.e_dash[27] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[28]$_DFF_P_  (.D(\hash.CA1.S1.X[28] ),
    .Q(\hash.CA2.e_dash[28] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[29]$_DFF_P_  (.D(\hash.CA1.S1.X[29] ),
    .Q(\hash.CA2.e_dash[29] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[2]$_DFF_P_  (.D(\hash.CA1.S1.X[2] ),
    .Q(\hash.CA2.e_dash[2] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[30]$_DFF_P_  (.D(\hash.CA1.S1.X[30] ),
    .Q(\hash.CA2.e_dash[30] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[31]$_DFF_P_  (.D(_06922_),
    .Q(\hash.CA2.e_dash[31] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[3]$_DFF_P_  (.D(\hash.CA1.S1.X[3] ),
    .Q(\hash.CA2.e_dash[3] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[4]$_DFF_P_  (.D(\hash.CA1.S1.X[4] ),
    .Q(\hash.CA2.e_dash[4] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[5]$_DFF_P_  (.D(\hash.CA1.S1.X[5] ),
    .Q(\hash.CA2.e_dash[5] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[6]$_DFF_P_  (.D(\hash.CA1.S1.X[6] ),
    .Q(\hash.CA2.e_dash[6] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[7]$_DFF_P_  (.D(\hash.CA1.S1.X[7] ),
    .Q(\hash.CA2.e_dash[7] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[8]$_DFF_P_  (.D(\hash.CA1.S1.X[8] ),
    .Q(\hash.CA2.e_dash[8] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[9]$_DFF_P_  (.D(\hash.CA1.S1.X[9] ),
    .Q(\hash.CA2.e_dash[9] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[0]$_DFF_P_  (.D(\hash.CA1.f[0] ),
    .Q(\hash.CA2.f_dash[0] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[10]$_DFF_P_  (.D(\hash.CA1.f[10] ),
    .Q(\hash.CA2.f_dash[10] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[11]$_DFF_P_  (.D(\hash.CA1.f[11] ),
    .Q(\hash.CA2.f_dash[11] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[12]$_DFF_P_  (.D(\hash.CA1.f[12] ),
    .Q(\hash.CA2.f_dash[12] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.f_cap[13]$_DFF_P_  (.D(\hash.CA1.f[13] ),
    .Q(\hash.CA2.f_dash[13] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.f_cap[14]$_DFF_P_  (.D(\hash.CA1.f[14] ),
    .Q(\hash.CA2.f_dash[14] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.f_cap[15]$_DFF_P_  (.D(\hash.CA1.f[15] ),
    .Q(\hash.CA2.f_dash[15] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[16]$_DFF_P_  (.D(\hash.CA1.f[16] ),
    .Q(\hash.CA2.f_dash[16] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[17]$_DFF_P_  (.D(\hash.CA1.f[17] ),
    .Q(\hash.CA2.f_dash[17] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[18]$_DFF_P_  (.D(\hash.CA1.f[18] ),
    .Q(\hash.CA2.f_dash[18] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[19]$_DFF_P_  (.D(\hash.CA1.f[19] ),
    .Q(\hash.CA2.f_dash[19] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[1]$_DFF_P_  (.D(\hash.CA1.f[1] ),
    .Q(\hash.CA2.f_dash[1] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[20]$_DFF_P_  (.D(\hash.CA1.f[20] ),
    .Q(\hash.CA2.f_dash[20] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[21]$_DFF_P_  (.D(\hash.CA1.f[21] ),
    .Q(\hash.CA2.f_dash[21] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[22]$_DFF_P_  (.D(\hash.CA1.f[22] ),
    .Q(\hash.CA2.f_dash[22] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[23]$_DFF_P_  (.D(\hash.CA1.f[23] ),
    .Q(\hash.CA2.f_dash[23] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[24]$_DFF_P_  (.D(_06668_),
    .Q(\hash.CA2.f_dash[24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[25]$_DFF_P_  (.D(\hash.CA1.f[25] ),
    .Q(\hash.CA2.f_dash[25] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[26]$_DFF_P_  (.D(\hash.CA1.f[26] ),
    .Q(\hash.CA2.f_dash[26] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[27]$_DFF_P_  (.D(\hash.CA1.f[27] ),
    .Q(\hash.CA2.f_dash[27] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[28]$_DFF_P_  (.D(\hash.CA1.f[28] ),
    .Q(\hash.CA2.f_dash[28] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[29]$_DFF_P_  (.D(\hash.CA1.f[29] ),
    .Q(\hash.CA2.f_dash[29] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[2]$_DFF_P_  (.D(\hash.CA1.f[2] ),
    .Q(\hash.CA2.f_dash[2] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[30]$_DFF_P_  (.D(\hash.CA1.f[30] ),
    .Q(\hash.CA2.f_dash[30] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.f_cap[31]$_DFF_P_  (.D(\hash.CA1.f[31] ),
    .Q(\hash.CA2.f_dash[31] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.f_cap[3]$_DFF_P_  (.D(\hash.CA1.f[3] ),
    .Q(\hash.CA2.f_dash[3] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[4]$_DFF_P_  (.D(\hash.CA1.f[4] ),
    .Q(\hash.CA2.f_dash[4] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[5]$_DFF_P_  (.D(\hash.CA1.f[5] ),
    .Q(\hash.CA2.f_dash[5] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.f_cap[6]$_DFF_P_  (.D(\hash.CA1.f[6] ),
    .Q(\hash.CA2.f_dash[6] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[7]$_DFF_P_  (.D(\hash.CA1.f[7] ),
    .Q(\hash.CA2.f_dash[7] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.f_cap[8]$_DFF_P_  (.D(\hash.CA1.f[8] ),
    .Q(\hash.CA2.f_dash[8] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[9]$_DFF_P_  (.D(\hash.CA1.f[9] ),
    .Q(\hash.CA2.f_dash[9] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[0]$_DFFE_PN_  (.D(_00658_),
    .DE(_00906_),
    .Q(net901),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[10]$_DFFE_PN_  (.D(_00659_),
    .DE(_00906_),
    .Q(net912),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[11]$_DFFE_PN_  (.D(_00660_),
    .DE(_00906_),
    .Q(net913),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[12]$_DFFE_PN_  (.D(_00661_),
    .DE(_00906_),
    .Q(net914),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[13]$_DFFE_PN_  (.D(_00662_),
    .DE(_00906_),
    .Q(net915),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[14]$_DFFE_PN_  (.D(_00663_),
    .DE(_00906_),
    .Q(net916),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[15]$_DFFE_PN_  (.D(_00664_),
    .DE(_00906_),
    .Q(net917),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[16]$_DFFE_PN_  (.D(_00665_),
    .DE(_00906_),
    .Q(net919),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[17]$_DFFE_PN_  (.D(_00666_),
    .DE(_00906_),
    .Q(net920),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[18]$_DFFE_PN_  (.D(_00667_),
    .DE(_00906_),
    .Q(net921),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[19]$_DFFE_PN_  (.D(_00668_),
    .DE(_00906_),
    .Q(net922),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[1]$_DFFE_PN_  (.D(_00669_),
    .DE(_00906_),
    .Q(net902),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[20]$_DFFE_PN_  (.D(_00670_),
    .DE(_00906_),
    .Q(net923),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[21]$_DFFE_PN_  (.D(_00671_),
    .DE(_00906_),
    .Q(net924),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[22]$_DFFE_PN_  (.D(_00672_),
    .DE(_00906_),
    .Q(net925),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[23]$_DFFE_PN_  (.D(_00673_),
    .DE(_00906_),
    .Q(net926),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[24]$_DFFE_PN_  (.D(_00674_),
    .DE(_00906_),
    .Q(net927),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[25]$_DFFE_PN_  (.D(_00675_),
    .DE(_00906_),
    .Q(net928),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[26]$_DFFE_PN_  (.D(_00676_),
    .DE(_00906_),
    .Q(net930),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[27]$_DFFE_PN_  (.D(_00677_),
    .DE(_00906_),
    .Q(net931),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[28]$_DFFE_PN_  (.D(_00678_),
    .DE(_00906_),
    .Q(net932),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[29]$_DFFE_PN_  (.D(_00679_),
    .DE(_00906_),
    .Q(net933),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[2]$_DFFE_PN_  (.D(_00680_),
    .DE(_00906_),
    .Q(net903),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[30]$_DFFE_PN_  (.D(_00681_),
    .DE(_00906_),
    .Q(net934),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[31]$_DFFE_PN_  (.D(_00682_),
    .DE(_00906_),
    .Q(net935),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[3]$_DFFE_PN_  (.D(_00683_),
    .DE(_00906_),
    .Q(net904),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[4]$_DFFE_PN_  (.D(_00684_),
    .DE(_00906_),
    .Q(net905),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[5]$_DFFE_PN_  (.D(_00685_),
    .DE(_00906_),
    .Q(net906),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[6]$_DFFE_PN_  (.D(_00686_),
    .DE(_00906_),
    .Q(net908),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[7]$_DFFE_PN_  (.D(_00687_),
    .DE(_00906_),
    .Q(net909),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[8]$_DFFE_PN_  (.D(_00688_),
    .DE(_00906_),
    .Q(net910),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[9]$_DFFE_PN_  (.D(_00689_),
    .DE(_00906_),
    .Q(net911),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[0]$_DFFE_PN_  (.D(_00690_),
    .DE(_00906_),
    .Q(net865),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[10]$_DFFE_PN_  (.D(_00691_),
    .DE(_00906_),
    .Q(net877),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[11]$_DFFE_PN_  (.D(_00692_),
    .DE(_00906_),
    .Q(net878),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[12]$_DFFE_PN_  (.D(_00693_),
    .DE(_00906_),
    .Q(net879),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[13]$_DFFE_PN_  (.D(_00694_),
    .DE(_00906_),
    .Q(net880),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[14]$_DFFE_PN_  (.D(_00695_),
    .DE(_00906_),
    .Q(net881),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[15]$_DFFE_PN_  (.D(_00696_),
    .DE(_00906_),
    .Q(net882),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[16]$_DFFE_PN_  (.D(_00697_),
    .DE(_00906_),
    .Q(net883),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[17]$_DFFE_PN_  (.D(_00698_),
    .DE(_00906_),
    .Q(net884),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[18]$_DFFE_PN_  (.D(_00699_),
    .DE(_00906_),
    .Q(net886),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[19]$_DFFE_PN_  (.D(_00700_),
    .DE(_00906_),
    .Q(net887),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[1]$_DFFE_PN_  (.D(_11746_),
    .DE(_00906_),
    .Q(net866),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[20]$_DFFE_PN_  (.D(_00701_),
    .DE(_00906_),
    .Q(net888),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[21]$_DFFE_PN_  (.D(_00702_),
    .DE(_00906_),
    .Q(net889),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[22]$_DFFE_PN_  (.D(_00703_),
    .DE(_00906_),
    .Q(net890),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[23]$_DFFE_PN_  (.D(_00704_),
    .DE(_00906_),
    .Q(net891),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[24]$_DFFE_PN_  (.D(_00705_),
    .DE(_00906_),
    .Q(net892),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[25]$_DFFE_PN_  (.D(_00706_),
    .DE(_00906_),
    .Q(net893),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[26]$_DFFE_PN_  (.D(_00707_),
    .DE(_00906_),
    .Q(net894),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[27]$_DFFE_PN_  (.D(_00708_),
    .DE(_00906_),
    .Q(net895),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[28]$_DFFE_PN_  (.D(_00709_),
    .DE(_00906_),
    .Q(net897),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[29]$_DFFE_PN_  (.D(_00710_),
    .DE(_00906_),
    .Q(net898),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[2]$_DFFE_PN_  (.D(_00711_),
    .DE(_00906_),
    .Q(net867),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[30]$_DFFE_PN_  (.D(_00712_),
    .DE(_00906_),
    .Q(net899),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[31]$_DFFE_PN_  (.D(_00713_),
    .DE(_00906_),
    .Q(net900),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[3]$_DFFE_PN_  (.D(_00714_),
    .DE(_00906_),
    .Q(net868),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[4]$_DFFE_PN_  (.D(_00715_),
    .DE(_00906_),
    .Q(net869),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[5]$_DFFE_PN_  (.D(_00716_),
    .DE(_00906_),
    .Q(net870),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[6]$_DFFE_PN_  (.D(_00717_),
    .DE(_00906_),
    .Q(net871),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[7]$_DFFE_PN_  (.D(_00718_),
    .DE(_00906_),
    .Q(net872),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[8]$_DFFE_PN_  (.D(_00719_),
    .DE(_00906_),
    .Q(net875),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[9]$_DFFE_PN_  (.D(_00720_),
    .DE(_00906_),
    .Q(net876),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[0]$_DFFE_PN_  (.D(\hash.CA1.c[0] ),
    .DE(_00906_),
    .Q(net830),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[10]$_DFFE_PN_  (.D(_00750_),
    .DE(_00906_),
    .Q(net841),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[11]$_DFFE_PN_  (.D(_00722_),
    .DE(_00906_),
    .Q(net842),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[12]$_DFFE_PN_  (.D(_00723_),
    .DE(_00906_),
    .Q(net843),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[13]$_DFFE_PN_  (.D(_00724_),
    .DE(_00906_),
    .Q(net844),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[14]$_DFFE_PN_  (.D(_00725_),
    .DE(_00906_),
    .Q(net845),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[15]$_DFFE_PN_  (.D(_00726_),
    .DE(_00906_),
    .Q(net846),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[16]$_DFFE_PN_  (.D(_00727_),
    .DE(_00906_),
    .Q(net847),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[17]$_DFFE_PN_  (.D(_00728_),
    .DE(_00906_),
    .Q(net848),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[18]$_DFFE_PN_  (.D(_00729_),
    .DE(_00906_),
    .Q(net849),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[19]$_DFFE_PN_  (.D(_00730_),
    .DE(_00906_),
    .Q(net850),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[1]$_DFFE_PN_  (.D(_00721_),
    .DE(_00906_),
    .Q(net831),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[20]$_DFFE_PN_  (.D(_00731_),
    .DE(_00906_),
    .Q(net852),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[21]$_DFFE_PN_  (.D(_00732_),
    .DE(_00906_),
    .Q(net853),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[22]$_DFFE_PN_  (.D(_00733_),
    .DE(_00906_),
    .Q(net854),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[23]$_DFFE_PN_  (.D(_00734_),
    .DE(_00906_),
    .Q(net855),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[24]$_DFFE_PN_  (.D(_00735_),
    .DE(_00906_),
    .Q(net856),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[25]$_DFFE_PN_  (.D(_00736_),
    .DE(_00906_),
    .Q(net857),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[26]$_DFFE_PN_  (.D(_00737_),
    .DE(_00906_),
    .Q(net858),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[27]$_DFFE_PN_  (.D(_00738_),
    .DE(_00906_),
    .Q(net859),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[28]$_DFFE_PN_  (.D(_00739_),
    .DE(_00906_),
    .Q(net860),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[29]$_DFFE_PN_  (.D(_00740_),
    .DE(_00906_),
    .Q(net861),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[2]$_DFFE_PN_  (.D(_11747_),
    .DE(_00906_),
    .Q(net832),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[30]$_DFFE_PN_  (.D(_00741_),
    .DE(_00906_),
    .Q(net863),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[31]$_DFFE_PN_  (.D(_00743_),
    .DE(_00906_),
    .Q(net864),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[3]$_DFFE_PN_  (.D(_00742_),
    .DE(_00906_),
    .Q(net833),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[4]$_DFFE_PN_  (.D(_00744_),
    .DE(_00906_),
    .Q(net834),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[5]$_DFFE_PN_  (.D(_00745_),
    .DE(_00906_),
    .Q(net835),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[6]$_DFFE_PN_  (.D(_00746_),
    .DE(_00906_),
    .Q(net836),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[7]$_DFFE_PN_  (.D(_00747_),
    .DE(_00906_),
    .Q(net837),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[8]$_DFFE_PN_  (.D(_00748_),
    .DE(_00906_),
    .Q(net838),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[9]$_DFFE_PN_  (.D(_00749_),
    .DE(_00906_),
    .Q(net839),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[0]$_DFFE_PN_  (.D(\hash.CA1.d[0] ),
    .DE(_00906_),
    .Q(net794),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[10]$_DFFE_PN_  (.D(_00780_),
    .DE(_00906_),
    .Q(net805),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[11]$_DFFE_PN_  (.D(_00752_),
    .DE(_00906_),
    .Q(net806),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[12]$_DFFE_PN_  (.D(_00753_),
    .DE(_00906_),
    .Q(net808),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[13]$_DFFE_PN_  (.D(_00754_),
    .DE(_00906_),
    .Q(net809),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[14]$_DFFE_PN_  (.D(_00755_),
    .DE(_00906_),
    .Q(net810),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[15]$_DFFE_PN_  (.D(_00756_),
    .DE(_00906_),
    .Q(net811),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[16]$_DFFE_PN_  (.D(_00757_),
    .DE(_00906_),
    .Q(net812),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[17]$_DFFE_PN_  (.D(_00758_),
    .DE(_00906_),
    .Q(net813),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[18]$_DFFE_PN_  (.D(_00759_),
    .DE(_00906_),
    .Q(net814),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[19]$_DFFE_PN_  (.D(_00760_),
    .DE(_00906_),
    .Q(net815),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[1]$_DFFE_PN_  (.D(_00751_),
    .DE(_00906_),
    .Q(net795),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[20]$_DFFE_PN_  (.D(_00761_),
    .DE(_00906_),
    .Q(net816),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[21]$_DFFE_PN_  (.D(_00762_),
    .DE(_00906_),
    .Q(net817),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[22]$_DFFE_PN_  (.D(_00763_),
    .DE(_00906_),
    .Q(net819),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[23]$_DFFE_PN_  (.D(_00764_),
    .DE(_00906_),
    .Q(net820),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[24]$_DFFE_PN_  (.D(_00765_),
    .DE(_00906_),
    .Q(net821),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[25]$_DFFE_PN_  (.D(_00766_),
    .DE(_00906_),
    .Q(net822),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[26]$_DFFE_PN_  (.D(_00767_),
    .DE(_00906_),
    .Q(net823),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[27]$_DFFE_PN_  (.D(_00768_),
    .DE(_00906_),
    .Q(net824),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[28]$_DFFE_PN_  (.D(_00769_),
    .DE(_00906_),
    .Q(net825),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[29]$_DFFE_PN_  (.D(_00770_),
    .DE(_00906_),
    .Q(net826),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[2]$_DFFE_PN_  (.D(_11748_),
    .DE(_00906_),
    .Q(net797),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[30]$_DFFE_PN_  (.D(_00771_),
    .DE(_00906_),
    .Q(net827),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[31]$_DFFE_PN_  (.D(_00773_),
    .DE(_00906_),
    .Q(net828),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[3]$_DFFE_PN_  (.D(_00772_),
    .DE(_00906_),
    .Q(net798),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[4]$_DFFE_PN_  (.D(_00774_),
    .DE(_00906_),
    .Q(net799),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[5]$_DFFE_PN_  (.D(_00775_),
    .DE(_00906_),
    .Q(net800),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[6]$_DFFE_PN_  (.D(_00776_),
    .DE(_00906_),
    .Q(net801),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[7]$_DFFE_PN_  (.D(_00777_),
    .DE(_00906_),
    .Q(net802),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[8]$_DFFE_PN_  (.D(_00778_),
    .DE(_00906_),
    .Q(net803),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[9]$_DFFE_PN_  (.D(_00779_),
    .DE(_00906_),
    .Q(net804),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[0]$_DFFE_PN_  (.D(_00781_),
    .DE(_00906_),
    .Q(net1014),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[10]$_DFFE_PN_  (.D(_00782_),
    .DE(_00906_),
    .Q(net770),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[11]$_DFFE_PN_  (.D(_00783_),
    .DE(_00906_),
    .Q(net771),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[12]$_DFFE_PN_  (.D(_00784_),
    .DE(_00906_),
    .Q(net772),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[13]$_DFFE_PN_  (.D(_00785_),
    .DE(_00906_),
    .Q(net773),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[14]$_DFFE_PN_  (.D(_00786_),
    .DE(_00906_),
    .Q(net775),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[15]$_DFFE_PN_  (.D(_00787_),
    .DE(_00906_),
    .Q(net776),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[16]$_DFFE_PN_  (.D(_00788_),
    .DE(_00906_),
    .Q(net777),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[17]$_DFFE_PN_  (.D(_00789_),
    .DE(_00906_),
    .Q(net778),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[18]$_DFFE_PN_  (.D(_00790_),
    .DE(_00906_),
    .Q(net779),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[19]$_DFFE_PN_  (.D(_00791_),
    .DE(_00906_),
    .Q(net780),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[1]$_DFFE_PN_  (.D(_00792_),
    .DE(_00906_),
    .Q(net1015),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[20]$_DFFE_PN_  (.D(_00793_),
    .DE(_00906_),
    .Q(net781),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[21]$_DFFE_PN_  (.D(_00794_),
    .DE(_00906_),
    .Q(net782),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[22]$_DFFE_PN_  (.D(_00795_),
    .DE(_00906_),
    .Q(net783),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[23]$_DFFE_PN_  (.D(_00796_),
    .DE(_00906_),
    .Q(net784),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[24]$_DFFE_PN_  (.D(_00797_),
    .DE(_00906_),
    .Q(net786),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[25]$_DFFE_PN_  (.D(_00798_),
    .DE(_00906_),
    .Q(net787),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[26]$_DFFE_PN_  (.D(_00799_),
    .DE(_00906_),
    .Q(net788),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[27]$_DFFE_PN_  (.D(_00800_),
    .DE(_00906_),
    .Q(net789),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[28]$_DFFE_PN_  (.D(_00801_),
    .DE(_00906_),
    .Q(net790),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[29]$_DFFE_PN_  (.D(_00802_),
    .DE(_00906_),
    .Q(net791),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[2]$_DFFE_PN_  (.D(_00803_),
    .DE(_00906_),
    .Q(net1016),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[30]$_DFFE_PN_  (.D(_00804_),
    .DE(_00906_),
    .Q(net792),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[31]$_DFFE_PN_  (.D(_00805_),
    .DE(_00906_),
    .Q(net793),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[3]$_DFFE_PN_  (.D(_00806_),
    .DE(_00906_),
    .Q(net1017),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[4]$_DFFE_PN_  (.D(_00807_),
    .DE(_00906_),
    .Q(net764),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[5]$_DFFE_PN_  (.D(_00808_),
    .DE(_00906_),
    .Q(net765),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[6]$_DFFE_PN_  (.D(_00809_),
    .DE(_00906_),
    .Q(net766),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[7]$_DFFE_PN_  (.D(_00810_),
    .DE(_00906_),
    .Q(net767),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[8]$_DFFE_PN_  (.D(_00811_),
    .DE(_00906_),
    .Q(net768),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[9]$_DFFE_PN_  (.D(_00812_),
    .DE(_00906_),
    .Q(net769),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[0]$_DFFE_PN_  (.D(\hash.CA1.f[0] ),
    .DE(_00906_),
    .Q(net979),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[10]$_DFFE_PN_  (.D(_00841_),
    .DE(_00906_),
    .Q(net990),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[11]$_DFFE_PN_  (.D(_00842_),
    .DE(_00906_),
    .Q(net991),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[12]$_DFFE_PN_  (.D(_00814_),
    .DE(_00906_),
    .Q(net992),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[13]$_DFFE_PN_  (.D(_00815_),
    .DE(_00906_),
    .Q(net993),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[14]$_DFFE_PN_  (.D(_00816_),
    .DE(_00906_),
    .Q(net994),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[15]$_DFFE_PN_  (.D(_00817_),
    .DE(_00906_),
    .Q(net995),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[16]$_DFFE_PN_  (.D(_00818_),
    .DE(_00906_),
    .Q(net997),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[17]$_DFFE_PN_  (.D(_00819_),
    .DE(_00906_),
    .Q(net998),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[18]$_DFFE_PN_  (.D(_00820_),
    .DE(_00906_),
    .Q(net999),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[19]$_DFFE_PN_  (.D(_00821_),
    .DE(_00906_),
    .Q(net1000),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[1]$_DFFE_PN_  (.D(\hash.CA1.f[1] ),
    .DE(_00906_),
    .Q(net980),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[20]$_DFFE_PN_  (.D(_00822_),
    .DE(_00906_),
    .Q(net1001),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[21]$_DFFE_PN_  (.D(_00823_),
    .DE(_00906_),
    .Q(net1002),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[22]$_DFFE_PN_  (.D(_00825_),
    .DE(_00906_),
    .Q(net1003),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[23]$_DFFE_PN_  (.D(_00826_),
    .DE(_00906_),
    .Q(net1004),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[24]$_DFFE_PN_  (.D(_00827_),
    .DE(_00906_),
    .Q(net1005),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[25]$_DFFE_PN_  (.D(_00828_),
    .DE(_00906_),
    .Q(net1006),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[26]$_DFFE_PN_  (.D(_00829_),
    .DE(_00906_),
    .Q(net1008),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[27]$_DFFE_PN_  (.D(_00830_),
    .DE(_00906_),
    .Q(net1009),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[28]$_DFFE_PN_  (.D(_00831_),
    .DE(_00906_),
    .Q(net1010),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[29]$_DFFE_PN_  (.D(_00832_),
    .DE(_00906_),
    .Q(net1011),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[2]$_DFFE_PN_  (.D(_00813_),
    .DE(_00906_),
    .Q(net981),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[30]$_DFFE_PN_  (.D(_00833_),
    .DE(_00906_),
    .Q(net1012),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[31]$_DFFE_PN_  (.D(_00834_),
    .DE(_00906_),
    .Q(net1013),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[3]$_DFFE_PN_  (.D(_00824_),
    .DE(_00906_),
    .Q(net982),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[4]$_DFFE_PN_  (.D(_00835_),
    .DE(_00906_),
    .Q(net983),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[5]$_DFFE_PN_  (.D(_00836_),
    .DE(_00906_),
    .Q(net984),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[6]$_DFFE_PN_  (.D(_00837_),
    .DE(_00906_),
    .Q(net986),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[7]$_DFFE_PN_  (.D(_00838_),
    .DE(_00906_),
    .Q(net987),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[8]$_DFFE_PN_  (.D(_00839_),
    .DE(_00906_),
    .Q(net988),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[9]$_DFFE_PN_  (.D(_00840_),
    .DE(_00906_),
    .Q(net989),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[0]$_DFFE_PN_  (.D(_00843_),
    .DE(_00906_),
    .Q(net944),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[10]$_DFFE_PN_  (.D(_00844_),
    .DE(_00906_),
    .Q(net955),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[11]$_DFFE_PN_  (.D(_00845_),
    .DE(_00906_),
    .Q(net956),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[12]$_DFFE_PN_  (.D(_00846_),
    .DE(_00906_),
    .Q(net957),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[13]$_DFFE_PN_  (.D(_00847_),
    .DE(_00906_),
    .Q(net958),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[14]$_DFFE_PN_  (.D(_00848_),
    .DE(_00906_),
    .Q(net959),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[15]$_DFFE_PN_  (.D(_00849_),
    .DE(_00906_),
    .Q(net960),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[16]$_DFFE_PN_  (.D(_00850_),
    .DE(_00906_),
    .Q(net961),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[17]$_DFFE_PN_  (.D(_00851_),
    .DE(_00906_),
    .Q(net962),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[18]$_DFFE_PN_  (.D(_00852_),
    .DE(_00906_),
    .Q(net964),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[19]$_DFFE_PN_  (.D(_00853_),
    .DE(_00906_),
    .Q(net965),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[1]$_DFFE_PN_  (.D(_00854_),
    .DE(_00906_),
    .Q(net945),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[20]$_DFFE_PN_  (.D(_00855_),
    .DE(_00906_),
    .Q(net966),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[21]$_DFFE_PN_  (.D(_00856_),
    .DE(_00906_),
    .Q(net967),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[22]$_DFFE_PN_  (.D(_00857_),
    .DE(_00906_),
    .Q(net968),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[23]$_DFFE_PN_  (.D(_00858_),
    .DE(_00906_),
    .Q(net969),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[24]$_DFFE_PN_  (.D(_00859_),
    .DE(_00906_),
    .Q(net970),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[25]$_DFFE_PN_  (.D(_00860_),
    .DE(_00906_),
    .Q(net971),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[26]$_DFFE_PN_  (.D(_00861_),
    .DE(_00906_),
    .Q(net972),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[27]$_DFFE_PN_  (.D(_00862_),
    .DE(_00906_),
    .Q(net973),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[28]$_DFFE_PN_  (.D(_00863_),
    .DE(_00906_),
    .Q(net975),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[29]$_DFFE_PN_  (.D(_00864_),
    .DE(_00906_),
    .Q(net976),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[2]$_DFFE_PN_  (.D(_00865_),
    .DE(_00906_),
    .Q(net946),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[30]$_DFFE_PN_  (.D(_00866_),
    .DE(_00906_),
    .Q(net977),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[31]$_DFFE_PN_  (.D(_00867_),
    .DE(_00906_),
    .Q(net978),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[3]$_DFFE_PN_  (.D(_00868_),
    .DE(_00906_),
    .Q(net947),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[4]$_DFFE_PN_  (.D(_00869_),
    .DE(_00906_),
    .Q(net948),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[5]$_DFFE_PN_  (.D(_00870_),
    .DE(_00906_),
    .Q(net949),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[6]$_DFFE_PN_  (.D(_00871_),
    .DE(_00906_),
    .Q(net950),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[7]$_DFFE_PN_  (.D(_00872_),
    .DE(_00906_),
    .Q(net951),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[8]$_DFFE_PN_  (.D(_00873_),
    .DE(_00906_),
    .Q(net953),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[9]$_DFFE_PN_  (.D(_00874_),
    .DE(_00906_),
    .Q(net954),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[0]$_DFFE_PN_  (.D(_00875_),
    .DE(_00906_),
    .Q(net763),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[10]$_DFFE_PN_  (.D(_00876_),
    .DE(_00906_),
    .Q(net774),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[11]$_DFFE_PN_  (.D(_00877_),
    .DE(_00906_),
    .Q(net785),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[12]$_DFFE_PN_  (.D(_00878_),
    .DE(_00906_),
    .Q(net796),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[13]$_DFFE_PN_  (.D(_00879_),
    .DE(_00906_),
    .Q(net807),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[14]$_DFFE_PN_  (.D(_00880_),
    .DE(_00906_),
    .Q(net818),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[15]$_DFFE_PN_  (.D(_00881_),
    .DE(_00906_),
    .Q(net829),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[16]$_DFFE_PN_  (.D(_00882_),
    .DE(_00906_),
    .Q(net840),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[17]$_DFFE_PN_  (.D(_00883_),
    .DE(_00906_),
    .Q(net851),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[18]$_DFFE_PN_  (.D(_00884_),
    .DE(_00906_),
    .Q(net862),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[19]$_DFFE_PN_  (.D(_00885_),
    .DE(_00906_),
    .Q(net873),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[1]$_DFFE_PN_  (.D(_11749_),
    .DE(_00906_),
    .Q(net874),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[20]$_DFFE_PN_  (.D(_00886_),
    .DE(_00906_),
    .Q(net885),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[21]$_DFFE_PN_  (.D(_00887_),
    .DE(_00906_),
    .Q(net896),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[22]$_DFFE_PN_  (.D(_00888_),
    .DE(_00906_),
    .Q(net907),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[23]$_DFFE_PN_  (.D(_00889_),
    .DE(_00906_),
    .Q(net918),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[24]$_DFFE_PN_  (.D(_00890_),
    .DE(_00906_),
    .Q(net929),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[25]$_DFFE_PN_  (.D(_00891_),
    .DE(_00906_),
    .Q(net936),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[26]$_DFFE_PN_  (.D(_00892_),
    .DE(_00906_),
    .Q(net937),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[27]$_DFFE_PN_  (.D(_00893_),
    .DE(_00906_),
    .Q(net938),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[28]$_DFFE_PN_  (.D(_00894_),
    .DE(_00906_),
    .Q(net939),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[29]$_DFFE_PN_  (.D(_00895_),
    .DE(_00906_),
    .Q(net940),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[2]$_DFFE_PN_  (.D(_00896_),
    .DE(_00906_),
    .Q(net941),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[30]$_DFFE_PN_  (.D(_00897_),
    .DE(_00906_),
    .Q(net942),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[31]$_DFFE_PN_  (.D(_00898_),
    .DE(_00906_),
    .Q(net943),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[3]$_DFFE_PN_  (.D(_00899_),
    .DE(_00906_),
    .Q(net952),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[4]$_DFFE_PN_  (.D(_00900_),
    .DE(_00906_),
    .Q(net963),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[5]$_DFFE_PN_  (.D(_00901_),
    .DE(_00906_),
    .Q(net974),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[6]$_DFFE_PN_  (.D(_00902_),
    .DE(_00906_),
    .Q(net985),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[7]$_DFFE_PN_  (.D(_00903_),
    .DE(_00906_),
    .Q(net996),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[8]$_DFFE_PN_  (.D(_00904_),
    .DE(_00906_),
    .Q(net1007),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[9]$_DFFE_PN_  (.D(_00905_),
    .DE(_00906_),
    .Q(net1018),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p1_cap[0]$_DFF_P_  (.D(\hash.CA1.p1[0] ),
    .Q(\hash.CA2.p1[0] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[10]$_DFF_P_  (.D(\hash.CA1.p1[10] ),
    .Q(\hash.CA2.p1[10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[11]$_DFF_P_  (.D(\hash.CA1.p1[11] ),
    .Q(\hash.CA2.p1[11] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[12]$_DFF_P_  (.D(\hash.CA1.p1[12] ),
    .Q(\hash.CA2.p1[12] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[13]$_DFF_P_  (.D(\hash.CA1.p1[13] ),
    .Q(\hash.CA2.p1[13] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[14]$_DFF_P_  (.D(\hash.CA1.p1[14] ),
    .Q(\hash.CA2.p1[14] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[15]$_DFF_P_  (.D(\hash.CA1.p1[15] ),
    .Q(\hash.CA2.p1[15] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[16]$_DFF_P_  (.D(\hash.CA1.p1[16] ),
    .Q(\hash.CA2.p1[16] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[17]$_DFF_P_  (.D(\hash.CA1.p1[17] ),
    .Q(\hash.CA2.p1[17] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[18]$_DFF_P_  (.D(\hash.CA1.p1[18] ),
    .Q(\hash.CA2.p1[18] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[19]$_DFF_P_  (.D(\hash.CA1.p1[19] ),
    .Q(\hash.CA2.p1[19] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[1]$_DFF_P_  (.D(\hash.CA1.p1[1] ),
    .Q(\hash.CA2.p1[1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[20]$_DFF_P_  (.D(\hash.CA1.p1[20] ),
    .Q(\hash.CA2.p1[20] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[21]$_DFF_P_  (.D(\hash.CA1.p1[21] ),
    .Q(\hash.CA2.p1[21] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[22]$_DFF_P_  (.D(\hash.CA1.p1[22] ),
    .Q(\hash.CA2.p1[22] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[23]$_DFF_P_  (.D(\hash.CA1.p1[23] ),
    .Q(\hash.CA2.p1[23] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[24]$_DFF_P_  (.D(\hash.CA1.p1[24] ),
    .Q(\hash.CA2.p1[24] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[25]$_DFF_P_  (.D(\hash.CA1.p1[25] ),
    .Q(\hash.CA2.p1[25] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[26]$_DFF_P_  (.D(\hash.CA1.p1[26] ),
    .Q(\hash.CA2.p1[26] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[27]$_DFF_P_  (.D(\hash.CA1.p1[27] ),
    .Q(\hash.CA2.p1[27] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[28]$_DFF_P_  (.D(\hash.CA1.p1[28] ),
    .Q(\hash.CA2.p1[28] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[29]$_DFF_P_  (.D(\hash.CA1.p1[29] ),
    .Q(\hash.CA2.p1[29] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[2]$_DFF_P_  (.D(\hash.CA1.p1[2] ),
    .Q(\hash.CA2.p1[2] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[30]$_DFF_P_  (.D(\hash.CA1.p1[30] ),
    .Q(\hash.CA2.p1[30] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[31]$_DFF_P_  (.D(\hash.CA1.p1[31] ),
    .Q(\hash.CA2.p1[31] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[3]$_DFF_P_  (.D(\hash.CA1.p1[3] ),
    .Q(\hash.CA2.p1[3] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[4]$_DFF_P_  (.D(\hash.CA1.p1[4] ),
    .Q(\hash.CA2.p1[4] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[5]$_DFF_P_  (.D(\hash.CA1.p1[5] ),
    .Q(\hash.CA2.p1[5] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[6]$_DFF_P_  (.D(\hash.CA1.p1[6] ),
    .Q(\hash.CA2.p1[6] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[7]$_DFF_P_  (.D(\hash.CA1.p1[7] ),
    .Q(\hash.CA2.p1[7] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[8]$_DFF_P_  (.D(\hash.CA1.p1[8] ),
    .Q(\hash.CA2.p1[8] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[9]$_DFF_P_  (.D(\hash.CA1.p1[9] ),
    .Q(\hash.CA2.p1[9] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[0]$_DFF_P_  (.D(\hash.CA1.p2[0] ),
    .Q(\hash.CA2.S1.X[0] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[10]$_DFF_P_  (.D(\hash.CA1.p2[10] ),
    .Q(\hash.CA2.S1.X[10] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[11]$_DFF_P_  (.D(\hash.CA1.p2[11] ),
    .Q(\hash.CA2.S1.X[11] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[12]$_DFF_P_  (.D(\hash.CA1.p2[12] ),
    .Q(\hash.CA2.S1.X[12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[13]$_DFF_P_  (.D(\hash.CA1.p2[13] ),
    .Q(\hash.CA2.S1.X[13] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[14]$_DFF_P_  (.D(\hash.CA1.p2[14] ),
    .Q(\hash.CA2.S1.X[14] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[15]$_DFF_P_  (.D(\hash.CA1.p2[15] ),
    .Q(\hash.CA2.S1.X[15] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[16]$_DFF_P_  (.D(\hash.CA1.p2[16] ),
    .Q(\hash.CA2.S1.X[16] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[17]$_DFF_P_  (.D(\hash.CA1.p2[17] ),
    .Q(\hash.CA2.S1.X[17] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[18]$_DFF_P_  (.D(\hash.CA1.p2[18] ),
    .Q(\hash.CA2.S1.X[18] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[19]$_DFF_P_  (.D(\hash.CA1.p2[19] ),
    .Q(\hash.CA2.S1.X[19] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[1]$_DFF_P_  (.D(\hash.CA1.p2[1] ),
    .Q(\hash.CA2.S1.X[1] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[20]$_DFF_P_  (.D(\hash.CA1.p2[20] ),
    .Q(\hash.CA2.S1.X[20] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[21]$_DFF_P_  (.D(\hash.CA1.p2[21] ),
    .Q(\hash.CA2.S1.X[21] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[22]$_DFF_P_  (.D(\hash.CA1.p2[22] ),
    .Q(\hash.CA2.S1.X[22] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[23]$_DFF_P_  (.D(\hash.CA1.p2[23] ),
    .Q(\hash.CA2.S1.X[23] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[24]$_DFF_P_  (.D(\hash.CA1.p2[24] ),
    .Q(\hash.CA2.S1.X[24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[25]$_DFF_P_  (.D(\hash.CA1.p2[25] ),
    .Q(\hash.CA2.S1.X[25] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[26]$_DFF_P_  (.D(\hash.CA1.p2[26] ),
    .Q(\hash.CA2.S1.X[26] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[27]$_DFF_P_  (.D(\hash.CA1.p2[27] ),
    .Q(\hash.CA2.S1.X[27] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[28]$_DFF_P_  (.D(\hash.CA1.p2[28] ),
    .Q(\hash.CA2.S1.X[28] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[29]$_DFF_P_  (.D(\hash.CA1.p2[29] ),
    .Q(\hash.CA2.S1.X[29] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[2]$_DFF_P_  (.D(\hash.CA1.p2[2] ),
    .Q(\hash.CA2.S1.X[2] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[30]$_DFF_P_  (.D(\hash.CA1.p2[30] ),
    .Q(\hash.CA2.S1.X[30] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[31]$_DFF_P_  (.D(\hash.CA1.p2[31] ),
    .Q(\hash.CA2.S1.X[31] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[3]$_DFF_P_  (.D(\hash.CA1.p2[3] ),
    .Q(\hash.CA2.S1.X[3] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[4]$_DFF_P_  (.D(\hash.CA1.p2[4] ),
    .Q(\hash.CA2.S1.X[4] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[5]$_DFF_P_  (.D(\hash.CA1.p2[5] ),
    .Q(\hash.CA2.S1.X[5] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[6]$_DFF_P_  (.D(\hash.CA1.p2[6] ),
    .Q(\hash.CA2.S1.X[6] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[7]$_DFF_P_  (.D(\hash.CA1.p2[7] ),
    .Q(\hash.CA2.S1.X[7] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[8]$_DFF_P_  (.D(\hash.CA1.p2[8] ),
    .Q(\hash.CA2.S1.X[8] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[9]$_DFF_P_  (.D(\hash.CA1.p2[9] ),
    .Q(\hash.CA2.S1.X[9] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[0]$_DFF_P_  (.D(\hash.CA1.p3[0] ),
    .Q(\hash.CA2.p3[0] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[10]$_DFF_P_  (.D(\hash.CA1.p3[10] ),
    .Q(\hash.CA2.p3[10] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[11]$_DFF_P_  (.D(\hash.CA1.p3[11] ),
    .Q(\hash.CA2.p3[11] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[12]$_DFF_P_  (.D(\hash.CA1.p3[12] ),
    .Q(\hash.CA2.p3[12] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[13]$_DFF_P_  (.D(\hash.CA1.p3[13] ),
    .Q(\hash.CA2.p3[13] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[14]$_DFF_P_  (.D(\hash.CA1.p3[14] ),
    .Q(\hash.CA2.p3[14] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[15]$_DFF_P_  (.D(\hash.CA1.p3[15] ),
    .Q(\hash.CA2.p3[15] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[16]$_DFF_P_  (.D(\hash.CA1.p3[16] ),
    .Q(\hash.CA2.p3[16] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[17]$_DFF_P_  (.D(\hash.CA1.p3[17] ),
    .Q(\hash.CA2.p3[17] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[18]$_DFF_P_  (.D(\hash.CA1.p3[18] ),
    .Q(\hash.CA2.p3[18] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[19]$_DFF_P_  (.D(\hash.CA1.p3[19] ),
    .Q(\hash.CA2.p3[19] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[1]$_DFF_P_  (.D(\hash.CA1.p3[1] ),
    .Q(\hash.CA2.p3[1] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[20]$_DFF_P_  (.D(\hash.CA1.p3[20] ),
    .Q(\hash.CA2.p3[20] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[21]$_DFF_P_  (.D(\hash.CA1.p3[21] ),
    .Q(\hash.CA2.p3[21] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[22]$_DFF_P_  (.D(\hash.CA1.p3[22] ),
    .Q(\hash.CA2.p3[22] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[23]$_DFF_P_  (.D(\hash.CA1.p3[23] ),
    .Q(\hash.CA2.p3[23] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[24]$_DFF_P_  (.D(\hash.CA1.p3[24] ),
    .Q(\hash.CA2.p3[24] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[25]$_DFF_P_  (.D(\hash.CA1.p3[25] ),
    .Q(\hash.CA2.p3[25] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[26]$_DFF_P_  (.D(\hash.CA1.p3[26] ),
    .Q(\hash.CA2.p3[26] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[27]$_DFF_P_  (.D(\hash.CA1.p3[27] ),
    .Q(\hash.CA2.p3[27] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[28]$_DFF_P_  (.D(\hash.CA1.p3[28] ),
    .Q(\hash.CA2.p3[28] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[29]$_DFF_P_  (.D(\hash.CA1.p3[29] ),
    .Q(\hash.CA2.p3[29] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[2]$_DFF_P_  (.D(\hash.CA1.p3[2] ),
    .Q(\hash.CA2.p3[2] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[30]$_DFF_P_  (.D(\hash.CA1.p3[30] ),
    .Q(\hash.CA2.p3[30] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[31]$_DFF_P_  (.D(\hash.CA1.p3[31] ),
    .Q(\hash.CA2.p3[31] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[3]$_DFF_P_  (.D(\hash.CA1.p3[3] ),
    .Q(\hash.CA2.p3[3] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[4]$_DFF_P_  (.D(\hash.CA1.p3[4] ),
    .Q(\hash.CA2.p3[4] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[5]$_DFF_P_  (.D(\hash.CA1.p3[5] ),
    .Q(\hash.CA2.p3[5] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[6]$_DFF_P_  (.D(\hash.CA1.p3[6] ),
    .Q(\hash.CA2.p3[6] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[7]$_DFF_P_  (.D(\hash.CA1.p3[7] ),
    .Q(\hash.CA2.p3[7] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[8]$_DFF_P_  (.D(\hash.CA1.p3[8] ),
    .Q(\hash.CA2.p3[8] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[9]$_DFF_P_  (.D(\hash.CA1.p3[9] ),
    .Q(\hash.CA2.p3[9] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[0]$_DFF_P_  (.D(\hash.CA1.p4[0] ),
    .Q(\hash.CA2.p4[0] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[10]$_DFF_P_  (.D(\hash.CA1.p4[10] ),
    .Q(\hash.CA2.p4[10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[11]$_DFF_P_  (.D(\hash.CA1.p4[11] ),
    .Q(\hash.CA2.p4[11] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[12]$_DFF_P_  (.D(\hash.CA1.p4[12] ),
    .Q(\hash.CA2.p4[12] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[13]$_DFF_P_  (.D(\hash.CA1.p4[13] ),
    .Q(\hash.CA2.p4[13] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[14]$_DFF_P_  (.D(\hash.CA1.p4[14] ),
    .Q(\hash.CA2.p4[14] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[15]$_DFF_P_  (.D(\hash.CA1.p4[15] ),
    .Q(\hash.CA2.p4[15] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[16]$_DFF_P_  (.D(\hash.CA1.p4[16] ),
    .Q(\hash.CA2.p4[16] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[17]$_DFF_P_  (.D(\hash.CA1.p4[17] ),
    .Q(\hash.CA2.p4[17] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[18]$_DFF_P_  (.D(\hash.CA1.p4[18] ),
    .Q(\hash.CA2.p4[18] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[19]$_DFF_P_  (.D(\hash.CA1.p4[19] ),
    .Q(\hash.CA2.p4[19] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[1]$_DFF_P_  (.D(\hash.CA1.p4[1] ),
    .Q(\hash.CA2.p4[1] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[20]$_DFF_P_  (.D(\hash.CA1.p4[20] ),
    .Q(\hash.CA2.p4[20] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[21]$_DFF_P_  (.D(\hash.CA1.p4[21] ),
    .Q(\hash.CA2.p4[21] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[22]$_DFF_P_  (.D(\hash.CA1.p4[22] ),
    .Q(\hash.CA2.p4[22] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[23]$_DFF_P_  (.D(\hash.CA1.p4[23] ),
    .Q(\hash.CA2.p4[23] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[24]$_DFF_P_  (.D(\hash.CA1.p4[24] ),
    .Q(\hash.CA2.p4[24] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[25]$_DFF_P_  (.D(\hash.CA1.p4[25] ),
    .Q(\hash.CA2.p4[25] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[26]$_DFF_P_  (.D(\hash.CA1.p4[26] ),
    .Q(\hash.CA2.p4[26] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[27]$_DFF_P_  (.D(\hash.CA1.p4[27] ),
    .Q(\hash.CA2.p4[27] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[28]$_DFF_P_  (.D(\hash.CA1.p4[28] ),
    .Q(\hash.CA2.p4[28] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[29]$_DFF_P_  (.D(\hash.CA1.p4[29] ),
    .Q(\hash.CA2.p4[29] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[2]$_DFF_P_  (.D(\hash.CA1.p4[2] ),
    .Q(\hash.CA2.p4[2] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[30]$_DFF_P_  (.D(\hash.CA1.p4[30] ),
    .Q(\hash.CA2.p4[30] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[31]$_DFF_P_  (.D(\hash.CA1.p4[31] ),
    .Q(\hash.CA2.p4[31] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[3]$_DFF_P_  (.D(\hash.CA1.p4[3] ),
    .Q(\hash.CA2.p4[3] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[4]$_DFF_P_  (.D(\hash.CA1.p4[4] ),
    .Q(\hash.CA2.p4[4] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[5]$_DFF_P_  (.D(\hash.CA1.p4[5] ),
    .Q(\hash.CA2.p4[5] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[6]$_DFF_P_  (.D(\hash.CA1.p4[6] ),
    .Q(\hash.CA2.p4[6] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[7]$_DFF_P_  (.D(\hash.CA1.p4[7] ),
    .Q(\hash.CA2.p4[7] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[8]$_DFF_P_  (.D(\hash.CA1.p4[8] ),
    .Q(\hash.CA2.p4[8] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[9]$_DFF_P_  (.D(\hash.CA1.p4[9] ),
    .Q(\hash.CA2.p4[9] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[0]$_DFF_P_  (.D(\hash.CA1.p5[0] ),
    .Q(\hash.CA2.p5[0] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[10]$_DFF_P_  (.D(\hash.CA1.p5[10] ),
    .Q(\hash.CA2.p5[10] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[11]$_DFF_P_  (.D(\hash.CA1.p5[11] ),
    .Q(\hash.CA2.p5[11] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[12]$_DFF_P_  (.D(\hash.CA1.p5[12] ),
    .Q(\hash.CA2.p5[12] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[13]$_DFF_P_  (.D(\hash.CA1.p5[13] ),
    .Q(\hash.CA2.p5[13] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[14]$_DFF_P_  (.D(\hash.CA1.p5[14] ),
    .Q(\hash.CA2.p5[14] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[15]$_DFF_P_  (.D(\hash.CA1.p5[15] ),
    .Q(\hash.CA2.p5[15] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[16]$_DFF_P_  (.D(\hash.CA1.p5[16] ),
    .Q(\hash.CA2.p5[16] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[17]$_DFF_P_  (.D(\hash.CA1.p5[17] ),
    .Q(\hash.CA2.p5[17] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[18]$_DFF_P_  (.D(\hash.CA1.p5[18] ),
    .Q(\hash.CA2.p5[18] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[19]$_DFF_P_  (.D(\hash.CA1.p5[19] ),
    .Q(\hash.CA2.p5[19] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[1]$_DFF_P_  (.D(\hash.CA1.p5[1] ),
    .Q(\hash.CA2.p5[1] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[20]$_DFF_P_  (.D(\hash.CA1.p5[20] ),
    .Q(\hash.CA2.p5[20] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[21]$_DFF_P_  (.D(\hash.CA1.p5[21] ),
    .Q(\hash.CA2.p5[21] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[22]$_DFF_P_  (.D(\hash.CA1.p5[22] ),
    .Q(\hash.CA2.p5[22] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[23]$_DFF_P_  (.D(\hash.CA1.p5[23] ),
    .Q(\hash.CA2.p5[23] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[24]$_DFF_P_  (.D(\hash.CA1.p5[24] ),
    .Q(\hash.CA2.p5[24] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[25]$_DFF_P_  (.D(\hash.CA1.p5[25] ),
    .Q(\hash.CA2.p5[25] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[26]$_DFF_P_  (.D(\hash.CA1.p5[26] ),
    .Q(\hash.CA2.p5[26] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[27]$_DFF_P_  (.D(\hash.CA1.p5[27] ),
    .Q(\hash.CA2.p5[27] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[28]$_DFF_P_  (.D(\hash.CA1.p5[28] ),
    .Q(\hash.CA2.p5[28] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[29]$_DFF_P_  (.D(\hash.CA1.p5[29] ),
    .Q(\hash.CA2.p5[29] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[2]$_DFF_P_  (.D(\hash.CA1.p5[2] ),
    .Q(\hash.CA2.p5[2] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[30]$_DFF_P_  (.D(\hash.CA1.p5[30] ),
    .Q(\hash.CA2.p5[30] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[31]$_DFF_P_  (.D(\hash.CA1.p5[31] ),
    .Q(\hash.CA2.p5[31] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[3]$_DFF_P_  (.D(\hash.CA1.p5[3] ),
    .Q(\hash.CA2.p5[3] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[4]$_DFF_P_  (.D(\hash.CA1.p5[4] ),
    .Q(\hash.CA2.p5[4] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[5]$_DFF_P_  (.D(\hash.CA1.p5[5] ),
    .Q(\hash.CA2.p5[5] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[6]$_DFF_P_  (.D(\hash.CA1.p5[6] ),
    .Q(\hash.CA2.p5[6] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[7]$_DFF_P_  (.D(\hash.CA1.p5[7] ),
    .Q(\hash.CA2.p5[7] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[8]$_DFF_P_  (.D(\hash.CA1.p5[8] ),
    .Q(\hash.CA2.p5[8] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[9]$_DFF_P_  (.D(\hash.CA1.p5[9] ),
    .Q(\hash.CA2.p5[9] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[0]$_SDFF_PP0_  (.D(_00969_),
    .Q(\hash.CA1.k_i1[0] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[10]$_SDFF_PP1_  (.D(_00970_),
    .Q(\hash.CA1.k_i1[10] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[11]$_SDFF_PP1_  (.D(_00971_),
    .Q(\hash.CA1.k_i1[11] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[12]$_SDFF_PP0_  (.D(_00972_),
    .Q(\hash.CA1.k_i1[12] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[13]$_SDFF_PP1_  (.D(_00973_),
    .Q(\hash.CA1.k_i1[13] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[14]$_SDFF_PP0_  (.D(_00974_),
    .Q(\hash.CA1.k_i1[14] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[15]$_SDFF_PP0_  (.D(_00975_),
    .Q(\hash.CA1.k_i1[15] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[16]$_SDFF_PP0_  (.D(_00976_),
    .Q(\hash.CA1.k_i1[16] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[17]$_SDFF_PP1_  (.D(_00977_),
    .Q(\hash.CA1.k_i1[17] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[18]$_SDFF_PP0_  (.D(_00978_),
    .Q(\hash.CA1.k_i1[18] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[19]$_SDFF_PP1_  (.D(_00979_),
    .Q(\hash.CA1.k_i1[19] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[1]$_SDFF_PP0_  (.D(_00980_),
    .Q(\hash.CA1.k_i1[1] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[20]$_SDFF_PP0_  (.D(_00981_),
    .Q(\hash.CA1.k_i1[20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[21]$_SDFF_PP0_  (.D(_00982_),
    .Q(\hash.CA1.k_i1[21] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[22]$_SDFF_PP0_  (.D(_00983_),
    .Q(\hash.CA1.k_i1[22] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[23]$_SDFF_PP1_  (.D(_00984_),
    .Q(\hash.CA1.k_i1[23] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[24]$_SDFF_PP0_  (.D(_00985_),
    .Q(\hash.CA1.k_i1[24] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[25]$_SDFF_PP1_  (.D(_00986_),
    .Q(\hash.CA1.k_i1[25] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[26]$_SDFF_PP0_  (.D(_00987_),
    .Q(\hash.CA1.k_i1[26] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[27]$_SDFF_PP0_  (.D(_00988_),
    .Q(\hash.CA1.k_i1[27] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[28]$_SDFF_PP0_  (.D(_00989_),
    .Q(\hash.CA1.k_i1[28] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[29]$_SDFF_PP0_  (.D(_00990_),
    .Q(\hash.CA1.k_i1[29] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[2]$_SDFF_PP0_  (.D(_00991_),
    .Q(\hash.CA1.k_i1[2] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[30]$_SDFF_PP1_  (.D(_00992_),
    .Q(\hash.CA1.k_i1[30] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[31]$_SDFF_PP0_  (.D(_00993_),
    .Q(\hash.CA1.k_i1[31] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[3]$_SDFF_PP1_  (.D(_00994_),
    .Q(\hash.CA1.k_i1[3] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[4]$_SDFF_PP1_  (.D(_00995_),
    .Q(\hash.CA1.k_i1[4] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[5]$_SDFF_PP0_  (.D(_00996_),
    .Q(\hash.CA1.k_i1[5] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[6]$_SDFF_PP0_  (.D(_00997_),
    .Q(\hash.CA1.k_i1[6] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[7]$_SDFF_PP1_  (.D(_00998_),
    .Q(\hash.CA1.k_i1[7] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[8]$_SDFF_PP1_  (.D(_00999_),
    .Q(\hash.CA1.k_i1[8] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[9]$_SDFF_PP1_  (.D(_01000_),
    .Q(\hash.CA1.k_i1[9] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[0]$_SDFF_PP1_  (.D(_01001_),
    .Q(\hash.CA1.k_i2[0] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[10]$_SDFF_PP1_  (.D(_01002_),
    .Q(\hash.CA1.k_i2[10] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[11]$_SDFF_PP0_  (.D(_01003_),
    .Q(\hash.CA1.k_i2[11] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[12]$_SDFF_PP0_  (.D(_01004_),
    .Q(\hash.CA1.k_i2[12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[13]$_SDFF_PP0_  (.D(_01005_),
    .Q(\hash.CA1.k_i2[13] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[14]$_SDFF_PP1_  (.D(_01006_),
    .Q(\hash.CA1.k_i2[14] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[15]$_SDFF_PP0_  (.D(_01007_),
    .Q(\hash.CA1.k_i2[15] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[16]$_SDFF_PP1_  (.D(_01008_),
    .Q(\hash.CA1.k_i2[16] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[17]$_SDFF_PP1_  (.D(_01009_),
    .Q(\hash.CA1.k_i2[17] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[18]$_SDFF_PP1_  (.D(_01010_),
    .Q(\hash.CA1.k_i2[18] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[19]$_SDFF_PP0_  (.D(_01011_),
    .Q(\hash.CA1.k_i2[19] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[1]$_SDFF_PP0_  (.D(_01012_),
    .Q(\hash.CA1.k_i2[1] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[20]$_SDFF_PP1_  (.D(_01013_),
    .Q(\hash.CA1.k_i2[20] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[21]$_SDFF_PP1_  (.D(_01014_),
    .Q(\hash.CA1.k_i2[21] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[22]$_SDFF_PP0_  (.D(_01015_),
    .Q(\hash.CA1.k_i2[22] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[23]$_SDFF_PP0_  (.D(_01016_),
    .Q(\hash.CA1.k_i2[23] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[24]$_SDFF_PP1_  (.D(_01017_),
    .Q(\hash.CA1.k_i2[24] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[25]$_SDFF_PP0_  (.D(_01018_),
    .Q(\hash.CA1.k_i2[25] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[26]$_SDFF_PP0_  (.D(_01019_),
    .Q(\hash.CA1.k_i2[26] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[27]$_SDFF_PP0_  (.D(_01020_),
    .Q(\hash.CA1.k_i2[27] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[28]$_SDFF_PP1_  (.D(_01021_),
    .Q(\hash.CA1.k_i2[28] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[29]$_SDFF_PP1_  (.D(_01022_),
    .Q(\hash.CA1.k_i2[29] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[2]$_SDFF_PP0_  (.D(_01023_),
    .Q(\hash.CA1.k_i2[2] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[30]$_SDFF_PP1_  (.D(_01024_),
    .Q(\hash.CA1.k_i2[30] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[31]$_SDFF_PP0_  (.D(_01025_),
    .Q(\hash.CA1.k_i2[31] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[3]$_SDFF_PP0_  (.D(_01026_),
    .Q(\hash.CA1.k_i2[3] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[4]$_SDFF_PP1_  (.D(_01027_),
    .Q(\hash.CA1.k_i2[4] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[5]$_SDFF_PP0_  (.D(_01028_),
    .Q(\hash.CA1.k_i2[5] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[6]$_SDFF_PP0_  (.D(_01029_),
    .Q(\hash.CA1.k_i2[6] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[7]$_SDFF_PP1_  (.D(_01030_),
    .Q(\hash.CA1.k_i2[7] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[8]$_SDFF_PP0_  (.D(_01031_),
    .Q(\hash.CA1.k_i2[8] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[9]$_SDFF_PP0_  (.D(_01032_),
    .Q(\hash.CA1.k_i2[9] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_4 \ready$_DFF_P_  (.D(ready_dash),
    .Q(net1019),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \ready_dash$_SDFF_PP0_  (.D(_01033_),
    .Q(ready_dash),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_4 \reset_hash$_DFF_P_  (.D(net762),
    .Q(reset_hash),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_4 \reset_hash_dash$_DFF_P_  (.D(net525),
    .Q(\hash.reset ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][0]$_DFFE_PP_  (.D(_00129_),
    .DE(_00127_),
    .Q(\w[0][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][10]$_DFFE_PP_  (.D(_00130_),
    .DE(_00127_),
    .Q(\w[0][10] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][11]$_DFFE_PP_  (.D(_00131_),
    .DE(_00127_),
    .Q(\w[0][11] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][12]$_DFFE_PP_  (.D(_00132_),
    .DE(_00127_),
    .Q(\w[0][12] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][13]$_DFFE_PP_  (.D(_00133_),
    .DE(_00127_),
    .Q(\w[0][13] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][14]$_DFFE_PP_  (.D(_00134_),
    .DE(_00127_),
    .Q(\w[0][14] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][15]$_DFFE_PP_  (.D(_00135_),
    .DE(_00127_),
    .Q(\w[0][15] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][16]$_DFFE_PP_  (.D(_00136_),
    .DE(_00127_),
    .Q(\w[0][16] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][17]$_DFFE_PP_  (.D(_00137_),
    .DE(_00127_),
    .Q(\w[0][17] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][18]$_DFFE_PP_  (.D(_00138_),
    .DE(_00127_),
    .Q(\w[0][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][19]$_DFFE_PP_  (.D(_00139_),
    .DE(_00127_),
    .Q(\w[0][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][1]$_DFFE_PP_  (.D(_00140_),
    .DE(_00127_),
    .Q(\w[0][1] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][20]$_DFFE_PP_  (.D(_00141_),
    .DE(_00127_),
    .Q(\w[0][20] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][21]$_DFFE_PP_  (.D(_00142_),
    .DE(_00127_),
    .Q(\w[0][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][22]$_DFFE_PP_  (.D(_00143_),
    .DE(_00127_),
    .Q(\w[0][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][23]$_DFFE_PP_  (.D(_00144_),
    .DE(_00127_),
    .Q(\w[0][23] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][24]$_DFFE_PP_  (.D(_00145_),
    .DE(_00127_),
    .Q(\w[0][24] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][25]$_DFFE_PP_  (.D(_00146_),
    .DE(_00127_),
    .Q(\w[0][25] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][26]$_DFFE_PP_  (.D(_00147_),
    .DE(_00127_),
    .Q(\w[0][26] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][27]$_DFFE_PP_  (.D(_00148_),
    .DE(_00127_),
    .Q(\w[0][27] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][28]$_DFFE_PP_  (.D(_00149_),
    .DE(_00127_),
    .Q(\w[0][28] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][29]$_DFFE_PP_  (.D(_00150_),
    .DE(_00127_),
    .Q(\w[0][29] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][2]$_DFFE_PP_  (.D(_00151_),
    .DE(_00127_),
    .Q(\w[0][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][30]$_DFFE_PP_  (.D(_00152_),
    .DE(_00127_),
    .Q(\w[0][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][31]$_DFFE_PP_  (.D(_00153_),
    .DE(_00127_),
    .Q(\w[0][31] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][3]$_DFFE_PP_  (.D(_00154_),
    .DE(_00127_),
    .Q(\w[0][3] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][4]$_DFFE_PP_  (.D(_00155_),
    .DE(_00127_),
    .Q(\w[0][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][5]$_DFFE_PP_  (.D(_00156_),
    .DE(_00127_),
    .Q(\w[0][5] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][6]$_DFFE_PP_  (.D(_00157_),
    .DE(_00127_),
    .Q(\w[0][6] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][7]$_DFFE_PP_  (.D(_00158_),
    .DE(_00127_),
    .Q(\w[0][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][8]$_DFFE_PP_  (.D(_00159_),
    .DE(_00127_),
    .Q(\w[0][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][9]$_DFFE_PP_  (.D(_00160_),
    .DE(_00127_),
    .Q(\w[0][9] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][0]$_DFFE_PP_  (.D(_00161_),
    .DE(_00126_),
    .Q(\w[10][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][10]$_DFFE_PP_  (.D(_00162_),
    .DE(_00126_),
    .Q(\w[10][10] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][11]$_DFFE_PP_  (.D(_00163_),
    .DE(_00126_),
    .Q(\w[10][11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][12]$_DFFE_PP_  (.D(_00164_),
    .DE(_00126_),
    .Q(\w[10][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][13]$_DFFE_PP_  (.D(_00165_),
    .DE(_00126_),
    .Q(\w[10][13] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][14]$_DFFE_PP_  (.D(_00166_),
    .DE(_00126_),
    .Q(\w[10][14] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][15]$_DFFE_PP_  (.D(_00167_),
    .DE(_00126_),
    .Q(\w[10][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][16]$_DFFE_PP_  (.D(_00168_),
    .DE(_00126_),
    .Q(\w[10][16] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][17]$_DFFE_PP_  (.D(_00169_),
    .DE(_00126_),
    .Q(\w[10][17] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][18]$_DFFE_PP_  (.D(_00170_),
    .DE(_00126_),
    .Q(\w[10][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][19]$_DFFE_PP_  (.D(_00171_),
    .DE(_00126_),
    .Q(\w[10][19] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][1]$_DFFE_PP_  (.D(_00172_),
    .DE(_00126_),
    .Q(\w[10][1] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][20]$_DFFE_PP_  (.D(_00173_),
    .DE(_00126_),
    .Q(\w[10][20] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][21]$_DFFE_PP_  (.D(_00174_),
    .DE(_00126_),
    .Q(\w[10][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][22]$_DFFE_PP_  (.D(_00175_),
    .DE(_00126_),
    .Q(\w[10][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][23]$_DFFE_PP_  (.D(_00176_),
    .DE(_00126_),
    .Q(\w[10][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][24]$_DFFE_PP_  (.D(_00177_),
    .DE(_00126_),
    .Q(\w[10][24] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][25]$_DFFE_PP_  (.D(_00178_),
    .DE(_00126_),
    .Q(\w[10][25] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][26]$_DFFE_PP_  (.D(_00179_),
    .DE(_00126_),
    .Q(\w[10][26] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][27]$_DFFE_PP_  (.D(_00180_),
    .DE(_00126_),
    .Q(\w[10][27] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][28]$_DFFE_PP_  (.D(_00181_),
    .DE(_00126_),
    .Q(\w[10][28] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][29]$_DFFE_PP_  (.D(_00182_),
    .DE(_00126_),
    .Q(\w[10][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][2]$_DFFE_PP_  (.D(_00183_),
    .DE(_00126_),
    .Q(\w[10][2] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][30]$_DFFE_PP_  (.D(_00184_),
    .DE(_00126_),
    .Q(\w[10][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][31]$_DFFE_PP_  (.D(_00185_),
    .DE(_00126_),
    .Q(\w[10][31] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][3]$_DFFE_PP_  (.D(_00186_),
    .DE(_00126_),
    .Q(\w[10][3] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][4]$_DFFE_PP_  (.D(_00187_),
    .DE(_00126_),
    .Q(\w[10][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][5]$_DFFE_PP_  (.D(_00188_),
    .DE(_00126_),
    .Q(\w[10][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][6]$_DFFE_PP_  (.D(_00189_),
    .DE(_00126_),
    .Q(\w[10][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][7]$_DFFE_PP_  (.D(_00190_),
    .DE(_00126_),
    .Q(\w[10][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][8]$_DFFE_PP_  (.D(_00191_),
    .DE(_00126_),
    .Q(\w[10][8] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][9]$_DFFE_PP_  (.D(_00192_),
    .DE(_00126_),
    .Q(\w[10][9] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][0]$_DFFE_PP_  (.D(_00193_),
    .DE(_00095_),
    .Q(\w[11][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][10]$_DFFE_PP_  (.D(_00194_),
    .DE(_00095_),
    .Q(\w[11][10] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][11]$_DFFE_PP_  (.D(_00195_),
    .DE(_00095_),
    .Q(\w[11][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][12]$_DFFE_PP_  (.D(_00196_),
    .DE(_00095_),
    .Q(\w[11][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][13]$_DFFE_PP_  (.D(_00197_),
    .DE(_00095_),
    .Q(\w[11][13] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][14]$_DFFE_PP_  (.D(_00198_),
    .DE(_00095_),
    .Q(\w[11][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][15]$_DFFE_PP_  (.D(_00199_),
    .DE(_00095_),
    .Q(\w[11][15] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][16]$_DFFE_PP_  (.D(_00200_),
    .DE(_00095_),
    .Q(\w[11][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][17]$_DFFE_PP_  (.D(_00201_),
    .DE(_00095_),
    .Q(\w[11][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][18]$_DFFE_PP_  (.D(_00202_),
    .DE(_00095_),
    .Q(\w[11][18] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][19]$_DFFE_PP_  (.D(_00203_),
    .DE(_00095_),
    .Q(\w[11][19] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][1]$_DFFE_PP_  (.D(_00204_),
    .DE(_00095_),
    .Q(\w[11][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][20]$_DFFE_PP_  (.D(_00205_),
    .DE(_00095_),
    .Q(\w[11][20] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][21]$_DFFE_PP_  (.D(_00206_),
    .DE(_00095_),
    .Q(\w[11][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][22]$_DFFE_PP_  (.D(_00207_),
    .DE(_00095_),
    .Q(\w[11][22] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][23]$_DFFE_PP_  (.D(_00208_),
    .DE(_00095_),
    .Q(\w[11][23] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][24]$_DFFE_PP_  (.D(_00209_),
    .DE(_00095_),
    .Q(\w[11][24] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][25]$_DFFE_PP_  (.D(_00210_),
    .DE(_00095_),
    .Q(\w[11][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][26]$_DFFE_PP_  (.D(_00211_),
    .DE(_00095_),
    .Q(\w[11][26] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][27]$_DFFE_PP_  (.D(_00212_),
    .DE(_00095_),
    .Q(\w[11][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][28]$_DFFE_PP_  (.D(_00213_),
    .DE(_00095_),
    .Q(\w[11][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][29]$_DFFE_PP_  (.D(_00214_),
    .DE(_00095_),
    .Q(\w[11][29] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][2]$_DFFE_PP_  (.D(_00215_),
    .DE(_00095_),
    .Q(\w[11][2] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][30]$_DFFE_PP_  (.D(_00216_),
    .DE(_00095_),
    .Q(\w[11][30] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][31]$_DFFE_PP_  (.D(_00217_),
    .DE(_00095_),
    .Q(\w[11][31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][3]$_DFFE_PP_  (.D(_00218_),
    .DE(_00095_),
    .Q(\w[11][3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][4]$_DFFE_PP_  (.D(_00219_),
    .DE(_00095_),
    .Q(\w[11][4] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][5]$_DFFE_PP_  (.D(_00220_),
    .DE(_00095_),
    .Q(\w[11][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][6]$_DFFE_PP_  (.D(_00221_),
    .DE(_00095_),
    .Q(\w[11][6] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][7]$_DFFE_PP_  (.D(_00222_),
    .DE(_00095_),
    .Q(\w[11][7] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][8]$_DFFE_PP_  (.D(_00223_),
    .DE(_00095_),
    .Q(\w[11][8] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][9]$_DFFE_PP_  (.D(_00224_),
    .DE(_00095_),
    .Q(\w[11][9] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][0]$_DFFE_PP_  (.D(_00225_),
    .DE(_00125_),
    .Q(\w[12][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][10]$_DFFE_PP_  (.D(_00226_),
    .DE(_00125_),
    .Q(\w[12][10] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][11]$_DFFE_PP_  (.D(_00227_),
    .DE(_00125_),
    .Q(\w[12][11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][12]$_DFFE_PP_  (.D(_00228_),
    .DE(_00125_),
    .Q(\w[12][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][13]$_DFFE_PP_  (.D(_00229_),
    .DE(_00125_),
    .Q(\w[12][13] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][14]$_DFFE_PP_  (.D(_00230_),
    .DE(_00125_),
    .Q(\w[12][14] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][15]$_DFFE_PP_  (.D(_00231_),
    .DE(_00125_),
    .Q(\w[12][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][16]$_DFFE_PP_  (.D(_00232_),
    .DE(_00125_),
    .Q(\w[12][16] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][17]$_DFFE_PP_  (.D(_00233_),
    .DE(_00125_),
    .Q(\w[12][17] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][18]$_DFFE_PP_  (.D(_00234_),
    .DE(_00125_),
    .Q(\w[12][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][19]$_DFFE_PP_  (.D(_00235_),
    .DE(_00125_),
    .Q(\w[12][19] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][1]$_DFFE_PP_  (.D(_00236_),
    .DE(_00125_),
    .Q(\w[12][1] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][20]$_DFFE_PP_  (.D(_00237_),
    .DE(_00125_),
    .Q(\w[12][20] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][21]$_DFFE_PP_  (.D(_00238_),
    .DE(_00125_),
    .Q(\w[12][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][22]$_DFFE_PP_  (.D(_00239_),
    .DE(_00125_),
    .Q(\w[12][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][23]$_DFFE_PP_  (.D(_00240_),
    .DE(_00125_),
    .Q(\w[12][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][24]$_DFFE_PP_  (.D(_00241_),
    .DE(_00125_),
    .Q(\w[12][24] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][25]$_DFFE_PP_  (.D(_00242_),
    .DE(_00125_),
    .Q(\w[12][25] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][26]$_DFFE_PP_  (.D(_00243_),
    .DE(_00125_),
    .Q(\w[12][26] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][27]$_DFFE_PP_  (.D(_00244_),
    .DE(_00125_),
    .Q(\w[12][27] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][28]$_DFFE_PP_  (.D(_00245_),
    .DE(_00125_),
    .Q(\w[12][28] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][29]$_DFFE_PP_  (.D(_00246_),
    .DE(_00125_),
    .Q(\w[12][29] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][2]$_DFFE_PP_  (.D(_00247_),
    .DE(_00125_),
    .Q(\w[12][2] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][30]$_DFFE_PP_  (.D(_00248_),
    .DE(_00125_),
    .Q(\w[12][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][31]$_DFFE_PP_  (.D(_00249_),
    .DE(_00125_),
    .Q(\w[12][31] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][3]$_DFFE_PP_  (.D(_00250_),
    .DE(_00125_),
    .Q(\w[12][3] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][4]$_DFFE_PP_  (.D(_00251_),
    .DE(_00125_),
    .Q(\w[12][4] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][5]$_DFFE_PP_  (.D(_00252_),
    .DE(_00125_),
    .Q(\w[12][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][6]$_DFFE_PP_  (.D(_00253_),
    .DE(_00125_),
    .Q(\w[12][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][7]$_DFFE_PP_  (.D(_00254_),
    .DE(_00125_),
    .Q(\w[12][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][8]$_DFFE_PP_  (.D(_00255_),
    .DE(_00125_),
    .Q(\w[12][8] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][9]$_DFFE_PP_  (.D(_00256_),
    .DE(_00125_),
    .Q(\w[12][9] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][0]$_DFFE_PP_  (.D(_00257_),
    .DE(_00094_),
    .Q(\w[13][0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][10]$_DFFE_PP_  (.D(_00258_),
    .DE(_00094_),
    .Q(\w[13][10] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][11]$_DFFE_PP_  (.D(_00259_),
    .DE(_00094_),
    .Q(\w[13][11] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][12]$_DFFE_PP_  (.D(_00260_),
    .DE(_00094_),
    .Q(\w[13][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][13]$_DFFE_PP_  (.D(_00261_),
    .DE(_00094_),
    .Q(\w[13][13] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][14]$_DFFE_PP_  (.D(_00262_),
    .DE(_00094_),
    .Q(\w[13][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][15]$_DFFE_PP_  (.D(_00263_),
    .DE(_00094_),
    .Q(\w[13][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][16]$_DFFE_PP_  (.D(_00264_),
    .DE(_00094_),
    .Q(\w[13][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][17]$_DFFE_PP_  (.D(_00265_),
    .DE(_00094_),
    .Q(\w[13][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][18]$_DFFE_PP_  (.D(_00266_),
    .DE(_00094_),
    .Q(\w[13][18] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][19]$_DFFE_PP_  (.D(_00267_),
    .DE(_00094_),
    .Q(\w[13][19] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][1]$_DFFE_PP_  (.D(_00268_),
    .DE(_00094_),
    .Q(\w[13][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][20]$_DFFE_PP_  (.D(_00269_),
    .DE(_00094_),
    .Q(\w[13][20] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][21]$_DFFE_PP_  (.D(_00270_),
    .DE(_00094_),
    .Q(\w[13][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][22]$_DFFE_PP_  (.D(_00271_),
    .DE(_00094_),
    .Q(\w[13][22] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][23]$_DFFE_PP_  (.D(_00272_),
    .DE(_00094_),
    .Q(\w[13][23] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][24]$_DFFE_PP_  (.D(_00273_),
    .DE(_00094_),
    .Q(\w[13][24] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][25]$_DFFE_PP_  (.D(_00274_),
    .DE(_00094_),
    .Q(\w[13][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][26]$_DFFE_PP_  (.D(_00275_),
    .DE(_00094_),
    .Q(\w[13][26] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][27]$_DFFE_PP_  (.D(_00276_),
    .DE(_00094_),
    .Q(\w[13][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][28]$_DFFE_PP_  (.D(_00277_),
    .DE(_00094_),
    .Q(\w[13][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][29]$_DFFE_PP_  (.D(_00278_),
    .DE(_00094_),
    .Q(\w[13][29] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][2]$_DFFE_PP_  (.D(_00279_),
    .DE(_00094_),
    .Q(\w[13][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][30]$_DFFE_PP_  (.D(_00280_),
    .DE(_00094_),
    .Q(\w[13][30] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][31]$_DFFE_PP_  (.D(_00281_),
    .DE(_00094_),
    .Q(\w[13][31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][3]$_DFFE_PP_  (.D(_00282_),
    .DE(_00094_),
    .Q(\w[13][3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][4]$_DFFE_PP_  (.D(_00283_),
    .DE(_00094_),
    .Q(\w[13][4] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][5]$_DFFE_PP_  (.D(_00284_),
    .DE(_00094_),
    .Q(\w[13][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][6]$_DFFE_PP_  (.D(_00285_),
    .DE(_00094_),
    .Q(\w[13][6] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][7]$_DFFE_PP_  (.D(_00286_),
    .DE(_00094_),
    .Q(\w[13][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][8]$_DFFE_PP_  (.D(_00287_),
    .DE(_00094_),
    .Q(\w[13][8] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][9]$_DFFE_PP_  (.D(_00288_),
    .DE(_00094_),
    .Q(\w[13][9] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][0]$_DFFE_PP_  (.D(_00289_),
    .DE(_00124_),
    .Q(\w[14][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][10]$_DFFE_PP_  (.D(_00290_),
    .DE(_00124_),
    .Q(\w[14][10] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][11]$_DFFE_PP_  (.D(_00291_),
    .DE(_00124_),
    .Q(\w[14][11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][12]$_DFFE_PP_  (.D(_00292_),
    .DE(_00124_),
    .Q(\w[14][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][13]$_DFFE_PP_  (.D(_00293_),
    .DE(_00124_),
    .Q(\w[14][13] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][14]$_DFFE_PP_  (.D(_00294_),
    .DE(_00124_),
    .Q(\w[14][14] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][15]$_DFFE_PP_  (.D(_00295_),
    .DE(_00124_),
    .Q(\w[14][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][16]$_DFFE_PP_  (.D(_00296_),
    .DE(_00124_),
    .Q(\w[14][16] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][17]$_DFFE_PP_  (.D(_00297_),
    .DE(_00124_),
    .Q(\w[14][17] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][18]$_DFFE_PP_  (.D(_00298_),
    .DE(_00124_),
    .Q(\w[14][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][19]$_DFFE_PP_  (.D(_00299_),
    .DE(_00124_),
    .Q(\w[14][19] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][1]$_DFFE_PP_  (.D(_00300_),
    .DE(_00124_),
    .Q(\w[14][1] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][20]$_DFFE_PP_  (.D(_00301_),
    .DE(_00124_),
    .Q(\w[14][20] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][21]$_DFFE_PP_  (.D(_00302_),
    .DE(_00124_),
    .Q(\w[14][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][22]$_DFFE_PP_  (.D(_00303_),
    .DE(_00124_),
    .Q(\w[14][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][23]$_DFFE_PP_  (.D(_00304_),
    .DE(_00124_),
    .Q(\w[14][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][24]$_DFFE_PP_  (.D(_00305_),
    .DE(_00124_),
    .Q(\w[14][24] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][25]$_DFFE_PP_  (.D(_00306_),
    .DE(_00124_),
    .Q(\w[14][25] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][26]$_DFFE_PP_  (.D(_00307_),
    .DE(_00124_),
    .Q(\w[14][26] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][27]$_DFFE_PP_  (.D(_00308_),
    .DE(_00124_),
    .Q(\w[14][27] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][28]$_DFFE_PP_  (.D(_00309_),
    .DE(_00124_),
    .Q(\w[14][28] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][29]$_DFFE_PP_  (.D(_00310_),
    .DE(_00124_),
    .Q(\w[14][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][2]$_DFFE_PP_  (.D(_00311_),
    .DE(_00124_),
    .Q(\w[14][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][30]$_DFFE_PP_  (.D(_00312_),
    .DE(_00124_),
    .Q(\w[14][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][31]$_DFFE_PP_  (.D(_00313_),
    .DE(_00124_),
    .Q(\w[14][31] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][3]$_DFFE_PP_  (.D(_00314_),
    .DE(_00124_),
    .Q(\w[14][3] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][4]$_DFFE_PP_  (.D(_00315_),
    .DE(_00124_),
    .Q(\w[14][4] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][5]$_DFFE_PP_  (.D(_00316_),
    .DE(_00124_),
    .Q(\w[14][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][6]$_DFFE_PP_  (.D(_00317_),
    .DE(_00124_),
    .Q(\w[14][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][7]$_DFFE_PP_  (.D(_00318_),
    .DE(_00124_),
    .Q(\w[14][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][8]$_DFFE_PP_  (.D(_00319_),
    .DE(_00124_),
    .Q(\w[14][8] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][9]$_DFFE_PP_  (.D(_00320_),
    .DE(_00124_),
    .Q(\w[14][9] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][0]$_DFFE_PP_  (.D(_00321_),
    .DE(_00093_),
    .Q(\w[15][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][10]$_DFFE_PP_  (.D(_00322_),
    .DE(_00093_),
    .Q(\w[15][10] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][11]$_DFFE_PP_  (.D(_00323_),
    .DE(_00093_),
    .Q(\w[15][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][12]$_DFFE_PP_  (.D(_00324_),
    .DE(_00093_),
    .Q(\w[15][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][13]$_DFFE_PP_  (.D(_00325_),
    .DE(_00093_),
    .Q(\w[15][13] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][14]$_DFFE_PP_  (.D(_00326_),
    .DE(_00093_),
    .Q(\w[15][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][15]$_DFFE_PP_  (.D(_00327_),
    .DE(_00093_),
    .Q(\w[15][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][16]$_DFFE_PP_  (.D(_00328_),
    .DE(_00093_),
    .Q(\w[15][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][17]$_DFFE_PP_  (.D(_00329_),
    .DE(_00093_),
    .Q(\w[15][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][18]$_DFFE_PP_  (.D(_00330_),
    .DE(_00093_),
    .Q(\w[15][18] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][19]$_DFFE_PP_  (.D(_00331_),
    .DE(_00093_),
    .Q(\w[15][19] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][1]$_DFFE_PP_  (.D(_00332_),
    .DE(_00093_),
    .Q(\w[15][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][20]$_DFFE_PP_  (.D(_00333_),
    .DE(_00093_),
    .Q(\w[15][20] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][21]$_DFFE_PP_  (.D(_00334_),
    .DE(_00093_),
    .Q(\w[15][21] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][22]$_DFFE_PP_  (.D(_00335_),
    .DE(_00093_),
    .Q(\w[15][22] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][23]$_DFFE_PP_  (.D(_00336_),
    .DE(_00093_),
    .Q(\w[15][23] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][24]$_DFFE_PP_  (.D(_00337_),
    .DE(_00093_),
    .Q(\w[15][24] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][25]$_DFFE_PP_  (.D(_00338_),
    .DE(_00093_),
    .Q(\w[15][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][26]$_DFFE_PP_  (.D(_00339_),
    .DE(_00093_),
    .Q(\w[15][26] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][27]$_DFFE_PP_  (.D(_00340_),
    .DE(_00093_),
    .Q(\w[15][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][28]$_DFFE_PP_  (.D(_00341_),
    .DE(_00093_),
    .Q(\w[15][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][29]$_DFFE_PP_  (.D(_00342_),
    .DE(_00093_),
    .Q(\w[15][29] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][2]$_DFFE_PP_  (.D(_00343_),
    .DE(_00093_),
    .Q(\w[15][2] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][30]$_DFFE_PP_  (.D(_00344_),
    .DE(_00093_),
    .Q(\w[15][30] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][31]$_DFFE_PP_  (.D(_00345_),
    .DE(_00093_),
    .Q(\w[15][31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][3]$_DFFE_PP_  (.D(_00346_),
    .DE(_00093_),
    .Q(\w[15][3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][4]$_DFFE_PP_  (.D(_00347_),
    .DE(_00093_),
    .Q(\w[15][4] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][5]$_DFFE_PP_  (.D(_00348_),
    .DE(_00093_),
    .Q(\w[15][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][6]$_DFFE_PP_  (.D(_00349_),
    .DE(_00093_),
    .Q(\w[15][6] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][7]$_DFFE_PP_  (.D(_00350_),
    .DE(_00093_),
    .Q(\w[15][7] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][8]$_DFFE_PP_  (.D(_00351_),
    .DE(_00093_),
    .Q(\w[15][8] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][9]$_DFFE_PP_  (.D(_00352_),
    .DE(_00093_),
    .Q(\w[15][9] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][0]$_SDFFCE_PN0P_  (.D(_01034_),
    .DE(_00123_),
    .Q(\w[16][0] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][10]$_SDFFCE_PN0P_  (.D(_01035_),
    .DE(_00123_),
    .Q(\w[16][10] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][11]$_SDFFCE_PN0P_  (.D(_01036_),
    .DE(_00123_),
    .Q(\w[16][11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][12]$_SDFFCE_PN0P_  (.D(_01037_),
    .DE(_00123_),
    .Q(\w[16][12] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][13]$_SDFFCE_PN0P_  (.D(_01038_),
    .DE(_00123_),
    .Q(\w[16][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][14]$_SDFFCE_PN0P_  (.D(_01039_),
    .DE(_00123_),
    .Q(\w[16][14] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][15]$_SDFFCE_PN0P_  (.D(_01040_),
    .DE(_00123_),
    .Q(\w[16][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][16]$_SDFFCE_PN0P_  (.D(_01041_),
    .DE(_00123_),
    .Q(\w[16][16] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][17]$_SDFFCE_PN0P_  (.D(_01042_),
    .DE(_00123_),
    .Q(\w[16][17] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][18]$_SDFFCE_PN0P_  (.D(_01043_),
    .DE(_00123_),
    .Q(\w[16][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][19]$_SDFFCE_PN0P_  (.D(_01044_),
    .DE(_00123_),
    .Q(\w[16][19] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][1]$_SDFFCE_PN0P_  (.D(_01045_),
    .DE(_00123_),
    .Q(\w[16][1] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][20]$_SDFFCE_PN0P_  (.D(_01046_),
    .DE(_00123_),
    .Q(\w[16][20] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][21]$_SDFFCE_PN0P_  (.D(_01047_),
    .DE(_00123_),
    .Q(\w[16][21] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][22]$_SDFFCE_PN0P_  (.D(_01048_),
    .DE(_00123_),
    .Q(\w[16][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][23]$_SDFFCE_PN0P_  (.D(_01049_),
    .DE(_00123_),
    .Q(\w[16][23] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][24]$_SDFFCE_PN0P_  (.D(_01050_),
    .DE(_00123_),
    .Q(\w[16][24] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][25]$_SDFFCE_PN0P_  (.D(_01051_),
    .DE(_00123_),
    .Q(\w[16][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][26]$_SDFFCE_PN0P_  (.D(_01052_),
    .DE(_00123_),
    .Q(\w[16][26] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][27]$_SDFFCE_PN0P_  (.D(_01053_),
    .DE(_00123_),
    .Q(\w[16][27] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][28]$_SDFFCE_PN0P_  (.D(_01054_),
    .DE(_00123_),
    .Q(\w[16][28] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][29]$_SDFFCE_PN0P_  (.D(_01055_),
    .DE(_00123_),
    .Q(\w[16][29] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][2]$_SDFFCE_PN0P_  (.D(_01056_),
    .DE(_00123_),
    .Q(\w[16][2] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][30]$_SDFFCE_PN0P_  (.D(_01057_),
    .DE(_00123_),
    .Q(\w[16][30] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][31]$_SDFFCE_PN0P_  (.D(_01058_),
    .DE(_00123_),
    .Q(\w[16][31] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][3]$_SDFFCE_PN0P_  (.D(_01059_),
    .DE(_00123_),
    .Q(\w[16][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][4]$_SDFFCE_PN0P_  (.D(_01060_),
    .DE(_00123_),
    .Q(\w[16][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][5]$_SDFFCE_PN0P_  (.D(_01061_),
    .DE(_00123_),
    .Q(\w[16][5] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][6]$_SDFFCE_PN0P_  (.D(_01062_),
    .DE(_00123_),
    .Q(\w[16][6] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][7]$_SDFFCE_PN0P_  (.D(_01063_),
    .DE(_00123_),
    .Q(\w[16][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][8]$_SDFFCE_PN0P_  (.D(_01064_),
    .DE(_00123_),
    .Q(\w[16][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][9]$_SDFFCE_PN0P_  (.D(_01065_),
    .DE(_00123_),
    .Q(\w[16][9] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][0]$_SDFFCE_PN0P_  (.D(_01066_),
    .DE(_00092_),
    .Q(\w[17][0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][10]$_SDFFCE_PN0P_  (.D(_01067_),
    .DE(_00092_),
    .Q(\w[17][10] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][11]$_SDFFCE_PN0P_  (.D(_01068_),
    .DE(_00092_),
    .Q(\w[17][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][12]$_SDFFCE_PN0P_  (.D(_01069_),
    .DE(_00092_),
    .Q(\w[17][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][13]$_SDFFCE_PN0P_  (.D(_01070_),
    .DE(_00092_),
    .Q(\w[17][13] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][14]$_SDFFCE_PN0P_  (.D(_01071_),
    .DE(_00092_),
    .Q(\w[17][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][15]$_SDFFCE_PN0P_  (.D(_01072_),
    .DE(_00092_),
    .Q(\w[17][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][16]$_SDFFCE_PN0P_  (.D(_01073_),
    .DE(_00092_),
    .Q(\w[17][16] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][17]$_SDFFCE_PN0P_  (.D(_01074_),
    .DE(_00092_),
    .Q(\w[17][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][18]$_SDFFCE_PN0P_  (.D(_01075_),
    .DE(_00092_),
    .Q(\w[17][18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][19]$_SDFFCE_PN0P_  (.D(_01076_),
    .DE(_00092_),
    .Q(\w[17][19] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][1]$_SDFFCE_PN0P_  (.D(_01077_),
    .DE(_00092_),
    .Q(\w[17][1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][20]$_SDFFCE_PN0P_  (.D(_01078_),
    .DE(_00092_),
    .Q(\w[17][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][21]$_SDFFCE_PN0P_  (.D(_01079_),
    .DE(_00092_),
    .Q(\w[17][21] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][22]$_SDFFCE_PN0P_  (.D(_01080_),
    .DE(_00092_),
    .Q(\w[17][22] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][23]$_SDFFCE_PN0P_  (.D(_01081_),
    .DE(_00092_),
    .Q(\w[17][23] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][24]$_SDFFCE_PN0P_  (.D(_01082_),
    .DE(_00092_),
    .Q(\w[17][24] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][25]$_SDFFCE_PN0P_  (.D(_01083_),
    .DE(_00092_),
    .Q(\w[17][25] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][26]$_SDFFCE_PN0P_  (.D(_01084_),
    .DE(_00092_),
    .Q(\w[17][26] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][27]$_SDFFCE_PN0P_  (.D(_01085_),
    .DE(_00092_),
    .Q(\w[17][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][28]$_SDFFCE_PN0P_  (.D(_01086_),
    .DE(_00092_),
    .Q(\w[17][28] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][29]$_SDFFCE_PN0P_  (.D(_01087_),
    .DE(_00092_),
    .Q(\w[17][29] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][2]$_SDFFCE_PN0P_  (.D(_01088_),
    .DE(_00092_),
    .Q(\w[17][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][30]$_SDFFCE_PN0P_  (.D(_01089_),
    .DE(_00092_),
    .Q(\w[17][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][31]$_SDFFCE_PN0P_  (.D(_01090_),
    .DE(_00092_),
    .Q(\w[17][31] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][3]$_SDFFCE_PN0P_  (.D(_01091_),
    .DE(_00092_),
    .Q(\w[17][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][4]$_SDFFCE_PN0P_  (.D(_01092_),
    .DE(_00092_),
    .Q(\w[17][4] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][5]$_SDFFCE_PN0P_  (.D(_01093_),
    .DE(_00092_),
    .Q(\w[17][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][6]$_SDFFCE_PN0P_  (.D(_01094_),
    .DE(_00092_),
    .Q(\w[17][6] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][7]$_SDFFCE_PN0P_  (.D(_01095_),
    .DE(_00092_),
    .Q(\w[17][7] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][8]$_SDFFCE_PN0P_  (.D(_01096_),
    .DE(_00092_),
    .Q(\w[17][8] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][9]$_SDFFCE_PN0P_  (.D(_01097_),
    .DE(_00092_),
    .Q(\w[17][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][0]$_SDFFCE_PN0P_  (.D(_01098_),
    .DE(_00122_),
    .Q(\w[18][0] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][10]$_SDFFCE_PN0P_  (.D(_01099_),
    .DE(_00122_),
    .Q(\w[18][10] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][11]$_SDFFCE_PN0P_  (.D(_01100_),
    .DE(_00122_),
    .Q(\w[18][11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][12]$_SDFFCE_PN0P_  (.D(_01101_),
    .DE(_00122_),
    .Q(\w[18][12] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][13]$_SDFFCE_PN0P_  (.D(_01102_),
    .DE(_00122_),
    .Q(\w[18][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][14]$_SDFFCE_PN0P_  (.D(_01103_),
    .DE(_00122_),
    .Q(\w[18][14] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][15]$_SDFFCE_PN0P_  (.D(_01104_),
    .DE(_00122_),
    .Q(\w[18][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][16]$_SDFFCE_PN0P_  (.D(_01105_),
    .DE(_00122_),
    .Q(\w[18][16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][17]$_SDFFCE_PN0P_  (.D(_01106_),
    .DE(_00122_),
    .Q(\w[18][17] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][18]$_SDFFCE_PN0P_  (.D(_01107_),
    .DE(_00122_),
    .Q(\w[18][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][19]$_SDFFCE_PN0P_  (.D(_01108_),
    .DE(_00122_),
    .Q(\w[18][19] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][1]$_SDFFCE_PN0P_  (.D(_01109_),
    .DE(_00122_),
    .Q(\w[18][1] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][20]$_SDFFCE_PN0P_  (.D(_01110_),
    .DE(_00122_),
    .Q(\w[18][20] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][21]$_SDFFCE_PN0P_  (.D(_01111_),
    .DE(_00122_),
    .Q(\w[18][21] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][22]$_SDFFCE_PN0P_  (.D(_01112_),
    .DE(_00122_),
    .Q(\w[18][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][23]$_SDFFCE_PN0P_  (.D(_01113_),
    .DE(_00122_),
    .Q(\w[18][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][24]$_SDFFCE_PN0P_  (.D(_01114_),
    .DE(_00122_),
    .Q(\w[18][24] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][25]$_SDFFCE_PN0P_  (.D(_01115_),
    .DE(_00122_),
    .Q(\w[18][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][26]$_SDFFCE_PN0P_  (.D(_01116_),
    .DE(_00122_),
    .Q(\w[18][26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][27]$_SDFFCE_PN0P_  (.D(_01117_),
    .DE(_00122_),
    .Q(\w[18][27] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][28]$_SDFFCE_PN0P_  (.D(_01118_),
    .DE(_00122_),
    .Q(\w[18][28] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][29]$_SDFFCE_PN0P_  (.D(_01119_),
    .DE(_00122_),
    .Q(\w[18][29] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][2]$_SDFFCE_PN0P_  (.D(_01120_),
    .DE(_00122_),
    .Q(\w[18][2] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][30]$_SDFFCE_PN0P_  (.D(_01121_),
    .DE(_00122_),
    .Q(\w[18][30] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][31]$_SDFFCE_PN0P_  (.D(_01122_),
    .DE(_00122_),
    .Q(\w[18][31] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][3]$_SDFFCE_PN0P_  (.D(_01123_),
    .DE(_00122_),
    .Q(\w[18][3] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][4]$_SDFFCE_PN0P_  (.D(_01124_),
    .DE(_00122_),
    .Q(\w[18][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][5]$_SDFFCE_PN0P_  (.D(_01125_),
    .DE(_00122_),
    .Q(\w[18][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][6]$_SDFFCE_PN0P_  (.D(_01126_),
    .DE(_00122_),
    .Q(\w[18][6] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][7]$_SDFFCE_PN0P_  (.D(_01127_),
    .DE(_00122_),
    .Q(\w[18][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][8]$_SDFFCE_PN0P_  (.D(_01128_),
    .DE(_00122_),
    .Q(\w[18][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][9]$_SDFFCE_PN0P_  (.D(_01129_),
    .DE(_00122_),
    .Q(\w[18][9] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][0]$_SDFFCE_PN0P_  (.D(_01130_),
    .DE(_00091_),
    .Q(\w[19][0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][10]$_SDFFCE_PN0P_  (.D(_01131_),
    .DE(_00091_),
    .Q(\w[19][10] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][11]$_SDFFCE_PN0P_  (.D(_01132_),
    .DE(_00091_),
    .Q(\w[19][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][12]$_SDFFCE_PN0P_  (.D(_01133_),
    .DE(_00091_),
    .Q(\w[19][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][13]$_SDFFCE_PN0P_  (.D(_01134_),
    .DE(_00091_),
    .Q(\w[19][13] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][14]$_SDFFCE_PN0P_  (.D(_01135_),
    .DE(_00091_),
    .Q(\w[19][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][15]$_SDFFCE_PN0P_  (.D(_01136_),
    .DE(_00091_),
    .Q(\w[19][15] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][16]$_SDFFCE_PN0P_  (.D(_01137_),
    .DE(_00091_),
    .Q(\w[19][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][17]$_SDFFCE_PN0P_  (.D(_01138_),
    .DE(_00091_),
    .Q(\w[19][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][18]$_SDFFCE_PN0P_  (.D(_01139_),
    .DE(_00091_),
    .Q(\w[19][18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][19]$_SDFFCE_PN0P_  (.D(_01140_),
    .DE(_00091_),
    .Q(\w[19][19] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][1]$_SDFFCE_PN0P_  (.D(_01141_),
    .DE(_00091_),
    .Q(\w[19][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][20]$_SDFFCE_PN0P_  (.D(_01142_),
    .DE(_00091_),
    .Q(\w[19][20] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][21]$_SDFFCE_PN0P_  (.D(_01143_),
    .DE(_00091_),
    .Q(\w[19][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][22]$_SDFFCE_PN0P_  (.D(_01144_),
    .DE(_00091_),
    .Q(\w[19][22] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][23]$_SDFFCE_PN0P_  (.D(_01145_),
    .DE(_00091_),
    .Q(\w[19][23] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][24]$_SDFFCE_PN0P_  (.D(_01146_),
    .DE(_00091_),
    .Q(\w[19][24] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][25]$_SDFFCE_PN0P_  (.D(_01147_),
    .DE(_00091_),
    .Q(\w[19][25] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][26]$_SDFFCE_PN0P_  (.D(_01148_),
    .DE(_00091_),
    .Q(\w[19][26] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][27]$_SDFFCE_PN0P_  (.D(_01149_),
    .DE(_00091_),
    .Q(\w[19][27] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][28]$_SDFFCE_PN0P_  (.D(_01150_),
    .DE(_00091_),
    .Q(\w[19][28] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][29]$_SDFFCE_PN0P_  (.D(_01151_),
    .DE(_00091_),
    .Q(\w[19][29] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][2]$_SDFFCE_PN0P_  (.D(_01152_),
    .DE(_00091_),
    .Q(\w[19][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][30]$_SDFFCE_PN0P_  (.D(_01153_),
    .DE(_00091_),
    .Q(\w[19][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][31]$_SDFFCE_PN0P_  (.D(_01154_),
    .DE(_00091_),
    .Q(\w[19][31] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][3]$_SDFFCE_PN0P_  (.D(_01155_),
    .DE(_00091_),
    .Q(\w[19][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][4]$_SDFFCE_PN0P_  (.D(_01156_),
    .DE(_00091_),
    .Q(\w[19][4] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][5]$_SDFFCE_PN0P_  (.D(_01157_),
    .DE(_00091_),
    .Q(\w[19][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][6]$_SDFFCE_PN0P_  (.D(_01158_),
    .DE(_00091_),
    .Q(\w[19][6] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][7]$_SDFFCE_PN0P_  (.D(_01159_),
    .DE(_00091_),
    .Q(\w[19][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][8]$_SDFFCE_PN0P_  (.D(_01160_),
    .DE(_00091_),
    .Q(\w[19][8] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][9]$_SDFFCE_PN0P_  (.D(_01161_),
    .DE(_00091_),
    .Q(\w[19][9] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][0]$_DFFE_PP_  (.D(_00353_),
    .DE(_00090_),
    .Q(\w[1][0] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][10]$_DFFE_PP_  (.D(_00354_),
    .DE(_00090_),
    .Q(\w[1][10] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][11]$_DFFE_PP_  (.D(_00355_),
    .DE(_00090_),
    .Q(\w[1][11] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][12]$_DFFE_PP_  (.D(_00356_),
    .DE(_00090_),
    .Q(\w[1][12] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][13]$_DFFE_PP_  (.D(_00357_),
    .DE(_00090_),
    .Q(\w[1][13] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][14]$_DFFE_PP_  (.D(_00358_),
    .DE(_00090_),
    .Q(\w[1][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][15]$_DFFE_PP_  (.D(_00359_),
    .DE(_00090_),
    .Q(\w[1][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][16]$_DFFE_PP_  (.D(_00360_),
    .DE(_00090_),
    .Q(\w[1][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][17]$_DFFE_PP_  (.D(_00361_),
    .DE(_00090_),
    .Q(\w[1][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][18]$_DFFE_PP_  (.D(_00362_),
    .DE(_00090_),
    .Q(\w[1][18] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][19]$_DFFE_PP_  (.D(_00363_),
    .DE(_00090_),
    .Q(\w[1][19] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][1]$_DFFE_PP_  (.D(_00364_),
    .DE(_00090_),
    .Q(\w[1][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][20]$_DFFE_PP_  (.D(_00365_),
    .DE(_00090_),
    .Q(\w[1][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][21]$_DFFE_PP_  (.D(_00366_),
    .DE(_00090_),
    .Q(\w[1][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][22]$_DFFE_PP_  (.D(_00367_),
    .DE(_00090_),
    .Q(\w[1][22] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][23]$_DFFE_PP_  (.D(_00368_),
    .DE(_00090_),
    .Q(\w[1][23] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][24]$_DFFE_PP_  (.D(_00369_),
    .DE(_00090_),
    .Q(\w[1][24] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][25]$_DFFE_PP_  (.D(_00370_),
    .DE(_00090_),
    .Q(\w[1][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][26]$_DFFE_PP_  (.D(_00371_),
    .DE(_00090_),
    .Q(\w[1][26] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][27]$_DFFE_PP_  (.D(_00372_),
    .DE(_00090_),
    .Q(\w[1][27] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][28]$_DFFE_PP_  (.D(_00373_),
    .DE(_00090_),
    .Q(\w[1][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][29]$_DFFE_PP_  (.D(_00374_),
    .DE(_00090_),
    .Q(\w[1][29] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][2]$_DFFE_PP_  (.D(_00375_),
    .DE(_00090_),
    .Q(\w[1][2] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][30]$_DFFE_PP_  (.D(_00376_),
    .DE(_00090_),
    .Q(\w[1][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][31]$_DFFE_PP_  (.D(_00377_),
    .DE(_00090_),
    .Q(\w[1][31] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][3]$_DFFE_PP_  (.D(_00378_),
    .DE(_00090_),
    .Q(\w[1][3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][4]$_DFFE_PP_  (.D(_00379_),
    .DE(_00090_),
    .Q(\w[1][4] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][5]$_DFFE_PP_  (.D(_00380_),
    .DE(_00090_),
    .Q(\w[1][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][6]$_DFFE_PP_  (.D(_00381_),
    .DE(_00090_),
    .Q(\w[1][6] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][7]$_DFFE_PP_  (.D(_00382_),
    .DE(_00090_),
    .Q(\w[1][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][8]$_DFFE_PP_  (.D(_00383_),
    .DE(_00090_),
    .Q(\w[1][8] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][9]$_DFFE_PP_  (.D(_00384_),
    .DE(_00090_),
    .Q(\w[1][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][0]$_SDFFCE_PN0P_  (.D(_01162_),
    .DE(_00121_),
    .Q(\w[20][0] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][10]$_SDFFCE_PN0P_  (.D(_01163_),
    .DE(_00121_),
    .Q(\w[20][10] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][11]$_SDFFCE_PN0P_  (.D(_01164_),
    .DE(_00121_),
    .Q(\w[20][11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][12]$_SDFFCE_PN0P_  (.D(_01165_),
    .DE(_00121_),
    .Q(\w[20][12] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][13]$_SDFFCE_PN0P_  (.D(_01166_),
    .DE(_00121_),
    .Q(\w[20][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][14]$_SDFFCE_PN0P_  (.D(_01167_),
    .DE(_00121_),
    .Q(\w[20][14] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][15]$_SDFFCE_PN0P_  (.D(_01168_),
    .DE(_00121_),
    .Q(\w[20][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][16]$_SDFFCE_PN0P_  (.D(_01169_),
    .DE(_00121_),
    .Q(\w[20][16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][17]$_SDFFCE_PN0P_  (.D(_01170_),
    .DE(_00121_),
    .Q(\w[20][17] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][18]$_SDFFCE_PN0P_  (.D(_01171_),
    .DE(_00121_),
    .Q(\w[20][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][19]$_SDFFCE_PN0P_  (.D(_01172_),
    .DE(_00121_),
    .Q(\w[20][19] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][1]$_SDFFCE_PN0P_  (.D(_01173_),
    .DE(_00121_),
    .Q(\w[20][1] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][20]$_SDFFCE_PN0P_  (.D(_01174_),
    .DE(_00121_),
    .Q(\w[20][20] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][21]$_SDFFCE_PN0P_  (.D(_01175_),
    .DE(_00121_),
    .Q(\w[20][21] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][22]$_SDFFCE_PN0P_  (.D(_01176_),
    .DE(_00121_),
    .Q(\w[20][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][23]$_SDFFCE_PN0P_  (.D(_01177_),
    .DE(_00121_),
    .Q(\w[20][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][24]$_SDFFCE_PN0P_  (.D(_01178_),
    .DE(_00121_),
    .Q(\w[20][24] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][25]$_SDFFCE_PN0P_  (.D(_01179_),
    .DE(_00121_),
    .Q(\w[20][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][26]$_SDFFCE_PN0P_  (.D(_01180_),
    .DE(_00121_),
    .Q(\w[20][26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][27]$_SDFFCE_PN0P_  (.D(_01181_),
    .DE(_00121_),
    .Q(\w[20][27] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][28]$_SDFFCE_PN0P_  (.D(_01182_),
    .DE(_00121_),
    .Q(\w[20][28] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][29]$_SDFFCE_PN0P_  (.D(_01183_),
    .DE(_00121_),
    .Q(\w[20][29] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][2]$_SDFFCE_PN0P_  (.D(_01184_),
    .DE(_00121_),
    .Q(\w[20][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][30]$_SDFFCE_PN0P_  (.D(_01185_),
    .DE(_00121_),
    .Q(\w[20][30] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][31]$_SDFFCE_PN0P_  (.D(_01186_),
    .DE(_00121_),
    .Q(\w[20][31] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][3]$_SDFFCE_PN0P_  (.D(_01187_),
    .DE(_00121_),
    .Q(\w[20][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][4]$_SDFFCE_PN0P_  (.D(_01188_),
    .DE(_00121_),
    .Q(\w[20][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][5]$_SDFFCE_PN0P_  (.D(_01189_),
    .DE(_00121_),
    .Q(\w[20][5] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][6]$_SDFFCE_PN0P_  (.D(_01190_),
    .DE(_00121_),
    .Q(\w[20][6] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][7]$_SDFFCE_PN0P_  (.D(_01191_),
    .DE(_00121_),
    .Q(\w[20][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][8]$_SDFFCE_PN0P_  (.D(_01192_),
    .DE(_00121_),
    .Q(\w[20][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][9]$_SDFFCE_PN0P_  (.D(_01193_),
    .DE(_00121_),
    .Q(\w[20][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][0]$_SDFFCE_PN0P_  (.D(_01194_),
    .DE(_00089_),
    .Q(\w[21][0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][10]$_SDFFCE_PN0P_  (.D(_01195_),
    .DE(_00089_),
    .Q(\w[21][10] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][11]$_SDFFCE_PN0P_  (.D(_01196_),
    .DE(_00089_),
    .Q(\w[21][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][12]$_SDFFCE_PN0P_  (.D(_01197_),
    .DE(_00089_),
    .Q(\w[21][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][13]$_SDFFCE_PN0P_  (.D(_01198_),
    .DE(_00089_),
    .Q(\w[21][13] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][14]$_SDFFCE_PN0P_  (.D(_01199_),
    .DE(_00089_),
    .Q(\w[21][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][15]$_SDFFCE_PN0P_  (.D(_01200_),
    .DE(_00089_),
    .Q(\w[21][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][16]$_SDFFCE_PN0P_  (.D(_01201_),
    .DE(_00089_),
    .Q(\w[21][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][17]$_SDFFCE_PN0P_  (.D(_01202_),
    .DE(_00089_),
    .Q(\w[21][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][18]$_SDFFCE_PN0P_  (.D(_01203_),
    .DE(_00089_),
    .Q(\w[21][18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][19]$_SDFFCE_PN0P_  (.D(_01204_),
    .DE(_00089_),
    .Q(\w[21][19] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][1]$_SDFFCE_PN0P_  (.D(_01205_),
    .DE(_00089_),
    .Q(\w[21][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][20]$_SDFFCE_PN0P_  (.D(_01206_),
    .DE(_00089_),
    .Q(\w[21][20] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][21]$_SDFFCE_PN0P_  (.D(_01207_),
    .DE(_00089_),
    .Q(\w[21][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][22]$_SDFFCE_PN0P_  (.D(_01208_),
    .DE(_00089_),
    .Q(\w[21][22] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][23]$_SDFFCE_PN0P_  (.D(_01209_),
    .DE(_00089_),
    .Q(\w[21][23] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][24]$_SDFFCE_PN0P_  (.D(_01210_),
    .DE(_00089_),
    .Q(\w[21][24] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][25]$_SDFFCE_PN0P_  (.D(_01211_),
    .DE(_00089_),
    .Q(\w[21][25] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][26]$_SDFFCE_PN0P_  (.D(_01212_),
    .DE(_00089_),
    .Q(\w[21][26] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][27]$_SDFFCE_PN0P_  (.D(_01213_),
    .DE(_00089_),
    .Q(\w[21][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][28]$_SDFFCE_PN0P_  (.D(_01214_),
    .DE(_00089_),
    .Q(\w[21][28] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][29]$_SDFFCE_PN0P_  (.D(_01215_),
    .DE(_00089_),
    .Q(\w[21][29] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][2]$_SDFFCE_PN0P_  (.D(_01216_),
    .DE(_00089_),
    .Q(\w[21][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][30]$_SDFFCE_PN0P_  (.D(_01217_),
    .DE(_00089_),
    .Q(\w[21][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][31]$_SDFFCE_PN0P_  (.D(_01218_),
    .DE(_00089_),
    .Q(\w[21][31] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][3]$_SDFFCE_PN0P_  (.D(_01219_),
    .DE(_00089_),
    .Q(\w[21][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][4]$_SDFFCE_PN0P_  (.D(_01220_),
    .DE(_00089_),
    .Q(\w[21][4] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][5]$_SDFFCE_PN0P_  (.D(_01221_),
    .DE(_00089_),
    .Q(\w[21][5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][6]$_SDFFCE_PN0P_  (.D(_01222_),
    .DE(_00089_),
    .Q(\w[21][6] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][7]$_SDFFCE_PN0P_  (.D(_01223_),
    .DE(_00089_),
    .Q(\w[21][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][8]$_SDFFCE_PN0P_  (.D(_01224_),
    .DE(_00089_),
    .Q(\w[21][8] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][9]$_SDFFCE_PN0P_  (.D(_01225_),
    .DE(_00089_),
    .Q(\w[21][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][0]$_SDFFCE_PN0P_  (.D(_01226_),
    .DE(_00120_),
    .Q(\w[22][0] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][10]$_SDFFCE_PN0P_  (.D(_01227_),
    .DE(_00120_),
    .Q(\w[22][10] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][11]$_SDFFCE_PN0P_  (.D(_01228_),
    .DE(_00120_),
    .Q(\w[22][11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][12]$_SDFFCE_PN0P_  (.D(_01229_),
    .DE(_00120_),
    .Q(\w[22][12] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][13]$_SDFFCE_PN0P_  (.D(_01230_),
    .DE(_00120_),
    .Q(\w[22][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][14]$_SDFFCE_PN0P_  (.D(_01231_),
    .DE(_00120_),
    .Q(\w[22][14] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][15]$_SDFFCE_PN0P_  (.D(_01232_),
    .DE(_00120_),
    .Q(\w[22][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][16]$_SDFFCE_PN0P_  (.D(_01233_),
    .DE(_00120_),
    .Q(\w[22][16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][17]$_SDFFCE_PN0P_  (.D(_01234_),
    .DE(_00120_),
    .Q(\w[22][17] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][18]$_SDFFCE_PN0P_  (.D(_01235_),
    .DE(_00120_),
    .Q(\w[22][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][19]$_SDFFCE_PN0P_  (.D(_01236_),
    .DE(_00120_),
    .Q(\w[22][19] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][1]$_SDFFCE_PN0P_  (.D(_01237_),
    .DE(_00120_),
    .Q(\w[22][1] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][20]$_SDFFCE_PN0P_  (.D(_01238_),
    .DE(_00120_),
    .Q(\w[22][20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][21]$_SDFFCE_PN0P_  (.D(_01239_),
    .DE(_00120_),
    .Q(\w[22][21] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][22]$_SDFFCE_PN0P_  (.D(_01240_),
    .DE(_00120_),
    .Q(\w[22][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][23]$_SDFFCE_PN0P_  (.D(_01241_),
    .DE(_00120_),
    .Q(\w[22][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][24]$_SDFFCE_PN0P_  (.D(_01242_),
    .DE(_00120_),
    .Q(\w[22][24] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][25]$_SDFFCE_PN0P_  (.D(_01243_),
    .DE(_00120_),
    .Q(\w[22][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][26]$_SDFFCE_PN0P_  (.D(_01244_),
    .DE(_00120_),
    .Q(\w[22][26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][27]$_SDFFCE_PN0P_  (.D(_01245_),
    .DE(_00120_),
    .Q(\w[22][27] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][28]$_SDFFCE_PN0P_  (.D(_01246_),
    .DE(_00120_),
    .Q(\w[22][28] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][29]$_SDFFCE_PN0P_  (.D(_01247_),
    .DE(_00120_),
    .Q(\w[22][29] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][2]$_SDFFCE_PN0P_  (.D(_01248_),
    .DE(_00120_),
    .Q(\w[22][2] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][30]$_SDFFCE_PN0P_  (.D(_01249_),
    .DE(_00120_),
    .Q(\w[22][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][31]$_SDFFCE_PN0P_  (.D(_01250_),
    .DE(_00120_),
    .Q(\w[22][31] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][3]$_SDFFCE_PN0P_  (.D(_01251_),
    .DE(_00120_),
    .Q(\w[22][3] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][4]$_SDFFCE_PN0P_  (.D(_01252_),
    .DE(_00120_),
    .Q(\w[22][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][5]$_SDFFCE_PN0P_  (.D(_01253_),
    .DE(_00120_),
    .Q(\w[22][5] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][6]$_SDFFCE_PN0P_  (.D(_01254_),
    .DE(_00120_),
    .Q(\w[22][6] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][7]$_SDFFCE_PN0P_  (.D(_01255_),
    .DE(_00120_),
    .Q(\w[22][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][8]$_SDFFCE_PN0P_  (.D(_01256_),
    .DE(_00120_),
    .Q(\w[22][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][9]$_SDFFCE_PN0P_  (.D(_01257_),
    .DE(_00120_),
    .Q(\w[22][9] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][0]$_SDFFCE_PN0P_  (.D(_01258_),
    .DE(net475),
    .Q(\w[23][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][10]$_SDFFCE_PN0P_  (.D(_01259_),
    .DE(net476),
    .Q(\w[23][10] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][11]$_SDFFCE_PN0P_  (.D(_01260_),
    .DE(net476),
    .Q(\w[23][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][12]$_SDFFCE_PN0P_  (.D(_01261_),
    .DE(net475),
    .Q(\w[23][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][13]$_SDFFCE_PN0P_  (.D(_01262_),
    .DE(net476),
    .Q(\w[23][13] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][14]$_SDFFCE_PN0P_  (.D(_01263_),
    .DE(net475),
    .Q(\w[23][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][15]$_SDFFCE_PN0P_  (.D(_01264_),
    .DE(net475),
    .Q(\w[23][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][16]$_SDFFCE_PN0P_  (.D(_01265_),
    .DE(net475),
    .Q(\w[23][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][17]$_SDFFCE_PN0P_  (.D(_01266_),
    .DE(net475),
    .Q(\w[23][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][18]$_SDFFCE_PN0P_  (.D(_01267_),
    .DE(net476),
    .Q(\w[23][18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][19]$_SDFFCE_PN0P_  (.D(_01268_),
    .DE(net476),
    .Q(\w[23][19] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][1]$_SDFFCE_PN0P_  (.D(_01269_),
    .DE(net475),
    .Q(\w[23][1] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][20]$_SDFFCE_PN0P_  (.D(_01270_),
    .DE(net476),
    .Q(\w[23][20] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][21]$_SDFFCE_PN0P_  (.D(_01271_),
    .DE(net476),
    .Q(\w[23][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][22]$_SDFFCE_PN0P_  (.D(_01272_),
    .DE(net476),
    .Q(\w[23][22] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][23]$_SDFFCE_PN0P_  (.D(_01273_),
    .DE(net475),
    .Q(\w[23][23] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][24]$_SDFFCE_PN0P_  (.D(_01274_),
    .DE(net475),
    .Q(\w[23][24] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][25]$_SDFFCE_PN0P_  (.D(_01275_),
    .DE(net475),
    .Q(\w[23][25] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][26]$_SDFFCE_PN0P_  (.D(_01276_),
    .DE(net475),
    .Q(\w[23][26] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][27]$_SDFFCE_PN0P_  (.D(_01277_),
    .DE(net475),
    .Q(\w[23][27] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][28]$_SDFFCE_PN0P_  (.D(_01278_),
    .DE(net476),
    .Q(\w[23][28] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][29]$_SDFFCE_PN0P_  (.D(_01279_),
    .DE(net476),
    .Q(\w[23][29] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][2]$_SDFFCE_PN0P_  (.D(_01280_),
    .DE(net475),
    .Q(\w[23][2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][30]$_SDFFCE_PN0P_  (.D(_01281_),
    .DE(net476),
    .Q(\w[23][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][31]$_SDFFCE_PN0P_  (.D(_01282_),
    .DE(net476),
    .Q(\w[23][31] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][3]$_SDFFCE_PN0P_  (.D(_01283_),
    .DE(net475),
    .Q(\w[23][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][4]$_SDFFCE_PN0P_  (.D(_01284_),
    .DE(_00088_),
    .Q(\w[23][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][5]$_SDFFCE_PN0P_  (.D(_01285_),
    .DE(net475),
    .Q(\w[23][5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][6]$_SDFFCE_PN0P_  (.D(_01286_),
    .DE(net476),
    .Q(\w[23][6] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][7]$_SDFFCE_PN0P_  (.D(_01287_),
    .DE(net475),
    .Q(\w[23][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][8]$_SDFFCE_PN0P_  (.D(_01288_),
    .DE(net475),
    .Q(\w[23][8] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][9]$_SDFFCE_PN0P_  (.D(_01289_),
    .DE(net476),
    .Q(\w[23][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][0]$_SDFFCE_PN0P_  (.D(_01290_),
    .DE(_00119_),
    .Q(\w[24][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][10]$_SDFFCE_PN0P_  (.D(_01291_),
    .DE(_00119_),
    .Q(\w[24][10] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][11]$_SDFFCE_PN0P_  (.D(_01292_),
    .DE(_00119_),
    .Q(\w[24][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][12]$_SDFFCE_PN0P_  (.D(_01293_),
    .DE(_00119_),
    .Q(\w[24][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][13]$_SDFFCE_PN0P_  (.D(_01294_),
    .DE(_00119_),
    .Q(\w[24][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][14]$_SDFFCE_PN0P_  (.D(_01295_),
    .DE(_00119_),
    .Q(\w[24][14] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][15]$_SDFFCE_PN0P_  (.D(_01296_),
    .DE(_00119_),
    .Q(\w[24][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][16]$_SDFFCE_PN0P_  (.D(_01297_),
    .DE(_00119_),
    .Q(\w[24][16] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][17]$_SDFFCE_PN0P_  (.D(_01298_),
    .DE(_00119_),
    .Q(\w[24][17] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][18]$_SDFFCE_PN0P_  (.D(_01299_),
    .DE(_00119_),
    .Q(\w[24][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][19]$_SDFFCE_PN0P_  (.D(_01300_),
    .DE(_00119_),
    .Q(\w[24][19] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][1]$_SDFFCE_PN0P_  (.D(_01301_),
    .DE(_00119_),
    .Q(\w[24][1] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][20]$_SDFFCE_PN0P_  (.D(_01302_),
    .DE(_00119_),
    .Q(\w[24][20] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][21]$_SDFFCE_PN0P_  (.D(_01303_),
    .DE(_00119_),
    .Q(\w[24][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][22]$_SDFFCE_PN0P_  (.D(_01304_),
    .DE(_00119_),
    .Q(\w[24][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][23]$_SDFFCE_PN0P_  (.D(_01305_),
    .DE(_00119_),
    .Q(\w[24][23] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][24]$_SDFFCE_PN0P_  (.D(_01306_),
    .DE(_00119_),
    .Q(\w[24][24] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][25]$_SDFFCE_PN0P_  (.D(_01307_),
    .DE(_00119_),
    .Q(\w[24][25] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][26]$_SDFFCE_PN0P_  (.D(_01308_),
    .DE(_00119_),
    .Q(\w[24][26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][27]$_SDFFCE_PN0P_  (.D(_01309_),
    .DE(_00119_),
    .Q(\w[24][27] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][28]$_SDFFCE_PN0P_  (.D(_01310_),
    .DE(_00119_),
    .Q(\w[24][28] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][29]$_SDFFCE_PN0P_  (.D(_01311_),
    .DE(_00119_),
    .Q(\w[24][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][2]$_SDFFCE_PN0P_  (.D(_01312_),
    .DE(_00119_),
    .Q(\w[24][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][30]$_SDFFCE_PN0P_  (.D(_01313_),
    .DE(_00119_),
    .Q(\w[24][30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][31]$_SDFFCE_PN0P_  (.D(_01314_),
    .DE(_00119_),
    .Q(\w[24][31] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][3]$_SDFFCE_PN0P_  (.D(_01315_),
    .DE(_00119_),
    .Q(\w[24][3] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][4]$_SDFFCE_PN0P_  (.D(_01316_),
    .DE(_00119_),
    .Q(\w[24][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][5]$_SDFFCE_PN0P_  (.D(_01317_),
    .DE(_00119_),
    .Q(\w[24][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][6]$_SDFFCE_PN0P_  (.D(_01318_),
    .DE(_00119_),
    .Q(\w[24][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][7]$_SDFFCE_PN0P_  (.D(_01319_),
    .DE(_00119_),
    .Q(\w[24][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][8]$_SDFFCE_PN0P_  (.D(_01320_),
    .DE(_00119_),
    .Q(\w[24][8] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][9]$_SDFFCE_PN0P_  (.D(_01321_),
    .DE(_00119_),
    .Q(\w[24][9] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][0]$_SDFFCE_PN0P_  (.D(_01322_),
    .DE(_00087_),
    .Q(\w[25][0] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][10]$_SDFFCE_PN0P_  (.D(_01323_),
    .DE(_00087_),
    .Q(\w[25][10] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][11]$_SDFFCE_PN0P_  (.D(_01324_),
    .DE(_00087_),
    .Q(\w[25][11] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][12]$_SDFFCE_PN0P_  (.D(_01325_),
    .DE(_00087_),
    .Q(\w[25][12] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][13]$_SDFFCE_PN0P_  (.D(_01326_),
    .DE(_00087_),
    .Q(\w[25][13] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][14]$_SDFFCE_PN0P_  (.D(_01327_),
    .DE(_00087_),
    .Q(\w[25][14] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][15]$_SDFFCE_PN0P_  (.D(_01328_),
    .DE(_00087_),
    .Q(\w[25][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][16]$_SDFFCE_PN0P_  (.D(_01329_),
    .DE(_00087_),
    .Q(\w[25][16] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][17]$_SDFFCE_PN0P_  (.D(_01330_),
    .DE(_00087_),
    .Q(\w[25][17] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][18]$_SDFFCE_PN0P_  (.D(_01331_),
    .DE(_00087_),
    .Q(\w[25][18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][19]$_SDFFCE_PN0P_  (.D(_01332_),
    .DE(_00087_),
    .Q(\w[25][19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][1]$_SDFFCE_PN0P_  (.D(_01333_),
    .DE(_00087_),
    .Q(\w[25][1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][20]$_SDFFCE_PN0P_  (.D(_01334_),
    .DE(_00087_),
    .Q(\w[25][20] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][21]$_SDFFCE_PN0P_  (.D(_01335_),
    .DE(_00087_),
    .Q(\w[25][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][22]$_SDFFCE_PN0P_  (.D(_01336_),
    .DE(_00087_),
    .Q(\w[25][22] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][23]$_SDFFCE_PN0P_  (.D(_01337_),
    .DE(_00087_),
    .Q(\w[25][23] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][24]$_SDFFCE_PN0P_  (.D(_01338_),
    .DE(_00087_),
    .Q(\w[25][24] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][25]$_SDFFCE_PN0P_  (.D(_01339_),
    .DE(_00087_),
    .Q(\w[25][25] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][26]$_SDFFCE_PN0P_  (.D(_01340_),
    .DE(_00087_),
    .Q(\w[25][26] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][27]$_SDFFCE_PN0P_  (.D(_01341_),
    .DE(_00087_),
    .Q(\w[25][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][28]$_SDFFCE_PN0P_  (.D(_01342_),
    .DE(_00087_),
    .Q(\w[25][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][29]$_SDFFCE_PN0P_  (.D(_01343_),
    .DE(_00087_),
    .Q(\w[25][29] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][2]$_SDFFCE_PN0P_  (.D(_01344_),
    .DE(_00087_),
    .Q(\w[25][2] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][30]$_SDFFCE_PN0P_  (.D(_01345_),
    .DE(_00087_),
    .Q(\w[25][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][31]$_SDFFCE_PN0P_  (.D(_01346_),
    .DE(_00087_),
    .Q(\w[25][31] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][3]$_SDFFCE_PN0P_  (.D(_01347_),
    .DE(_00087_),
    .Q(\w[25][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][4]$_SDFFCE_PN0P_  (.D(_01348_),
    .DE(_00087_),
    .Q(\w[25][4] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][5]$_SDFFCE_PN0P_  (.D(_01349_),
    .DE(_00087_),
    .Q(\w[25][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][6]$_SDFFCE_PN0P_  (.D(_01350_),
    .DE(_00087_),
    .Q(\w[25][6] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][7]$_SDFFCE_PN0P_  (.D(_01351_),
    .DE(_00087_),
    .Q(\w[25][7] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][8]$_SDFFCE_PN0P_  (.D(_01352_),
    .DE(_00087_),
    .Q(\w[25][8] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][9]$_SDFFCE_PN0P_  (.D(_01353_),
    .DE(_00087_),
    .Q(\w[25][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][0]$_SDFFCE_PN0P_  (.D(_01354_),
    .DE(_00118_),
    .Q(\w[26][0] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][10]$_SDFFCE_PN0P_  (.D(_01355_),
    .DE(_00118_),
    .Q(\w[26][10] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][11]$_SDFFCE_PN0P_  (.D(_01356_),
    .DE(_00118_),
    .Q(\w[26][11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][12]$_SDFFCE_PN0P_  (.D(_01357_),
    .DE(_00118_),
    .Q(\w[26][12] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][13]$_SDFFCE_PN0P_  (.D(_01358_),
    .DE(_00118_),
    .Q(\w[26][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][14]$_SDFFCE_PN0P_  (.D(_01359_),
    .DE(_00118_),
    .Q(\w[26][14] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][15]$_SDFFCE_PN0P_  (.D(_01360_),
    .DE(_00118_),
    .Q(\w[26][15] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][16]$_SDFFCE_PN0P_  (.D(_01361_),
    .DE(_00118_),
    .Q(\w[26][16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][17]$_SDFFCE_PN0P_  (.D(_01362_),
    .DE(_00118_),
    .Q(\w[26][17] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][18]$_SDFFCE_PN0P_  (.D(_01363_),
    .DE(_00118_),
    .Q(\w[26][18] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][19]$_SDFFCE_PN0P_  (.D(_01364_),
    .DE(_00118_),
    .Q(\w[26][19] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][1]$_SDFFCE_PN0P_  (.D(_01365_),
    .DE(_00118_),
    .Q(\w[26][1] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][20]$_SDFFCE_PN0P_  (.D(_01366_),
    .DE(_00118_),
    .Q(\w[26][20] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][21]$_SDFFCE_PN0P_  (.D(_01367_),
    .DE(_00118_),
    .Q(\w[26][21] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][22]$_SDFFCE_PN0P_  (.D(_01368_),
    .DE(_00118_),
    .Q(\w[26][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][23]$_SDFFCE_PN0P_  (.D(_01369_),
    .DE(_00118_),
    .Q(\w[26][23] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][24]$_SDFFCE_PN0P_  (.D(_01370_),
    .DE(_00118_),
    .Q(\w[26][24] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][25]$_SDFFCE_PN0P_  (.D(_01371_),
    .DE(_00118_),
    .Q(\w[26][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][26]$_SDFFCE_PN0P_  (.D(_01372_),
    .DE(_00118_),
    .Q(\w[26][26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][27]$_SDFFCE_PN0P_  (.D(_01373_),
    .DE(_00118_),
    .Q(\w[26][27] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][28]$_SDFFCE_PN0P_  (.D(_01374_),
    .DE(_00118_),
    .Q(\w[26][28] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][29]$_SDFFCE_PN0P_  (.D(_01375_),
    .DE(_00118_),
    .Q(\w[26][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][2]$_SDFFCE_PN0P_  (.D(_01376_),
    .DE(_00118_),
    .Q(\w[26][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][30]$_SDFFCE_PN0P_  (.D(_01377_),
    .DE(_00118_),
    .Q(\w[26][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][31]$_SDFFCE_PN0P_  (.D(_01378_),
    .DE(_00118_),
    .Q(\w[26][31] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][3]$_SDFFCE_PN0P_  (.D(_01379_),
    .DE(_00118_),
    .Q(\w[26][3] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][4]$_SDFFCE_PN0P_  (.D(_01380_),
    .DE(_00118_),
    .Q(\w[26][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][5]$_SDFFCE_PN0P_  (.D(_01381_),
    .DE(_00118_),
    .Q(\w[26][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][6]$_SDFFCE_PN0P_  (.D(_01382_),
    .DE(_00118_),
    .Q(\w[26][6] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][7]$_SDFFCE_PN0P_  (.D(_01383_),
    .DE(_00118_),
    .Q(\w[26][7] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][8]$_SDFFCE_PN0P_  (.D(_01384_),
    .DE(_00118_),
    .Q(\w[26][8] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][9]$_SDFFCE_PN0P_  (.D(_01385_),
    .DE(_00118_),
    .Q(\w[26][9] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][0]$_SDFFCE_PN0P_  (.D(_01386_),
    .DE(_00086_),
    .Q(\w[27][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][10]$_SDFFCE_PN0P_  (.D(_01387_),
    .DE(_00086_),
    .Q(\w[27][10] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][11]$_SDFFCE_PN0P_  (.D(_01388_),
    .DE(_00086_),
    .Q(\w[27][11] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][12]$_SDFFCE_PN0P_  (.D(_01389_),
    .DE(_00086_),
    .Q(\w[27][12] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][13]$_SDFFCE_PN0P_  (.D(_01390_),
    .DE(_00086_),
    .Q(\w[27][13] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][14]$_SDFFCE_PN0P_  (.D(_01391_),
    .DE(_00086_),
    .Q(\w[27][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][15]$_SDFFCE_PN0P_  (.D(_01392_),
    .DE(_00086_),
    .Q(\w[27][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][16]$_SDFFCE_PN0P_  (.D(_01393_),
    .DE(_00086_),
    .Q(\w[27][16] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][17]$_SDFFCE_PN0P_  (.D(_01394_),
    .DE(_00086_),
    .Q(\w[27][17] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][18]$_SDFFCE_PN0P_  (.D(_01395_),
    .DE(_00086_),
    .Q(\w[27][18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][19]$_SDFFCE_PN0P_  (.D(_01396_),
    .DE(_00086_),
    .Q(\w[27][19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][1]$_SDFFCE_PN0P_  (.D(_01397_),
    .DE(_00086_),
    .Q(\w[27][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][20]$_SDFFCE_PN0P_  (.D(_01398_),
    .DE(_00086_),
    .Q(\w[27][20] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][21]$_SDFFCE_PN0P_  (.D(_01399_),
    .DE(_00086_),
    .Q(\w[27][21] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][22]$_SDFFCE_PN0P_  (.D(_01400_),
    .DE(_00086_),
    .Q(\w[27][22] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][23]$_SDFFCE_PN0P_  (.D(_01401_),
    .DE(_00086_),
    .Q(\w[27][23] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][24]$_SDFFCE_PN0P_  (.D(_01402_),
    .DE(_00086_),
    .Q(\w[27][24] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][25]$_SDFFCE_PN0P_  (.D(_01403_),
    .DE(_00086_),
    .Q(\w[27][25] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][26]$_SDFFCE_PN0P_  (.D(_01404_),
    .DE(_00086_),
    .Q(\w[27][26] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][27]$_SDFFCE_PN0P_  (.D(_01405_),
    .DE(_00086_),
    .Q(\w[27][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][28]$_SDFFCE_PN0P_  (.D(_01406_),
    .DE(_00086_),
    .Q(\w[27][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][29]$_SDFFCE_PN0P_  (.D(_01407_),
    .DE(_00086_),
    .Q(\w[27][29] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][2]$_SDFFCE_PN0P_  (.D(_01408_),
    .DE(_00086_),
    .Q(\w[27][2] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][30]$_SDFFCE_PN0P_  (.D(_01409_),
    .DE(_00086_),
    .Q(\w[27][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][31]$_SDFFCE_PN0P_  (.D(_01410_),
    .DE(_00086_),
    .Q(\w[27][31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][3]$_SDFFCE_PN0P_  (.D(_01411_),
    .DE(_00086_),
    .Q(\w[27][3] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][4]$_SDFFCE_PN0P_  (.D(_01412_),
    .DE(_00086_),
    .Q(\w[27][4] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][5]$_SDFFCE_PN0P_  (.D(_01413_),
    .DE(_00086_),
    .Q(\w[27][5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][6]$_SDFFCE_PN0P_  (.D(_01414_),
    .DE(_00086_),
    .Q(\w[27][6] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][7]$_SDFFCE_PN0P_  (.D(_01415_),
    .DE(_00086_),
    .Q(\w[27][7] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][8]$_SDFFCE_PN0P_  (.D(_01416_),
    .DE(_00086_),
    .Q(\w[27][8] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][9]$_SDFFCE_PN0P_  (.D(_01417_),
    .DE(_00086_),
    .Q(\w[27][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][0]$_SDFFCE_PN0P_  (.D(_01418_),
    .DE(_00117_),
    .Q(\w[28][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][10]$_SDFFCE_PN0P_  (.D(_01419_),
    .DE(_00117_),
    .Q(\w[28][10] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][11]$_SDFFCE_PN0P_  (.D(_01420_),
    .DE(_00117_),
    .Q(\w[28][11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][12]$_SDFFCE_PN0P_  (.D(_01421_),
    .DE(_00117_),
    .Q(\w[28][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][13]$_SDFFCE_PN0P_  (.D(_01422_),
    .DE(_00117_),
    .Q(\w[28][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][14]$_SDFFCE_PN0P_  (.D(_01423_),
    .DE(_00117_),
    .Q(\w[28][14] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][15]$_SDFFCE_PN0P_  (.D(_01424_),
    .DE(_00117_),
    .Q(\w[28][15] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][16]$_SDFFCE_PN0P_  (.D(_01425_),
    .DE(_00117_),
    .Q(\w[28][16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][17]$_SDFFCE_PN0P_  (.D(_01426_),
    .DE(_00117_),
    .Q(\w[28][17] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][18]$_SDFFCE_PN0P_  (.D(_01427_),
    .DE(_00117_),
    .Q(\w[28][18] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][19]$_SDFFCE_PN0P_  (.D(_01428_),
    .DE(_00117_),
    .Q(\w[28][19] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][1]$_SDFFCE_PN0P_  (.D(_01429_),
    .DE(_00117_),
    .Q(\w[28][1] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][20]$_SDFFCE_PN0P_  (.D(_01430_),
    .DE(_00117_),
    .Q(\w[28][20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][21]$_SDFFCE_PN0P_  (.D(_01431_),
    .DE(_00117_),
    .Q(\w[28][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][22]$_SDFFCE_PN0P_  (.D(_01432_),
    .DE(_00117_),
    .Q(\w[28][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][23]$_SDFFCE_PN0P_  (.D(_01433_),
    .DE(_00117_),
    .Q(\w[28][23] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][24]$_SDFFCE_PN0P_  (.D(_01434_),
    .DE(_00117_),
    .Q(\w[28][24] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][25]$_SDFFCE_PN0P_  (.D(_01435_),
    .DE(_00117_),
    .Q(\w[28][25] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][26]$_SDFFCE_PN0P_  (.D(_01436_),
    .DE(_00117_),
    .Q(\w[28][26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][27]$_SDFFCE_PN0P_  (.D(_01437_),
    .DE(_00117_),
    .Q(\w[28][27] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][28]$_SDFFCE_PN0P_  (.D(_01438_),
    .DE(_00117_),
    .Q(\w[28][28] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][29]$_SDFFCE_PN0P_  (.D(_01439_),
    .DE(_00117_),
    .Q(\w[28][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][2]$_SDFFCE_PN0P_  (.D(_01440_),
    .DE(_00117_),
    .Q(\w[28][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][30]$_SDFFCE_PN0P_  (.D(_01441_),
    .DE(_00117_),
    .Q(\w[28][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][31]$_SDFFCE_PN0P_  (.D(_01442_),
    .DE(_00117_),
    .Q(\w[28][31] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][3]$_SDFFCE_PN0P_  (.D(_01443_),
    .DE(_00117_),
    .Q(\w[28][3] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][4]$_SDFFCE_PN0P_  (.D(_01444_),
    .DE(_00117_),
    .Q(\w[28][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][5]$_SDFFCE_PN0P_  (.D(_01445_),
    .DE(_00117_),
    .Q(\w[28][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][6]$_SDFFCE_PN0P_  (.D(_01446_),
    .DE(_00117_),
    .Q(\w[28][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][7]$_SDFFCE_PN0P_  (.D(_01447_),
    .DE(_00117_),
    .Q(\w[28][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][8]$_SDFFCE_PN0P_  (.D(_01448_),
    .DE(_00117_),
    .Q(\w[28][8] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][9]$_SDFFCE_PN0P_  (.D(_01449_),
    .DE(_00117_),
    .Q(\w[28][9] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][0]$_SDFFCE_PN0P_  (.D(_01450_),
    .DE(_00085_),
    .Q(\w[29][0] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][10]$_SDFFCE_PN0P_  (.D(_01451_),
    .DE(_00085_),
    .Q(\w[29][10] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][11]$_SDFFCE_PN0P_  (.D(_01452_),
    .DE(_00085_),
    .Q(\w[29][11] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][12]$_SDFFCE_PN0P_  (.D(_01453_),
    .DE(_00085_),
    .Q(\w[29][12] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][13]$_SDFFCE_PN0P_  (.D(_01454_),
    .DE(_00085_),
    .Q(\w[29][13] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][14]$_SDFFCE_PN0P_  (.D(_01455_),
    .DE(_00085_),
    .Q(\w[29][14] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][15]$_SDFFCE_PN0P_  (.D(_01456_),
    .DE(_00085_),
    .Q(\w[29][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][16]$_SDFFCE_PN0P_  (.D(_01457_),
    .DE(_00085_),
    .Q(\w[29][16] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][17]$_SDFFCE_PN0P_  (.D(_01458_),
    .DE(_00085_),
    .Q(\w[29][17] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][18]$_SDFFCE_PN0P_  (.D(_01459_),
    .DE(_00085_),
    .Q(\w[29][18] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][19]$_SDFFCE_PN0P_  (.D(_01460_),
    .DE(_00085_),
    .Q(\w[29][19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][1]$_SDFFCE_PN0P_  (.D(_01461_),
    .DE(_00085_),
    .Q(\w[29][1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][20]$_SDFFCE_PN0P_  (.D(_01462_),
    .DE(_00085_),
    .Q(\w[29][20] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][21]$_SDFFCE_PN0P_  (.D(_01463_),
    .DE(_00085_),
    .Q(\w[29][21] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][22]$_SDFFCE_PN0P_  (.D(_01464_),
    .DE(_00085_),
    .Q(\w[29][22] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][23]$_SDFFCE_PN0P_  (.D(_01465_),
    .DE(_00085_),
    .Q(\w[29][23] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][24]$_SDFFCE_PN0P_  (.D(_01466_),
    .DE(_00085_),
    .Q(\w[29][24] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][25]$_SDFFCE_PN0P_  (.D(_01467_),
    .DE(_00085_),
    .Q(\w[29][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][26]$_SDFFCE_PN0P_  (.D(_01468_),
    .DE(_00085_),
    .Q(\w[29][26] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][27]$_SDFFCE_PN0P_  (.D(_01469_),
    .DE(_00085_),
    .Q(\w[29][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][28]$_SDFFCE_PN0P_  (.D(_01470_),
    .DE(_00085_),
    .Q(\w[29][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][29]$_SDFFCE_PN0P_  (.D(_01471_),
    .DE(_00085_),
    .Q(\w[29][29] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][2]$_SDFFCE_PN0P_  (.D(_01472_),
    .DE(_00085_),
    .Q(\w[29][2] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][30]$_SDFFCE_PN0P_  (.D(_01473_),
    .DE(_00085_),
    .Q(\w[29][30] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][31]$_SDFFCE_PN0P_  (.D(_01474_),
    .DE(_00085_),
    .Q(\w[29][31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][3]$_SDFFCE_PN0P_  (.D(_01475_),
    .DE(_00085_),
    .Q(\w[29][3] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][4]$_SDFFCE_PN0P_  (.D(_01476_),
    .DE(_00085_),
    .Q(\w[29][4] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][5]$_SDFFCE_PN0P_  (.D(_01477_),
    .DE(_00085_),
    .Q(\w[29][5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][6]$_SDFFCE_PN0P_  (.D(_01478_),
    .DE(_00085_),
    .Q(\w[29][6] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][7]$_SDFFCE_PN0P_  (.D(_01479_),
    .DE(_00085_),
    .Q(\w[29][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][8]$_SDFFCE_PN0P_  (.D(_01480_),
    .DE(_00085_),
    .Q(\w[29][8] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][9]$_SDFFCE_PN0P_  (.D(_01481_),
    .DE(_00085_),
    .Q(\w[29][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][0]$_DFFE_PP_  (.D(_00385_),
    .DE(_00116_),
    .Q(\w[2][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][10]$_DFFE_PP_  (.D(_00386_),
    .DE(_00116_),
    .Q(\w[2][10] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][11]$_DFFE_PP_  (.D(_00387_),
    .DE(_00116_),
    .Q(\w[2][11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][12]$_DFFE_PP_  (.D(_00388_),
    .DE(_00116_),
    .Q(\w[2][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][13]$_DFFE_PP_  (.D(_00389_),
    .DE(_00116_),
    .Q(\w[2][13] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][14]$_DFFE_PP_  (.D(_00390_),
    .DE(_00116_),
    .Q(\w[2][14] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][15]$_DFFE_PP_  (.D(_00391_),
    .DE(_00116_),
    .Q(\w[2][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][16]$_DFFE_PP_  (.D(_00392_),
    .DE(_00116_),
    .Q(\w[2][16] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][17]$_DFFE_PP_  (.D(_00393_),
    .DE(_00116_),
    .Q(\w[2][17] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][18]$_DFFE_PP_  (.D(_00394_),
    .DE(_00116_),
    .Q(\w[2][18] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][19]$_DFFE_PP_  (.D(_00395_),
    .DE(_00116_),
    .Q(\w[2][19] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][1]$_DFFE_PP_  (.D(_00396_),
    .DE(_00116_),
    .Q(\w[2][1] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][20]$_DFFE_PP_  (.D(_00397_),
    .DE(_00116_),
    .Q(\w[2][20] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][21]$_DFFE_PP_  (.D(_00398_),
    .DE(_00116_),
    .Q(\w[2][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][22]$_DFFE_PP_  (.D(_00399_),
    .DE(_00116_),
    .Q(\w[2][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][23]$_DFFE_PP_  (.D(_00400_),
    .DE(_00116_),
    .Q(\w[2][23] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][24]$_DFFE_PP_  (.D(_00401_),
    .DE(_00116_),
    .Q(\w[2][24] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][25]$_DFFE_PP_  (.D(_00402_),
    .DE(_00116_),
    .Q(\w[2][25] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][26]$_DFFE_PP_  (.D(_00403_),
    .DE(_00116_),
    .Q(\w[2][26] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][27]$_DFFE_PP_  (.D(_00404_),
    .DE(_00116_),
    .Q(\w[2][27] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][28]$_DFFE_PP_  (.D(_00405_),
    .DE(_00116_),
    .Q(\w[2][28] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][29]$_DFFE_PP_  (.D(_00406_),
    .DE(_00116_),
    .Q(\w[2][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][2]$_DFFE_PP_  (.D(_00407_),
    .DE(_00116_),
    .Q(\w[2][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][30]$_DFFE_PP_  (.D(_00408_),
    .DE(_00116_),
    .Q(\w[2][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][31]$_DFFE_PP_  (.D(_00409_),
    .DE(_00116_),
    .Q(\w[2][31] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][3]$_DFFE_PP_  (.D(_00410_),
    .DE(_00116_),
    .Q(\w[2][3] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][4]$_DFFE_PP_  (.D(_00411_),
    .DE(_00116_),
    .Q(\w[2][4] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][5]$_DFFE_PP_  (.D(_00412_),
    .DE(_00116_),
    .Q(\w[2][5] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][6]$_DFFE_PP_  (.D(_00413_),
    .DE(_00116_),
    .Q(\w[2][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][7]$_DFFE_PP_  (.D(_00414_),
    .DE(_00116_),
    .Q(\w[2][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][8]$_DFFE_PP_  (.D(_00415_),
    .DE(_00116_),
    .Q(\w[2][8] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][9]$_DFFE_PP_  (.D(_00416_),
    .DE(_00116_),
    .Q(\w[2][9] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][0]$_SDFFCE_PN0P_  (.D(_01482_),
    .DE(_00115_),
    .Q(\w[30][0] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][10]$_SDFFCE_PN0P_  (.D(_01483_),
    .DE(_00115_),
    .Q(\w[30][10] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][11]$_SDFFCE_PN0P_  (.D(_01484_),
    .DE(_00115_),
    .Q(\w[30][11] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][12]$_SDFFCE_PN0P_  (.D(_01485_),
    .DE(_00115_),
    .Q(\w[30][12] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][13]$_SDFFCE_PN0P_  (.D(_01486_),
    .DE(_00115_),
    .Q(\w[30][13] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][14]$_SDFFCE_PN0P_  (.D(_01487_),
    .DE(_00115_),
    .Q(\w[30][14] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][15]$_SDFFCE_PN0P_  (.D(_01488_),
    .DE(_00115_),
    .Q(\w[30][15] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][16]$_SDFFCE_PN0P_  (.D(_01489_),
    .DE(_00115_),
    .Q(\w[30][16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][17]$_SDFFCE_PN0P_  (.D(_01490_),
    .DE(_00115_),
    .Q(\w[30][17] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][18]$_SDFFCE_PN0P_  (.D(_01491_),
    .DE(_00115_),
    .Q(\w[30][18] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][19]$_SDFFCE_PN0P_  (.D(_01492_),
    .DE(_00115_),
    .Q(\w[30][19] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][1]$_SDFFCE_PN0P_  (.D(_01493_),
    .DE(_00115_),
    .Q(\w[30][1] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][20]$_SDFFCE_PN0P_  (.D(_01494_),
    .DE(_00115_),
    .Q(\w[30][20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][21]$_SDFFCE_PN0P_  (.D(_01495_),
    .DE(_00115_),
    .Q(\w[30][21] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][22]$_SDFFCE_PN0P_  (.D(_01496_),
    .DE(_00115_),
    .Q(\w[30][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][23]$_SDFFCE_PN0P_  (.D(_01497_),
    .DE(_00115_),
    .Q(\w[30][23] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][24]$_SDFFCE_PN0P_  (.D(_01498_),
    .DE(_00115_),
    .Q(\w[30][24] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][25]$_SDFFCE_PN0P_  (.D(_01499_),
    .DE(_00115_),
    .Q(\w[30][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][26]$_SDFFCE_PN0P_  (.D(_01500_),
    .DE(_00115_),
    .Q(\w[30][26] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][27]$_SDFFCE_PN0P_  (.D(_01501_),
    .DE(_00115_),
    .Q(\w[30][27] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][28]$_SDFFCE_PN0P_  (.D(_01502_),
    .DE(_00115_),
    .Q(\w[30][28] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][29]$_SDFFCE_PN0P_  (.D(_01503_),
    .DE(_00115_),
    .Q(\w[30][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][2]$_SDFFCE_PN0P_  (.D(_01504_),
    .DE(_00115_),
    .Q(\w[30][2] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][30]$_SDFFCE_PN0P_  (.D(_01505_),
    .DE(_00115_),
    .Q(\w[30][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][31]$_SDFFCE_PN0P_  (.D(_01506_),
    .DE(_00115_),
    .Q(\w[30][31] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][3]$_SDFFCE_PN0P_  (.D(_01507_),
    .DE(_00115_),
    .Q(\w[30][3] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][4]$_SDFFCE_PN0P_  (.D(_01508_),
    .DE(_00115_),
    .Q(\w[30][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][5]$_SDFFCE_PN0P_  (.D(_01509_),
    .DE(_00115_),
    .Q(\w[30][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][6]$_SDFFCE_PN0P_  (.D(_01510_),
    .DE(_00115_),
    .Q(\w[30][6] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][7]$_SDFFCE_PN0P_  (.D(_01511_),
    .DE(_00115_),
    .Q(\w[30][7] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][8]$_SDFFCE_PN0P_  (.D(_01512_),
    .DE(_00115_),
    .Q(\w[30][8] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][9]$_SDFFCE_PN0P_  (.D(_01513_),
    .DE(_00115_),
    .Q(\w[30][9] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][0]$_SDFFCE_PN0P_  (.D(_01514_),
    .DE(_00084_),
    .Q(\w[31][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][10]$_SDFFCE_PN0P_  (.D(_01515_),
    .DE(_00084_),
    .Q(\w[31][10] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][11]$_SDFFCE_PN0P_  (.D(_01516_),
    .DE(_00084_),
    .Q(\w[31][11] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][12]$_SDFFCE_PN0P_  (.D(_01517_),
    .DE(_00084_),
    .Q(\w[31][12] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][13]$_SDFFCE_PN0P_  (.D(_01518_),
    .DE(_00084_),
    .Q(\w[31][13] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][14]$_SDFFCE_PN0P_  (.D(_01519_),
    .DE(_00084_),
    .Q(\w[31][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][15]$_SDFFCE_PN0P_  (.D(_01520_),
    .DE(_00084_),
    .Q(\w[31][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][16]$_SDFFCE_PN0P_  (.D(_01521_),
    .DE(_00084_),
    .Q(\w[31][16] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][17]$_SDFFCE_PN0P_  (.D(_01522_),
    .DE(_00084_),
    .Q(\w[31][17] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][18]$_SDFFCE_PN0P_  (.D(_01523_),
    .DE(_00084_),
    .Q(\w[31][18] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][19]$_SDFFCE_PN0P_  (.D(_01524_),
    .DE(_00084_),
    .Q(\w[31][19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][1]$_SDFFCE_PN0P_  (.D(_01525_),
    .DE(_00084_),
    .Q(\w[31][1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][20]$_SDFFCE_PN0P_  (.D(_01526_),
    .DE(_00084_),
    .Q(\w[31][20] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][21]$_SDFFCE_PN0P_  (.D(_01527_),
    .DE(_00084_),
    .Q(\w[31][21] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][22]$_SDFFCE_PN0P_  (.D(_01528_),
    .DE(_00084_),
    .Q(\w[31][22] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][23]$_SDFFCE_PN0P_  (.D(_01529_),
    .DE(_00084_),
    .Q(\w[31][23] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][24]$_SDFFCE_PN0P_  (.D(_01530_),
    .DE(_00084_),
    .Q(\w[31][24] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][25]$_SDFFCE_PN0P_  (.D(_01531_),
    .DE(_00084_),
    .Q(\w[31][25] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][26]$_SDFFCE_PN0P_  (.D(_01532_),
    .DE(_00084_),
    .Q(\w[31][26] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][27]$_SDFFCE_PN0P_  (.D(_01533_),
    .DE(_00084_),
    .Q(\w[31][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][28]$_SDFFCE_PN0P_  (.D(_01534_),
    .DE(_00084_),
    .Q(\w[31][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][29]$_SDFFCE_PN0P_  (.D(_01535_),
    .DE(_00084_),
    .Q(\w[31][29] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][2]$_SDFFCE_PN0P_  (.D(_01536_),
    .DE(_00084_),
    .Q(\w[31][2] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][30]$_SDFFCE_PN0P_  (.D(_01537_),
    .DE(_00084_),
    .Q(\w[31][30] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][31]$_SDFFCE_PN0P_  (.D(_01538_),
    .DE(_00084_),
    .Q(\w[31][31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][3]$_SDFFCE_PN0P_  (.D(_01539_),
    .DE(_00084_),
    .Q(\w[31][3] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][4]$_SDFFCE_PN0P_  (.D(_01540_),
    .DE(_00084_),
    .Q(\w[31][4] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][5]$_SDFFCE_PN0P_  (.D(_01541_),
    .DE(_00084_),
    .Q(\w[31][5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][6]$_SDFFCE_PN0P_  (.D(_01542_),
    .DE(_00084_),
    .Q(\w[31][6] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][7]$_SDFFCE_PN0P_  (.D(_01543_),
    .DE(_00084_),
    .Q(\w[31][7] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][8]$_SDFFCE_PN0P_  (.D(_01544_),
    .DE(_00084_),
    .Q(\w[31][8] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][9]$_SDFFCE_PN0P_  (.D(_01545_),
    .DE(_00084_),
    .Q(\w[31][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][0]$_SDFFCE_PN0P_  (.D(_01546_),
    .DE(_00114_),
    .Q(\w[32][0] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][10]$_SDFFCE_PN0P_  (.D(_01547_),
    .DE(_00114_),
    .Q(\w[32][10] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][11]$_SDFFCE_PN0P_  (.D(_01548_),
    .DE(_00114_),
    .Q(\w[32][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][12]$_SDFFCE_PN0P_  (.D(_01549_),
    .DE(_00114_),
    .Q(\w[32][12] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][13]$_SDFFCE_PN0P_  (.D(_01550_),
    .DE(_00114_),
    .Q(\w[32][13] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][14]$_SDFFCE_PN0P_  (.D(_01551_),
    .DE(_00114_),
    .Q(\w[32][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][15]$_SDFFCE_PN0P_  (.D(_01552_),
    .DE(_00114_),
    .Q(\w[32][15] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][16]$_SDFFCE_PN0P_  (.D(_01553_),
    .DE(_00114_),
    .Q(\w[32][16] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][17]$_SDFFCE_PN0P_  (.D(_01554_),
    .DE(_00114_),
    .Q(\w[32][17] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][18]$_SDFFCE_PN0P_  (.D(_01555_),
    .DE(_00114_),
    .Q(\w[32][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][19]$_SDFFCE_PN0P_  (.D(_01556_),
    .DE(_00114_),
    .Q(\w[32][19] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][1]$_SDFFCE_PN0P_  (.D(_01557_),
    .DE(_00114_),
    .Q(\w[32][1] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][20]$_SDFFCE_PN0P_  (.D(_01558_),
    .DE(_00114_),
    .Q(\w[32][20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][21]$_SDFFCE_PN0P_  (.D(_01559_),
    .DE(_00114_),
    .Q(\w[32][21] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][22]$_SDFFCE_PN0P_  (.D(_01560_),
    .DE(_00114_),
    .Q(\w[32][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][23]$_SDFFCE_PN0P_  (.D(_01561_),
    .DE(_00114_),
    .Q(\w[32][23] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][24]$_SDFFCE_PN0P_  (.D(_01562_),
    .DE(_00114_),
    .Q(\w[32][24] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][25]$_SDFFCE_PN0P_  (.D(_01563_),
    .DE(_00114_),
    .Q(\w[32][25] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][26]$_SDFFCE_PN0P_  (.D(_01564_),
    .DE(_00114_),
    .Q(\w[32][26] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][27]$_SDFFCE_PN0P_  (.D(_01565_),
    .DE(_00114_),
    .Q(\w[32][27] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][28]$_SDFFCE_PN0P_  (.D(_01566_),
    .DE(_00114_),
    .Q(\w[32][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][29]$_SDFFCE_PN0P_  (.D(_01567_),
    .DE(_00114_),
    .Q(\w[32][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][2]$_SDFFCE_PN0P_  (.D(_01568_),
    .DE(_00114_),
    .Q(\w[32][2] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][30]$_SDFFCE_PN0P_  (.D(_01569_),
    .DE(_00114_),
    .Q(\w[32][30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][31]$_SDFFCE_PN0P_  (.D(_01570_),
    .DE(_00114_),
    .Q(\w[32][31] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][3]$_SDFFCE_PN0P_  (.D(_01571_),
    .DE(_00114_),
    .Q(\w[32][3] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][4]$_SDFFCE_PN0P_  (.D(_01572_),
    .DE(_00114_),
    .Q(\w[32][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][5]$_SDFFCE_PN0P_  (.D(_01573_),
    .DE(_00114_),
    .Q(\w[32][5] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][6]$_SDFFCE_PN0P_  (.D(_01574_),
    .DE(_00114_),
    .Q(\w[32][6] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][7]$_SDFFCE_PN0P_  (.D(_01575_),
    .DE(_00114_),
    .Q(\w[32][7] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][8]$_SDFFCE_PN0P_  (.D(_01576_),
    .DE(_00114_),
    .Q(\w[32][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][9]$_SDFFCE_PN0P_  (.D(_01577_),
    .DE(_00114_),
    .Q(\w[32][9] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][0]$_SDFFCE_PN0P_  (.D(_01578_),
    .DE(_00083_),
    .Q(\w[33][0] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][10]$_SDFFCE_PN0P_  (.D(_01579_),
    .DE(_00083_),
    .Q(\w[33][10] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][11]$_SDFFCE_PN0P_  (.D(_01580_),
    .DE(_00083_),
    .Q(\w[33][11] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][12]$_SDFFCE_PN0P_  (.D(_01581_),
    .DE(_00083_),
    .Q(\w[33][12] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][13]$_SDFFCE_PN0P_  (.D(_01582_),
    .DE(_00083_),
    .Q(\w[33][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][14]$_SDFFCE_PN0P_  (.D(_01583_),
    .DE(_00083_),
    .Q(\w[33][14] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][15]$_SDFFCE_PN0P_  (.D(_01584_),
    .DE(_00083_),
    .Q(\w[33][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][16]$_SDFFCE_PN0P_  (.D(_01585_),
    .DE(_00083_),
    .Q(\w[33][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][17]$_SDFFCE_PN0P_  (.D(_01586_),
    .DE(_00083_),
    .Q(\w[33][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][18]$_SDFFCE_PN0P_  (.D(_01587_),
    .DE(_00083_),
    .Q(\w[33][18] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][19]$_SDFFCE_PN0P_  (.D(_01588_),
    .DE(_00083_),
    .Q(\w[33][19] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][1]$_SDFFCE_PN0P_  (.D(_01589_),
    .DE(_00083_),
    .Q(\w[33][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][20]$_SDFFCE_PN0P_  (.D(_01590_),
    .DE(_00083_),
    .Q(\w[33][20] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][21]$_SDFFCE_PN0P_  (.D(_01591_),
    .DE(_00083_),
    .Q(\w[33][21] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][22]$_SDFFCE_PN0P_  (.D(_01592_),
    .DE(_00083_),
    .Q(\w[33][22] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][23]$_SDFFCE_PN0P_  (.D(_01593_),
    .DE(_00083_),
    .Q(\w[33][23] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][24]$_SDFFCE_PN0P_  (.D(_01594_),
    .DE(_00083_),
    .Q(\w[33][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][25]$_SDFFCE_PN0P_  (.D(_01595_),
    .DE(_00083_),
    .Q(\w[33][25] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][26]$_SDFFCE_PN0P_  (.D(_01596_),
    .DE(_00083_),
    .Q(\w[33][26] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][27]$_SDFFCE_PN0P_  (.D(_01597_),
    .DE(_00083_),
    .Q(\w[33][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][28]$_SDFFCE_PN0P_  (.D(_01598_),
    .DE(_00083_),
    .Q(\w[33][28] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][29]$_SDFFCE_PN0P_  (.D(_01599_),
    .DE(_00083_),
    .Q(\w[33][29] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][2]$_SDFFCE_PN0P_  (.D(_01600_),
    .DE(_00083_),
    .Q(\w[33][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][30]$_SDFFCE_PN0P_  (.D(_01601_),
    .DE(_00083_),
    .Q(\w[33][30] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][31]$_SDFFCE_PN0P_  (.D(_01602_),
    .DE(_00083_),
    .Q(\w[33][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][3]$_SDFFCE_PN0P_  (.D(_01603_),
    .DE(_00083_),
    .Q(\w[33][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][4]$_SDFFCE_PN0P_  (.D(_01604_),
    .DE(_00083_),
    .Q(\w[33][4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][5]$_SDFFCE_PN0P_  (.D(_01605_),
    .DE(_00083_),
    .Q(\w[33][5] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][6]$_SDFFCE_PN0P_  (.D(_01606_),
    .DE(_00083_),
    .Q(\w[33][6] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][7]$_SDFFCE_PN0P_  (.D(_01607_),
    .DE(_00083_),
    .Q(\w[33][7] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][8]$_SDFFCE_PN0P_  (.D(_01608_),
    .DE(_00083_),
    .Q(\w[33][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][9]$_SDFFCE_PN0P_  (.D(_01609_),
    .DE(_00083_),
    .Q(\w[33][9] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][0]$_SDFFCE_PN0P_  (.D(_01610_),
    .DE(_00113_),
    .Q(\w[34][0] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][10]$_SDFFCE_PN0P_  (.D(_01611_),
    .DE(_00113_),
    .Q(\w[34][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][11]$_SDFFCE_PN0P_  (.D(_01612_),
    .DE(_00113_),
    .Q(\w[34][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][12]$_SDFFCE_PN0P_  (.D(_01613_),
    .DE(_00113_),
    .Q(\w[34][12] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][13]$_SDFFCE_PN0P_  (.D(_01614_),
    .DE(_00113_),
    .Q(\w[34][13] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][14]$_SDFFCE_PN0P_  (.D(_01615_),
    .DE(_00113_),
    .Q(\w[34][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][15]$_SDFFCE_PN0P_  (.D(_01616_),
    .DE(_00113_),
    .Q(\w[34][15] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][16]$_SDFFCE_PN0P_  (.D(_01617_),
    .DE(_00113_),
    .Q(\w[34][16] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][17]$_SDFFCE_PN0P_  (.D(_01618_),
    .DE(_00113_),
    .Q(\w[34][17] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][18]$_SDFFCE_PN0P_  (.D(_01619_),
    .DE(_00113_),
    .Q(\w[34][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][19]$_SDFFCE_PN0P_  (.D(_01620_),
    .DE(_00113_),
    .Q(\w[34][19] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][1]$_SDFFCE_PN0P_  (.D(_01621_),
    .DE(_00113_),
    .Q(\w[34][1] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][20]$_SDFFCE_PN0P_  (.D(_01622_),
    .DE(_00113_),
    .Q(\w[34][20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][21]$_SDFFCE_PN0P_  (.D(_01623_),
    .DE(_00113_),
    .Q(\w[34][21] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][22]$_SDFFCE_PN0P_  (.D(_01624_),
    .DE(_00113_),
    .Q(\w[34][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][23]$_SDFFCE_PN0P_  (.D(_01625_),
    .DE(_00113_),
    .Q(\w[34][23] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][24]$_SDFFCE_PN0P_  (.D(_01626_),
    .DE(_00113_),
    .Q(\w[34][24] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][25]$_SDFFCE_PN0P_  (.D(_01627_),
    .DE(_00113_),
    .Q(\w[34][25] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][26]$_SDFFCE_PN0P_  (.D(_01628_),
    .DE(_00113_),
    .Q(\w[34][26] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][27]$_SDFFCE_PN0P_  (.D(_01629_),
    .DE(_00113_),
    .Q(\w[34][27] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][28]$_SDFFCE_PN0P_  (.D(_01630_),
    .DE(_00113_),
    .Q(\w[34][28] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][29]$_SDFFCE_PN0P_  (.D(_01631_),
    .DE(_00113_),
    .Q(\w[34][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][2]$_SDFFCE_PN0P_  (.D(_01632_),
    .DE(_00113_),
    .Q(\w[34][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][30]$_SDFFCE_PN0P_  (.D(_01633_),
    .DE(_00113_),
    .Q(\w[34][30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][31]$_SDFFCE_PN0P_  (.D(_01634_),
    .DE(_00113_),
    .Q(\w[34][31] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][3]$_SDFFCE_PN0P_  (.D(_01635_),
    .DE(_00113_),
    .Q(\w[34][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][4]$_SDFFCE_PN0P_  (.D(_01636_),
    .DE(_00113_),
    .Q(\w[34][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][5]$_SDFFCE_PN0P_  (.D(_01637_),
    .DE(_00113_),
    .Q(\w[34][5] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][6]$_SDFFCE_PN0P_  (.D(_01638_),
    .DE(_00113_),
    .Q(\w[34][6] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][7]$_SDFFCE_PN0P_  (.D(_01639_),
    .DE(_00113_),
    .Q(\w[34][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][8]$_SDFFCE_PN0P_  (.D(_01640_),
    .DE(_00113_),
    .Q(\w[34][8] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][9]$_SDFFCE_PN0P_  (.D(_01641_),
    .DE(_00113_),
    .Q(\w[34][9] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][0]$_SDFFCE_PN0P_  (.D(_01642_),
    .DE(_00082_),
    .Q(\w[35][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][10]$_SDFFCE_PN0P_  (.D(_01643_),
    .DE(_00082_),
    .Q(\w[35][10] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][11]$_SDFFCE_PN0P_  (.D(_01644_),
    .DE(_00082_),
    .Q(\w[35][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][12]$_SDFFCE_PN0P_  (.D(_01645_),
    .DE(_00082_),
    .Q(\w[35][12] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][13]$_SDFFCE_PN0P_  (.D(_01646_),
    .DE(_00082_),
    .Q(\w[35][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][14]$_SDFFCE_PN0P_  (.D(_01647_),
    .DE(_00082_),
    .Q(\w[35][14] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][15]$_SDFFCE_PN0P_  (.D(_01648_),
    .DE(_00082_),
    .Q(\w[35][15] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][16]$_SDFFCE_PN0P_  (.D(_01649_),
    .DE(_00082_),
    .Q(\w[35][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][17]$_SDFFCE_PN0P_  (.D(_01650_),
    .DE(_00082_),
    .Q(\w[35][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][18]$_SDFFCE_PN0P_  (.D(_01651_),
    .DE(_00082_),
    .Q(\w[35][18] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][19]$_SDFFCE_PN0P_  (.D(_01652_),
    .DE(_00082_),
    .Q(\w[35][19] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][1]$_SDFFCE_PN0P_  (.D(_01653_),
    .DE(_00082_),
    .Q(\w[35][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][20]$_SDFFCE_PN0P_  (.D(_01654_),
    .DE(_00082_),
    .Q(\w[35][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][21]$_SDFFCE_PN0P_  (.D(_01655_),
    .DE(_00082_),
    .Q(\w[35][21] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][22]$_SDFFCE_PN0P_  (.D(_01656_),
    .DE(_00082_),
    .Q(\w[35][22] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][23]$_SDFFCE_PN0P_  (.D(_01657_),
    .DE(_00082_),
    .Q(\w[35][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][24]$_SDFFCE_PN0P_  (.D(_01658_),
    .DE(_00082_),
    .Q(\w[35][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][25]$_SDFFCE_PN0P_  (.D(_01659_),
    .DE(_00082_),
    .Q(\w[35][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][26]$_SDFFCE_PN0P_  (.D(_01660_),
    .DE(_00082_),
    .Q(\w[35][26] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][27]$_SDFFCE_PN0P_  (.D(_01661_),
    .DE(_00082_),
    .Q(\w[35][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][28]$_SDFFCE_PN0P_  (.D(_01662_),
    .DE(_00082_),
    .Q(\w[35][28] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][29]$_SDFFCE_PN0P_  (.D(_01663_),
    .DE(_00082_),
    .Q(\w[35][29] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][2]$_SDFFCE_PN0P_  (.D(_01664_),
    .DE(_00082_),
    .Q(\w[35][2] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][30]$_SDFFCE_PN0P_  (.D(_01665_),
    .DE(_00082_),
    .Q(\w[35][30] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][31]$_SDFFCE_PN0P_  (.D(_01666_),
    .DE(_00082_),
    .Q(\w[35][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][3]$_SDFFCE_PN0P_  (.D(_01667_),
    .DE(_00082_),
    .Q(\w[35][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][4]$_SDFFCE_PN0P_  (.D(_01668_),
    .DE(_00082_),
    .Q(\w[35][4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][5]$_SDFFCE_PN0P_  (.D(_01669_),
    .DE(_00082_),
    .Q(\w[35][5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][6]$_SDFFCE_PN0P_  (.D(_01670_),
    .DE(_00082_),
    .Q(\w[35][6] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][7]$_SDFFCE_PN0P_  (.D(_01671_),
    .DE(_00082_),
    .Q(\w[35][7] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][8]$_SDFFCE_PN0P_  (.D(_01672_),
    .DE(_00082_),
    .Q(\w[35][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][9]$_SDFFCE_PN0P_  (.D(_01673_),
    .DE(_00082_),
    .Q(\w[35][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][0]$_SDFFCE_PN0P_  (.D(_01674_),
    .DE(_00112_),
    .Q(\w[36][0] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][10]$_SDFFCE_PN0P_  (.D(_01675_),
    .DE(_00112_),
    .Q(\w[36][10] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][11]$_SDFFCE_PN0P_  (.D(_01676_),
    .DE(_00112_),
    .Q(\w[36][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][12]$_SDFFCE_PN0P_  (.D(_01677_),
    .DE(_00112_),
    .Q(\w[36][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][13]$_SDFFCE_PN0P_  (.D(_01678_),
    .DE(_00112_),
    .Q(\w[36][13] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][14]$_SDFFCE_PN0P_  (.D(_01679_),
    .DE(_00112_),
    .Q(\w[36][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][15]$_SDFFCE_PN0P_  (.D(_01680_),
    .DE(_00112_),
    .Q(\w[36][15] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][16]$_SDFFCE_PN0P_  (.D(_01681_),
    .DE(_00112_),
    .Q(\w[36][16] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][17]$_SDFFCE_PN0P_  (.D(_01682_),
    .DE(_00112_),
    .Q(\w[36][17] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][18]$_SDFFCE_PN0P_  (.D(_01683_),
    .DE(_00112_),
    .Q(\w[36][18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][19]$_SDFFCE_PN0P_  (.D(_01684_),
    .DE(_00112_),
    .Q(\w[36][19] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][1]$_SDFFCE_PN0P_  (.D(_01685_),
    .DE(_00112_),
    .Q(\w[36][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][20]$_SDFFCE_PN0P_  (.D(_01686_),
    .DE(_00112_),
    .Q(\w[36][20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][21]$_SDFFCE_PN0P_  (.D(_01687_),
    .DE(_00112_),
    .Q(\w[36][21] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][22]$_SDFFCE_PN0P_  (.D(_01688_),
    .DE(_00112_),
    .Q(\w[36][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][23]$_SDFFCE_PN0P_  (.D(_01689_),
    .DE(_00112_),
    .Q(\w[36][23] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][24]$_SDFFCE_PN0P_  (.D(_01690_),
    .DE(_00112_),
    .Q(\w[36][24] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][25]$_SDFFCE_PN0P_  (.D(_01691_),
    .DE(_00112_),
    .Q(\w[36][25] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][26]$_SDFFCE_PN0P_  (.D(_01692_),
    .DE(_00112_),
    .Q(\w[36][26] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][27]$_SDFFCE_PN0P_  (.D(_01693_),
    .DE(_00112_),
    .Q(\w[36][27] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][28]$_SDFFCE_PN0P_  (.D(_01694_),
    .DE(_00112_),
    .Q(\w[36][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][29]$_SDFFCE_PN0P_  (.D(_01695_),
    .DE(_00112_),
    .Q(\w[36][29] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][2]$_SDFFCE_PN0P_  (.D(_01696_),
    .DE(_00112_),
    .Q(\w[36][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][30]$_SDFFCE_PN0P_  (.D(_01697_),
    .DE(_00112_),
    .Q(\w[36][30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][31]$_SDFFCE_PN0P_  (.D(_01698_),
    .DE(_00112_),
    .Q(\w[36][31] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][3]$_SDFFCE_PN0P_  (.D(_01699_),
    .DE(_00112_),
    .Q(\w[36][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][4]$_SDFFCE_PN0P_  (.D(_01700_),
    .DE(_00112_),
    .Q(\w[36][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][5]$_SDFFCE_PN0P_  (.D(_01701_),
    .DE(_00112_),
    .Q(\w[36][5] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][6]$_SDFFCE_PN0P_  (.D(_01702_),
    .DE(_00112_),
    .Q(\w[36][6] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][7]$_SDFFCE_PN0P_  (.D(_01703_),
    .DE(_00112_),
    .Q(\w[36][7] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][8]$_SDFFCE_PN0P_  (.D(_01704_),
    .DE(_00112_),
    .Q(\w[36][8] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][9]$_SDFFCE_PN0P_  (.D(_01705_),
    .DE(_00112_),
    .Q(\w[36][9] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][0]$_SDFFCE_PN0P_  (.D(_01706_),
    .DE(_00081_),
    .Q(\w[37][0] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][10]$_SDFFCE_PN0P_  (.D(_01707_),
    .DE(_00081_),
    .Q(\w[37][10] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][11]$_SDFFCE_PN0P_  (.D(_01708_),
    .DE(_00081_),
    .Q(\w[37][11] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][12]$_SDFFCE_PN0P_  (.D(_01709_),
    .DE(_00081_),
    .Q(\w[37][12] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][13]$_SDFFCE_PN0P_  (.D(_01710_),
    .DE(_00081_),
    .Q(\w[37][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][14]$_SDFFCE_PN0P_  (.D(_01711_),
    .DE(_00081_),
    .Q(\w[37][14] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][15]$_SDFFCE_PN0P_  (.D(_01712_),
    .DE(_00081_),
    .Q(\w[37][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][16]$_SDFFCE_PN0P_  (.D(_01713_),
    .DE(_00081_),
    .Q(\w[37][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][17]$_SDFFCE_PN0P_  (.D(_01714_),
    .DE(_00081_),
    .Q(\w[37][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][18]$_SDFFCE_PN0P_  (.D(_01715_),
    .DE(_00081_),
    .Q(\w[37][18] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][19]$_SDFFCE_PN0P_  (.D(_01716_),
    .DE(_00081_),
    .Q(\w[37][19] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][1]$_SDFFCE_PN0P_  (.D(_01717_),
    .DE(_00081_),
    .Q(\w[37][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][20]$_SDFFCE_PN0P_  (.D(_01718_),
    .DE(_00081_),
    .Q(\w[37][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][21]$_SDFFCE_PN0P_  (.D(_01719_),
    .DE(_00081_),
    .Q(\w[37][21] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][22]$_SDFFCE_PN0P_  (.D(_01720_),
    .DE(_00081_),
    .Q(\w[37][22] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][23]$_SDFFCE_PN0P_  (.D(_01721_),
    .DE(_00081_),
    .Q(\w[37][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][24]$_SDFFCE_PN0P_  (.D(_01722_),
    .DE(_00081_),
    .Q(\w[37][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][25]$_SDFFCE_PN0P_  (.D(_01723_),
    .DE(_00081_),
    .Q(\w[37][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][26]$_SDFFCE_PN0P_  (.D(_01724_),
    .DE(_00081_),
    .Q(\w[37][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][27]$_SDFFCE_PN0P_  (.D(_01725_),
    .DE(_00081_),
    .Q(\w[37][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][28]$_SDFFCE_PN0P_  (.D(_01726_),
    .DE(_00081_),
    .Q(\w[37][28] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][29]$_SDFFCE_PN0P_  (.D(_01727_),
    .DE(_00081_),
    .Q(\w[37][29] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][2]$_SDFFCE_PN0P_  (.D(_01728_),
    .DE(_00081_),
    .Q(\w[37][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][30]$_SDFFCE_PN0P_  (.D(_01729_),
    .DE(_00081_),
    .Q(\w[37][30] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][31]$_SDFFCE_PN0P_  (.D(_01730_),
    .DE(_00081_),
    .Q(\w[37][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][3]$_SDFFCE_PN0P_  (.D(_01731_),
    .DE(_00081_),
    .Q(\w[37][3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][4]$_SDFFCE_PN0P_  (.D(_01732_),
    .DE(_00081_),
    .Q(\w[37][4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][5]$_SDFFCE_PN0P_  (.D(_01733_),
    .DE(_00081_),
    .Q(\w[37][5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][6]$_SDFFCE_PN0P_  (.D(_01734_),
    .DE(_00081_),
    .Q(\w[37][6] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][7]$_SDFFCE_PN0P_  (.D(_01735_),
    .DE(_00081_),
    .Q(\w[37][7] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][8]$_SDFFCE_PN0P_  (.D(_01736_),
    .DE(_00081_),
    .Q(\w[37][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][9]$_SDFFCE_PN0P_  (.D(_01737_),
    .DE(_00081_),
    .Q(\w[37][9] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][0]$_SDFFCE_PN0P_  (.D(_01738_),
    .DE(_00111_),
    .Q(\w[38][0] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][10]$_SDFFCE_PN0P_  (.D(_01739_),
    .DE(_00111_),
    .Q(\w[38][10] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][11]$_SDFFCE_PN0P_  (.D(_01740_),
    .DE(_00111_),
    .Q(\w[38][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][12]$_SDFFCE_PN0P_  (.D(_01741_),
    .DE(_00111_),
    .Q(\w[38][12] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][13]$_SDFFCE_PN0P_  (.D(_01742_),
    .DE(_00111_),
    .Q(\w[38][13] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][14]$_SDFFCE_PN0P_  (.D(_01743_),
    .DE(_00111_),
    .Q(\w[38][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][15]$_SDFFCE_PN0P_  (.D(_01744_),
    .DE(_00111_),
    .Q(\w[38][15] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][16]$_SDFFCE_PN0P_  (.D(_01745_),
    .DE(_00111_),
    .Q(\w[38][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][17]$_SDFFCE_PN0P_  (.D(_01746_),
    .DE(_00111_),
    .Q(\w[38][17] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][18]$_SDFFCE_PN0P_  (.D(_01747_),
    .DE(_00111_),
    .Q(\w[38][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][19]$_SDFFCE_PN0P_  (.D(_01748_),
    .DE(_00111_),
    .Q(\w[38][19] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][1]$_SDFFCE_PN0P_  (.D(_01749_),
    .DE(_00111_),
    .Q(\w[38][1] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][20]$_SDFFCE_PN0P_  (.D(_01750_),
    .DE(_00111_),
    .Q(\w[38][20] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][21]$_SDFFCE_PN0P_  (.D(_01751_),
    .DE(_00111_),
    .Q(\w[38][21] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][22]$_SDFFCE_PN0P_  (.D(_01752_),
    .DE(_00111_),
    .Q(\w[38][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][23]$_SDFFCE_PN0P_  (.D(_01753_),
    .DE(_00111_),
    .Q(\w[38][23] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][24]$_SDFFCE_PN0P_  (.D(_01754_),
    .DE(_00111_),
    .Q(\w[38][24] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][25]$_SDFFCE_PN0P_  (.D(_01755_),
    .DE(_00111_),
    .Q(\w[38][25] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][26]$_SDFFCE_PN0P_  (.D(_01756_),
    .DE(_00111_),
    .Q(\w[38][26] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][27]$_SDFFCE_PN0P_  (.D(_01757_),
    .DE(_00111_),
    .Q(\w[38][27] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][28]$_SDFFCE_PN0P_  (.D(_01758_),
    .DE(_00111_),
    .Q(\w[38][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][29]$_SDFFCE_PN0P_  (.D(_01759_),
    .DE(_00111_),
    .Q(\w[38][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][2]$_SDFFCE_PN0P_  (.D(_01760_),
    .DE(_00111_),
    .Q(\w[38][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][30]$_SDFFCE_PN0P_  (.D(_01761_),
    .DE(_00111_),
    .Q(\w[38][30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][31]$_SDFFCE_PN0P_  (.D(_01762_),
    .DE(_00111_),
    .Q(\w[38][31] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][3]$_SDFFCE_PN0P_  (.D(_01763_),
    .DE(_00111_),
    .Q(\w[38][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][4]$_SDFFCE_PN0P_  (.D(_01764_),
    .DE(_00111_),
    .Q(\w[38][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][5]$_SDFFCE_PN0P_  (.D(_01765_),
    .DE(_00111_),
    .Q(\w[38][5] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][6]$_SDFFCE_PN0P_  (.D(_01766_),
    .DE(_00111_),
    .Q(\w[38][6] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][7]$_SDFFCE_PN0P_  (.D(_01767_),
    .DE(_00111_),
    .Q(\w[38][7] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][8]$_SDFFCE_PN0P_  (.D(_01768_),
    .DE(_00111_),
    .Q(\w[38][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][9]$_SDFFCE_PN0P_  (.D(_01769_),
    .DE(_00111_),
    .Q(\w[38][9] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][0]$_SDFFCE_PN0P_  (.D(_01770_),
    .DE(net474),
    .Q(\w[39][0] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][10]$_SDFFCE_PN0P_  (.D(_01771_),
    .DE(net472),
    .Q(\w[39][10] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][11]$_SDFFCE_PN0P_  (.D(_01772_),
    .DE(_00080_),
    .Q(\w[39][11] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][12]$_SDFFCE_PN0P_  (.D(_01773_),
    .DE(net474),
    .Q(\w[39][12] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][13]$_SDFFCE_PN0P_  (.D(_01774_),
    .DE(net472),
    .Q(\w[39][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][14]$_SDFFCE_PN0P_  (.D(_01775_),
    .DE(net473),
    .Q(\w[39][14] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][15]$_SDFFCE_PN0P_  (.D(_01776_),
    .DE(net473),
    .Q(\w[39][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][16]$_SDFFCE_PN0P_  (.D(_01777_),
    .DE(net473),
    .Q(\w[39][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][17]$_SDFFCE_PN0P_  (.D(_01778_),
    .DE(net473),
    .Q(\w[39][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][18]$_SDFFCE_PN0P_  (.D(_01779_),
    .DE(net472),
    .Q(\w[39][18] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][19]$_SDFFCE_PN0P_  (.D(_01780_),
    .DE(_00080_),
    .Q(\w[39][19] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][1]$_SDFFCE_PN0P_  (.D(_01781_),
    .DE(net473),
    .Q(\w[39][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][20]$_SDFFCE_PN0P_  (.D(_01782_),
    .DE(_00080_),
    .Q(\w[39][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][21]$_SDFFCE_PN0P_  (.D(_01783_),
    .DE(net472),
    .Q(\w[39][21] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][22]$_SDFFCE_PN0P_  (.D(_01784_),
    .DE(net472),
    .Q(\w[39][22] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][23]$_SDFFCE_PN0P_  (.D(_01785_),
    .DE(net474),
    .Q(\w[39][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][24]$_SDFFCE_PN0P_  (.D(_01786_),
    .DE(net473),
    .Q(\w[39][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][25]$_SDFFCE_PN0P_  (.D(_01787_),
    .DE(net473),
    .Q(\w[39][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][26]$_SDFFCE_PN0P_  (.D(_01788_),
    .DE(net474),
    .Q(\w[39][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][27]$_SDFFCE_PN0P_  (.D(_01789_),
    .DE(net473),
    .Q(\w[39][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][28]$_SDFFCE_PN0P_  (.D(_01790_),
    .DE(net472),
    .Q(\w[39][28] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][29]$_SDFFCE_PN0P_  (.D(_01791_),
    .DE(net472),
    .Q(\w[39][29] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][2]$_SDFFCE_PN0P_  (.D(_01792_),
    .DE(net473),
    .Q(\w[39][2] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][30]$_SDFFCE_PN0P_  (.D(_01793_),
    .DE(net472),
    .Q(\w[39][30] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][31]$_SDFFCE_PN0P_  (.D(_01794_),
    .DE(net474),
    .Q(\w[39][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][3]$_SDFFCE_PN0P_  (.D(_01795_),
    .DE(net473),
    .Q(\w[39][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][4]$_SDFFCE_PN0P_  (.D(_01796_),
    .DE(net474),
    .Q(\w[39][4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][5]$_SDFFCE_PN0P_  (.D(_01797_),
    .DE(net473),
    .Q(\w[39][5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][6]$_SDFFCE_PN0P_  (.D(_01798_),
    .DE(net472),
    .Q(\w[39][6] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][7]$_SDFFCE_PN0P_  (.D(_01799_),
    .DE(net473),
    .Q(\w[39][7] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][8]$_SDFFCE_PN0P_  (.D(_01800_),
    .DE(net474),
    .Q(\w[39][8] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][9]$_SDFFCE_PN0P_  (.D(_01801_),
    .DE(net472),
    .Q(\w[39][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][0]$_DFFE_PP_  (.D(_00417_),
    .DE(_00079_),
    .Q(\w[3][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][10]$_DFFE_PP_  (.D(_00418_),
    .DE(_00079_),
    .Q(\w[3][10] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][11]$_DFFE_PP_  (.D(_00419_),
    .DE(_00079_),
    .Q(\w[3][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][12]$_DFFE_PP_  (.D(_00420_),
    .DE(_00079_),
    .Q(\w[3][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][13]$_DFFE_PP_  (.D(_00421_),
    .DE(_00079_),
    .Q(\w[3][13] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][14]$_DFFE_PP_  (.D(_00422_),
    .DE(_00079_),
    .Q(\w[3][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][15]$_DFFE_PP_  (.D(_00423_),
    .DE(_00079_),
    .Q(\w[3][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][16]$_DFFE_PP_  (.D(_00424_),
    .DE(_00079_),
    .Q(\w[3][16] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][17]$_DFFE_PP_  (.D(_00425_),
    .DE(_00079_),
    .Q(\w[3][17] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][18]$_DFFE_PP_  (.D(_00426_),
    .DE(_00079_),
    .Q(\w[3][18] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][19]$_DFFE_PP_  (.D(_00427_),
    .DE(_00079_),
    .Q(\w[3][19] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][1]$_DFFE_PP_  (.D(_00428_),
    .DE(_00079_),
    .Q(\w[3][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][20]$_DFFE_PP_  (.D(_00429_),
    .DE(_00079_),
    .Q(\w[3][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][21]$_DFFE_PP_  (.D(_00430_),
    .DE(_00079_),
    .Q(\w[3][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][22]$_DFFE_PP_  (.D(_00431_),
    .DE(_00079_),
    .Q(\w[3][22] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][23]$_DFFE_PP_  (.D(_00432_),
    .DE(_00079_),
    .Q(\w[3][23] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][24]$_DFFE_PP_  (.D(_00433_),
    .DE(_00079_),
    .Q(\w[3][24] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][25]$_DFFE_PP_  (.D(_00434_),
    .DE(_00079_),
    .Q(\w[3][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][26]$_DFFE_PP_  (.D(_00435_),
    .DE(_00079_),
    .Q(\w[3][26] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][27]$_DFFE_PP_  (.D(_00436_),
    .DE(_00079_),
    .Q(\w[3][27] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][28]$_DFFE_PP_  (.D(_00437_),
    .DE(_00079_),
    .Q(\w[3][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][29]$_DFFE_PP_  (.D(_00438_),
    .DE(_00079_),
    .Q(\w[3][29] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][2]$_DFFE_PP_  (.D(_00439_),
    .DE(_00079_),
    .Q(\w[3][2] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][30]$_DFFE_PP_  (.D(_00440_),
    .DE(_00079_),
    .Q(\w[3][30] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][31]$_DFFE_PP_  (.D(_00441_),
    .DE(_00079_),
    .Q(\w[3][31] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][3]$_DFFE_PP_  (.D(_00442_),
    .DE(_00079_),
    .Q(\w[3][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][4]$_DFFE_PP_  (.D(_00443_),
    .DE(_00079_),
    .Q(\w[3][4] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][5]$_DFFE_PP_  (.D(_00444_),
    .DE(_00079_),
    .Q(\w[3][5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][6]$_DFFE_PP_  (.D(_00445_),
    .DE(_00079_),
    .Q(\w[3][6] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][7]$_DFFE_PP_  (.D(_00446_),
    .DE(_00079_),
    .Q(\w[3][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][8]$_DFFE_PP_  (.D(_00447_),
    .DE(_00079_),
    .Q(\w[3][8] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][9]$_DFFE_PP_  (.D(_00448_),
    .DE(_00079_),
    .Q(\w[3][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][0]$_SDFFCE_PN0P_  (.D(_01802_),
    .DE(_00110_),
    .Q(\w[40][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][10]$_SDFFCE_PN0P_  (.D(_01803_),
    .DE(_00110_),
    .Q(\w[40][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][11]$_SDFFCE_PN0P_  (.D(_01804_),
    .DE(_00110_),
    .Q(\w[40][11] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][12]$_SDFFCE_PN0P_  (.D(_01805_),
    .DE(_00110_),
    .Q(\w[40][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][13]$_SDFFCE_PN0P_  (.D(_01806_),
    .DE(_00110_),
    .Q(\w[40][13] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][14]$_SDFFCE_PN0P_  (.D(_01807_),
    .DE(_00110_),
    .Q(\w[40][14] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][15]$_SDFFCE_PN0P_  (.D(_01808_),
    .DE(_00110_),
    .Q(\w[40][15] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][16]$_SDFFCE_PN0P_  (.D(_01809_),
    .DE(_00110_),
    .Q(\w[40][16] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][17]$_SDFFCE_PN0P_  (.D(_01810_),
    .DE(_00110_),
    .Q(\w[40][17] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][18]$_SDFFCE_PN0P_  (.D(_01811_),
    .DE(_00110_),
    .Q(\w[40][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][19]$_SDFFCE_PN0P_  (.D(_01812_),
    .DE(_00110_),
    .Q(\w[40][19] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][1]$_SDFFCE_PN0P_  (.D(_01813_),
    .DE(_00110_),
    .Q(\w[40][1] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][20]$_SDFFCE_PN0P_  (.D(_01814_),
    .DE(_00110_),
    .Q(\w[40][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][21]$_SDFFCE_PN0P_  (.D(_01815_),
    .DE(_00110_),
    .Q(\w[40][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][22]$_SDFFCE_PN0P_  (.D(_01816_),
    .DE(_00110_),
    .Q(\w[40][22] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][23]$_SDFFCE_PN0P_  (.D(_01817_),
    .DE(_00110_),
    .Q(\w[40][23] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][24]$_SDFFCE_PN0P_  (.D(_01818_),
    .DE(_00110_),
    .Q(\w[40][24] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][25]$_SDFFCE_PN0P_  (.D(_01819_),
    .DE(_00110_),
    .Q(\w[40][25] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][26]$_SDFFCE_PN0P_  (.D(_01820_),
    .DE(_00110_),
    .Q(\w[40][26] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][27]$_SDFFCE_PN0P_  (.D(_01821_),
    .DE(_00110_),
    .Q(\w[40][27] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][28]$_SDFFCE_PN0P_  (.D(_01822_),
    .DE(_00110_),
    .Q(\w[40][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][29]$_SDFFCE_PN0P_  (.D(_01823_),
    .DE(_00110_),
    .Q(\w[40][29] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][2]$_SDFFCE_PN0P_  (.D(_01824_),
    .DE(_00110_),
    .Q(\w[40][2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][30]$_SDFFCE_PN0P_  (.D(_01825_),
    .DE(_00110_),
    .Q(\w[40][30] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][31]$_SDFFCE_PN0P_  (.D(_01826_),
    .DE(_00110_),
    .Q(\w[40][31] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][3]$_SDFFCE_PN0P_  (.D(_01827_),
    .DE(_00110_),
    .Q(\w[40][3] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][4]$_SDFFCE_PN0P_  (.D(_01828_),
    .DE(_00110_),
    .Q(\w[40][4] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][5]$_SDFFCE_PN0P_  (.D(_01829_),
    .DE(_00110_),
    .Q(\w[40][5] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][6]$_SDFFCE_PN0P_  (.D(_01830_),
    .DE(_00110_),
    .Q(\w[40][6] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][7]$_SDFFCE_PN0P_  (.D(_01831_),
    .DE(_00110_),
    .Q(\w[40][7] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][8]$_SDFFCE_PN0P_  (.D(_01832_),
    .DE(_00110_),
    .Q(\w[40][8] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][9]$_SDFFCE_PN0P_  (.D(_01833_),
    .DE(_00110_),
    .Q(\w[40][9] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][0]$_SDFFCE_PN0P_  (.D(_01834_),
    .DE(_00078_),
    .Q(\w[41][0] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][10]$_SDFFCE_PN0P_  (.D(_01835_),
    .DE(_00078_),
    .Q(\w[41][10] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][11]$_SDFFCE_PN0P_  (.D(_01836_),
    .DE(_00078_),
    .Q(\w[41][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][12]$_SDFFCE_PN0P_  (.D(_01837_),
    .DE(_00078_),
    .Q(\w[41][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][13]$_SDFFCE_PN0P_  (.D(_01838_),
    .DE(_00078_),
    .Q(\w[41][13] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][14]$_SDFFCE_PN0P_  (.D(_01839_),
    .DE(_00078_),
    .Q(\w[41][14] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][15]$_SDFFCE_PN0P_  (.D(_01840_),
    .DE(_00078_),
    .Q(\w[41][15] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][16]$_SDFFCE_PN0P_  (.D(_01841_),
    .DE(_00078_),
    .Q(\w[41][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][17]$_SDFFCE_PN0P_  (.D(_01842_),
    .DE(_00078_),
    .Q(\w[41][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][18]$_SDFFCE_PN0P_  (.D(_01843_),
    .DE(_00078_),
    .Q(\w[41][18] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][19]$_SDFFCE_PN0P_  (.D(_01844_),
    .DE(_00078_),
    .Q(\w[41][19] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][1]$_SDFFCE_PN0P_  (.D(_01845_),
    .DE(_00078_),
    .Q(\w[41][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][20]$_SDFFCE_PN0P_  (.D(_01846_),
    .DE(_00078_),
    .Q(\w[41][20] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][21]$_SDFFCE_PN0P_  (.D(_01847_),
    .DE(_00078_),
    .Q(\w[41][21] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][22]$_SDFFCE_PN0P_  (.D(_01848_),
    .DE(_00078_),
    .Q(\w[41][22] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][23]$_SDFFCE_PN0P_  (.D(_01849_),
    .DE(_00078_),
    .Q(\w[41][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][24]$_SDFFCE_PN0P_  (.D(_01850_),
    .DE(_00078_),
    .Q(\w[41][24] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][25]$_SDFFCE_PN0P_  (.D(_01851_),
    .DE(_00078_),
    .Q(\w[41][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][26]$_SDFFCE_PN0P_  (.D(_01852_),
    .DE(_00078_),
    .Q(\w[41][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][27]$_SDFFCE_PN0P_  (.D(_01853_),
    .DE(_00078_),
    .Q(\w[41][27] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][28]$_SDFFCE_PN0P_  (.D(_01854_),
    .DE(_00078_),
    .Q(\w[41][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][29]$_SDFFCE_PN0P_  (.D(_01855_),
    .DE(_00078_),
    .Q(\w[41][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][2]$_SDFFCE_PN0P_  (.D(_01856_),
    .DE(_00078_),
    .Q(\w[41][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][30]$_SDFFCE_PN0P_  (.D(_01857_),
    .DE(_00078_),
    .Q(\w[41][30] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][31]$_SDFFCE_PN0P_  (.D(_01858_),
    .DE(_00078_),
    .Q(\w[41][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][3]$_SDFFCE_PN0P_  (.D(_01859_),
    .DE(_00078_),
    .Q(\w[41][3] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][4]$_SDFFCE_PN0P_  (.D(_01860_),
    .DE(_00078_),
    .Q(\w[41][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][5]$_SDFFCE_PN0P_  (.D(_01861_),
    .DE(_00078_),
    .Q(\w[41][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][6]$_SDFFCE_PN0P_  (.D(_01862_),
    .DE(_00078_),
    .Q(\w[41][6] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][7]$_SDFFCE_PN0P_  (.D(_01863_),
    .DE(_00078_),
    .Q(\w[41][7] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][8]$_SDFFCE_PN0P_  (.D(_01864_),
    .DE(_00078_),
    .Q(\w[41][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][9]$_SDFFCE_PN0P_  (.D(_01865_),
    .DE(_00078_),
    .Q(\w[41][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][0]$_SDFFCE_PN0P_  (.D(_01866_),
    .DE(_00109_),
    .Q(\w[42][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][10]$_SDFFCE_PN0P_  (.D(_01867_),
    .DE(_00109_),
    .Q(\w[42][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][11]$_SDFFCE_PN0P_  (.D(_01868_),
    .DE(_00109_),
    .Q(\w[42][11] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][12]$_SDFFCE_PN0P_  (.D(_01869_),
    .DE(_00109_),
    .Q(\w[42][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][13]$_SDFFCE_PN0P_  (.D(_01870_),
    .DE(_00109_),
    .Q(\w[42][13] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][14]$_SDFFCE_PN0P_  (.D(_01871_),
    .DE(_00109_),
    .Q(\w[42][14] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][15]$_SDFFCE_PN0P_  (.D(_01872_),
    .DE(_00109_),
    .Q(\w[42][15] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][16]$_SDFFCE_PN0P_  (.D(_01873_),
    .DE(_00109_),
    .Q(\w[42][16] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][17]$_SDFFCE_PN0P_  (.D(_01874_),
    .DE(_00109_),
    .Q(\w[42][17] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][18]$_SDFFCE_PN0P_  (.D(_01875_),
    .DE(_00109_),
    .Q(\w[42][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][19]$_SDFFCE_PN0P_  (.D(_01876_),
    .DE(_00109_),
    .Q(\w[42][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][1]$_SDFFCE_PN0P_  (.D(_01877_),
    .DE(_00109_),
    .Q(\w[42][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][20]$_SDFFCE_PN0P_  (.D(_01878_),
    .DE(_00109_),
    .Q(\w[42][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][21]$_SDFFCE_PN0P_  (.D(_01879_),
    .DE(_00109_),
    .Q(\w[42][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][22]$_SDFFCE_PN0P_  (.D(_01880_),
    .DE(_00109_),
    .Q(\w[42][22] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][23]$_SDFFCE_PN0P_  (.D(_01881_),
    .DE(_00109_),
    .Q(\w[42][23] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][24]$_SDFFCE_PN0P_  (.D(_01882_),
    .DE(_00109_),
    .Q(\w[42][24] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][25]$_SDFFCE_PN0P_  (.D(_01883_),
    .DE(_00109_),
    .Q(\w[42][25] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][26]$_SDFFCE_PN0P_  (.D(_01884_),
    .DE(_00109_),
    .Q(\w[42][26] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][27]$_SDFFCE_PN0P_  (.D(_01885_),
    .DE(_00109_),
    .Q(\w[42][27] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][28]$_SDFFCE_PN0P_  (.D(_01886_),
    .DE(_00109_),
    .Q(\w[42][28] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][29]$_SDFFCE_PN0P_  (.D(_01887_),
    .DE(_00109_),
    .Q(\w[42][29] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][2]$_SDFFCE_PN0P_  (.D(_01888_),
    .DE(_00109_),
    .Q(\w[42][2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][30]$_SDFFCE_PN0P_  (.D(_01889_),
    .DE(_00109_),
    .Q(\w[42][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][31]$_SDFFCE_PN0P_  (.D(_01890_),
    .DE(_00109_),
    .Q(\w[42][31] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][3]$_SDFFCE_PN0P_  (.D(_01891_),
    .DE(_00109_),
    .Q(\w[42][3] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][4]$_SDFFCE_PN0P_  (.D(_01892_),
    .DE(_00109_),
    .Q(\w[42][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][5]$_SDFFCE_PN0P_  (.D(_01893_),
    .DE(_00109_),
    .Q(\w[42][5] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][6]$_SDFFCE_PN0P_  (.D(_01894_),
    .DE(_00109_),
    .Q(\w[42][6] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][7]$_SDFFCE_PN0P_  (.D(_01895_),
    .DE(_00109_),
    .Q(\w[42][7] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][8]$_SDFFCE_PN0P_  (.D(_01896_),
    .DE(_00109_),
    .Q(\w[42][8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][9]$_SDFFCE_PN0P_  (.D(_01897_),
    .DE(_00109_),
    .Q(\w[42][9] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][0]$_SDFFCE_PN0P_  (.D(_01898_),
    .DE(_00077_),
    .Q(\w[43][0] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][10]$_SDFFCE_PN0P_  (.D(_01899_),
    .DE(_00077_),
    .Q(\w[43][10] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][11]$_SDFFCE_PN0P_  (.D(_01900_),
    .DE(_00077_),
    .Q(\w[43][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][12]$_SDFFCE_PN0P_  (.D(_01901_),
    .DE(_00077_),
    .Q(\w[43][12] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][13]$_SDFFCE_PN0P_  (.D(_01902_),
    .DE(_00077_),
    .Q(\w[43][13] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][14]$_SDFFCE_PN0P_  (.D(_01903_),
    .DE(_00077_),
    .Q(\w[43][14] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][15]$_SDFFCE_PN0P_  (.D(_01904_),
    .DE(_00077_),
    .Q(\w[43][15] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][16]$_SDFFCE_PN0P_  (.D(_01905_),
    .DE(_00077_),
    .Q(\w[43][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][17]$_SDFFCE_PN0P_  (.D(_01906_),
    .DE(_00077_),
    .Q(\w[43][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][18]$_SDFFCE_PN0P_  (.D(_01907_),
    .DE(_00077_),
    .Q(\w[43][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][19]$_SDFFCE_PN0P_  (.D(_01908_),
    .DE(_00077_),
    .Q(\w[43][19] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][1]$_SDFFCE_PN0P_  (.D(_01909_),
    .DE(_00077_),
    .Q(\w[43][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][20]$_SDFFCE_PN0P_  (.D(_01910_),
    .DE(_00077_),
    .Q(\w[43][20] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][21]$_SDFFCE_PN0P_  (.D(_01911_),
    .DE(_00077_),
    .Q(\w[43][21] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][22]$_SDFFCE_PN0P_  (.D(_01912_),
    .DE(_00077_),
    .Q(\w[43][22] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][23]$_SDFFCE_PN0P_  (.D(_01913_),
    .DE(_00077_),
    .Q(\w[43][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][24]$_SDFFCE_PN0P_  (.D(_01914_),
    .DE(_00077_),
    .Q(\w[43][24] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][25]$_SDFFCE_PN0P_  (.D(_01915_),
    .DE(_00077_),
    .Q(\w[43][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][26]$_SDFFCE_PN0P_  (.D(_01916_),
    .DE(_00077_),
    .Q(\w[43][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][27]$_SDFFCE_PN0P_  (.D(_01917_),
    .DE(_00077_),
    .Q(\w[43][27] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][28]$_SDFFCE_PN0P_  (.D(_01918_),
    .DE(_00077_),
    .Q(\w[43][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][29]$_SDFFCE_PN0P_  (.D(_01919_),
    .DE(_00077_),
    .Q(\w[43][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][2]$_SDFFCE_PN0P_  (.D(_01920_),
    .DE(_00077_),
    .Q(\w[43][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][30]$_SDFFCE_PN0P_  (.D(_01921_),
    .DE(_00077_),
    .Q(\w[43][30] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][31]$_SDFFCE_PN0P_  (.D(_01922_),
    .DE(_00077_),
    .Q(\w[43][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][3]$_SDFFCE_PN0P_  (.D(_01923_),
    .DE(_00077_),
    .Q(\w[43][3] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][4]$_SDFFCE_PN0P_  (.D(_01924_),
    .DE(_00077_),
    .Q(\w[43][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][5]$_SDFFCE_PN0P_  (.D(_01925_),
    .DE(_00077_),
    .Q(\w[43][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][6]$_SDFFCE_PN0P_  (.D(_01926_),
    .DE(_00077_),
    .Q(\w[43][6] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][7]$_SDFFCE_PN0P_  (.D(_01927_),
    .DE(_00077_),
    .Q(\w[43][7] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][8]$_SDFFCE_PN0P_  (.D(_01928_),
    .DE(_00077_),
    .Q(\w[43][8] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][9]$_SDFFCE_PN0P_  (.D(_01929_),
    .DE(_00077_),
    .Q(\w[43][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][0]$_SDFFCE_PN0P_  (.D(_01930_),
    .DE(_00108_),
    .Q(\w[44][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][10]$_SDFFCE_PN0P_  (.D(_01931_),
    .DE(_00108_),
    .Q(\w[44][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][11]$_SDFFCE_PN0P_  (.D(_01932_),
    .DE(_00108_),
    .Q(\w[44][11] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][12]$_SDFFCE_PN0P_  (.D(_01933_),
    .DE(_00108_),
    .Q(\w[44][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][13]$_SDFFCE_PN0P_  (.D(_01934_),
    .DE(_00108_),
    .Q(\w[44][13] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][14]$_SDFFCE_PN0P_  (.D(_01935_),
    .DE(_00108_),
    .Q(\w[44][14] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][15]$_SDFFCE_PN0P_  (.D(_01936_),
    .DE(_00108_),
    .Q(\w[44][15] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][16]$_SDFFCE_PN0P_  (.D(_01937_),
    .DE(_00108_),
    .Q(\w[44][16] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][17]$_SDFFCE_PN0P_  (.D(_01938_),
    .DE(_00108_),
    .Q(\w[44][17] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][18]$_SDFFCE_PN0P_  (.D(_01939_),
    .DE(_00108_),
    .Q(\w[44][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][19]$_SDFFCE_PN0P_  (.D(_01940_),
    .DE(_00108_),
    .Q(\w[44][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][1]$_SDFFCE_PN0P_  (.D(_01941_),
    .DE(_00108_),
    .Q(\w[44][1] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][20]$_SDFFCE_PN0P_  (.D(_01942_),
    .DE(_00108_),
    .Q(\w[44][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][21]$_SDFFCE_PN0P_  (.D(_01943_),
    .DE(_00108_),
    .Q(\w[44][21] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][22]$_SDFFCE_PN0P_  (.D(_01944_),
    .DE(_00108_),
    .Q(\w[44][22] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][23]$_SDFFCE_PN0P_  (.D(_01945_),
    .DE(_00108_),
    .Q(\w[44][23] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][24]$_SDFFCE_PN0P_  (.D(_01946_),
    .DE(_00108_),
    .Q(\w[44][24] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][25]$_SDFFCE_PN0P_  (.D(_01947_),
    .DE(_00108_),
    .Q(\w[44][25] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][26]$_SDFFCE_PN0P_  (.D(_01948_),
    .DE(_00108_),
    .Q(\w[44][26] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][27]$_SDFFCE_PN0P_  (.D(_01949_),
    .DE(_00108_),
    .Q(\w[44][27] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][28]$_SDFFCE_PN0P_  (.D(_01950_),
    .DE(_00108_),
    .Q(\w[44][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][29]$_SDFFCE_PN0P_  (.D(_01951_),
    .DE(_00108_),
    .Q(\w[44][29] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][2]$_SDFFCE_PN0P_  (.D(_01952_),
    .DE(_00108_),
    .Q(\w[44][2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][30]$_SDFFCE_PN0P_  (.D(_01953_),
    .DE(_00108_),
    .Q(\w[44][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][31]$_SDFFCE_PN0P_  (.D(_01954_),
    .DE(_00108_),
    .Q(\w[44][31] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][3]$_SDFFCE_PN0P_  (.D(_01955_),
    .DE(_00108_),
    .Q(\w[44][3] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][4]$_SDFFCE_PN0P_  (.D(_01956_),
    .DE(_00108_),
    .Q(\w[44][4] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][5]$_SDFFCE_PN0P_  (.D(_01957_),
    .DE(_00108_),
    .Q(\w[44][5] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][6]$_SDFFCE_PN0P_  (.D(_01958_),
    .DE(_00108_),
    .Q(\w[44][6] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][7]$_SDFFCE_PN0P_  (.D(_01959_),
    .DE(_00108_),
    .Q(\w[44][7] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][8]$_SDFFCE_PN0P_  (.D(_01960_),
    .DE(_00108_),
    .Q(\w[44][8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][9]$_SDFFCE_PN0P_  (.D(_01961_),
    .DE(_00108_),
    .Q(\w[44][9] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][0]$_SDFFCE_PN0P_  (.D(_01962_),
    .DE(_00076_),
    .Q(\w[45][0] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][10]$_SDFFCE_PN0P_  (.D(_01963_),
    .DE(_00076_),
    .Q(\w[45][10] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][11]$_SDFFCE_PN0P_  (.D(_01964_),
    .DE(_00076_),
    .Q(\w[45][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][12]$_SDFFCE_PN0P_  (.D(_01965_),
    .DE(_00076_),
    .Q(\w[45][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][13]$_SDFFCE_PN0P_  (.D(_01966_),
    .DE(_00076_),
    .Q(\w[45][13] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][14]$_SDFFCE_PN0P_  (.D(_01967_),
    .DE(_00076_),
    .Q(\w[45][14] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][15]$_SDFFCE_PN0P_  (.D(_01968_),
    .DE(_00076_),
    .Q(\w[45][15] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][16]$_SDFFCE_PN0P_  (.D(_01969_),
    .DE(_00076_),
    .Q(\w[45][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][17]$_SDFFCE_PN0P_  (.D(_01970_),
    .DE(_00076_),
    .Q(\w[45][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][18]$_SDFFCE_PN0P_  (.D(_01971_),
    .DE(_00076_),
    .Q(\w[45][18] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][19]$_SDFFCE_PN0P_  (.D(_01972_),
    .DE(_00076_),
    .Q(\w[45][19] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][1]$_SDFFCE_PN0P_  (.D(_01973_),
    .DE(_00076_),
    .Q(\w[45][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][20]$_SDFFCE_PN0P_  (.D(_01974_),
    .DE(_00076_),
    .Q(\w[45][20] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][21]$_SDFFCE_PN0P_  (.D(_01975_),
    .DE(_00076_),
    .Q(\w[45][21] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][22]$_SDFFCE_PN0P_  (.D(_01976_),
    .DE(_00076_),
    .Q(\w[45][22] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][23]$_SDFFCE_PN0P_  (.D(_01977_),
    .DE(_00076_),
    .Q(\w[45][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][24]$_SDFFCE_PN0P_  (.D(_01978_),
    .DE(_00076_),
    .Q(\w[45][24] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][25]$_SDFFCE_PN0P_  (.D(_01979_),
    .DE(_00076_),
    .Q(\w[45][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][26]$_SDFFCE_PN0P_  (.D(_01980_),
    .DE(_00076_),
    .Q(\w[45][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][27]$_SDFFCE_PN0P_  (.D(_01981_),
    .DE(_00076_),
    .Q(\w[45][27] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][28]$_SDFFCE_PN0P_  (.D(_01982_),
    .DE(_00076_),
    .Q(\w[45][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][29]$_SDFFCE_PN0P_  (.D(_01983_),
    .DE(_00076_),
    .Q(\w[45][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][2]$_SDFFCE_PN0P_  (.D(_01984_),
    .DE(_00076_),
    .Q(\w[45][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][30]$_SDFFCE_PN0P_  (.D(_01985_),
    .DE(_00076_),
    .Q(\w[45][30] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][31]$_SDFFCE_PN0P_  (.D(_01986_),
    .DE(_00076_),
    .Q(\w[45][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][3]$_SDFFCE_PN0P_  (.D(_01987_),
    .DE(_00076_),
    .Q(\w[45][3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][4]$_SDFFCE_PN0P_  (.D(_01988_),
    .DE(_00076_),
    .Q(\w[45][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][5]$_SDFFCE_PN0P_  (.D(_01989_),
    .DE(_00076_),
    .Q(\w[45][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][6]$_SDFFCE_PN0P_  (.D(_01990_),
    .DE(_00076_),
    .Q(\w[45][6] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][7]$_SDFFCE_PN0P_  (.D(_01991_),
    .DE(_00076_),
    .Q(\w[45][7] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][8]$_SDFFCE_PN0P_  (.D(_01992_),
    .DE(_00076_),
    .Q(\w[45][8] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][9]$_SDFFCE_PN0P_  (.D(_01993_),
    .DE(_00076_),
    .Q(\w[45][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][0]$_SDFFCE_PN0P_  (.D(_01994_),
    .DE(_00107_),
    .Q(\w[46][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][10]$_SDFFCE_PN0P_  (.D(_01995_),
    .DE(_00107_),
    .Q(\w[46][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][11]$_SDFFCE_PN0P_  (.D(_01996_),
    .DE(_00107_),
    .Q(\w[46][11] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][12]$_SDFFCE_PN0P_  (.D(_01997_),
    .DE(_00107_),
    .Q(\w[46][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][13]$_SDFFCE_PN0P_  (.D(_01998_),
    .DE(_00107_),
    .Q(\w[46][13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][14]$_SDFFCE_PN0P_  (.D(_01999_),
    .DE(_00107_),
    .Q(\w[46][14] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][15]$_SDFFCE_PN0P_  (.D(_02000_),
    .DE(_00107_),
    .Q(\w[46][15] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][16]$_SDFFCE_PN0P_  (.D(_02001_),
    .DE(_00107_),
    .Q(\w[46][16] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][17]$_SDFFCE_PN0P_  (.D(_02002_),
    .DE(_00107_),
    .Q(\w[46][17] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][18]$_SDFFCE_PN0P_  (.D(_02003_),
    .DE(_00107_),
    .Q(\w[46][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][19]$_SDFFCE_PN0P_  (.D(_02004_),
    .DE(_00107_),
    .Q(\w[46][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][1]$_SDFFCE_PN0P_  (.D(_02005_),
    .DE(_00107_),
    .Q(\w[46][1] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][20]$_SDFFCE_PN0P_  (.D(_02006_),
    .DE(_00107_),
    .Q(\w[46][20] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][21]$_SDFFCE_PN0P_  (.D(_02007_),
    .DE(_00107_),
    .Q(\w[46][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][22]$_SDFFCE_PN0P_  (.D(_02008_),
    .DE(_00107_),
    .Q(\w[46][22] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][23]$_SDFFCE_PN0P_  (.D(_02009_),
    .DE(_00107_),
    .Q(\w[46][23] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][24]$_SDFFCE_PN0P_  (.D(_02010_),
    .DE(_00107_),
    .Q(\w[46][24] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][25]$_SDFFCE_PN0P_  (.D(_02011_),
    .DE(_00107_),
    .Q(\w[46][25] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][26]$_SDFFCE_PN0P_  (.D(_02012_),
    .DE(_00107_),
    .Q(\w[46][26] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][27]$_SDFFCE_PN0P_  (.D(_02013_),
    .DE(_00107_),
    .Q(\w[46][27] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][28]$_SDFFCE_PN0P_  (.D(_02014_),
    .DE(_00107_),
    .Q(\w[46][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][29]$_SDFFCE_PN0P_  (.D(_02015_),
    .DE(_00107_),
    .Q(\w[46][29] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][2]$_SDFFCE_PN0P_  (.D(_02016_),
    .DE(_00107_),
    .Q(\w[46][2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][30]$_SDFFCE_PN0P_  (.D(_02017_),
    .DE(_00107_),
    .Q(\w[46][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][31]$_SDFFCE_PN0P_  (.D(_02018_),
    .DE(_00107_),
    .Q(\w[46][31] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][3]$_SDFFCE_PN0P_  (.D(_02019_),
    .DE(_00107_),
    .Q(\w[46][3] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][4]$_SDFFCE_PN0P_  (.D(_02020_),
    .DE(_00107_),
    .Q(\w[46][4] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][5]$_SDFFCE_PN0P_  (.D(_02021_),
    .DE(_00107_),
    .Q(\w[46][5] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][6]$_SDFFCE_PN0P_  (.D(_02022_),
    .DE(_00107_),
    .Q(\w[46][6] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][7]$_SDFFCE_PN0P_  (.D(_02023_),
    .DE(_00107_),
    .Q(\w[46][7] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][8]$_SDFFCE_PN0P_  (.D(_02024_),
    .DE(_00107_),
    .Q(\w[46][8] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][9]$_SDFFCE_PN0P_  (.D(_02025_),
    .DE(_00107_),
    .Q(\w[46][9] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][0]$_SDFFCE_PN0P_  (.D(_02026_),
    .DE(_00075_),
    .Q(\w[47][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][10]$_SDFFCE_PN0P_  (.D(_02027_),
    .DE(_00075_),
    .Q(\w[47][10] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][11]$_SDFFCE_PN0P_  (.D(_02028_),
    .DE(_00075_),
    .Q(\w[47][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][12]$_SDFFCE_PN0P_  (.D(_02029_),
    .DE(_00075_),
    .Q(\w[47][12] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][13]$_SDFFCE_PN0P_  (.D(_02030_),
    .DE(_00075_),
    .Q(\w[47][13] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][14]$_SDFFCE_PN0P_  (.D(_02031_),
    .DE(_00075_),
    .Q(\w[47][14] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][15]$_SDFFCE_PN0P_  (.D(_02032_),
    .DE(_00075_),
    .Q(\w[47][15] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][16]$_SDFFCE_PN0P_  (.D(_02033_),
    .DE(_00075_),
    .Q(\w[47][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][17]$_SDFFCE_PN0P_  (.D(_02034_),
    .DE(_00075_),
    .Q(\w[47][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][18]$_SDFFCE_PN0P_  (.D(_02035_),
    .DE(_00075_),
    .Q(\w[47][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][19]$_SDFFCE_PN0P_  (.D(_02036_),
    .DE(_00075_),
    .Q(\w[47][19] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][1]$_SDFFCE_PN0P_  (.D(_02037_),
    .DE(_00075_),
    .Q(\w[47][1] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][20]$_SDFFCE_PN0P_  (.D(_02038_),
    .DE(_00075_),
    .Q(\w[47][20] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][21]$_SDFFCE_PN0P_  (.D(_02039_),
    .DE(_00075_),
    .Q(\w[47][21] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][22]$_SDFFCE_PN0P_  (.D(_02040_),
    .DE(_00075_),
    .Q(\w[47][22] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][23]$_SDFFCE_PN0P_  (.D(_02041_),
    .DE(_00075_),
    .Q(\w[47][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][24]$_SDFFCE_PN0P_  (.D(_02042_),
    .DE(_00075_),
    .Q(\w[47][24] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][25]$_SDFFCE_PN0P_  (.D(_02043_),
    .DE(_00075_),
    .Q(\w[47][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][26]$_SDFFCE_PN0P_  (.D(_02044_),
    .DE(_00075_),
    .Q(\w[47][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][27]$_SDFFCE_PN0P_  (.D(_02045_),
    .DE(_00075_),
    .Q(\w[47][27] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][28]$_SDFFCE_PN0P_  (.D(_02046_),
    .DE(_00075_),
    .Q(\w[47][28] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][29]$_SDFFCE_PN0P_  (.D(_02047_),
    .DE(_00075_),
    .Q(\w[47][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][2]$_SDFFCE_PN0P_  (.D(_02048_),
    .DE(_00075_),
    .Q(\w[47][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][30]$_SDFFCE_PN0P_  (.D(_02049_),
    .DE(_00075_),
    .Q(\w[47][30] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][31]$_SDFFCE_PN0P_  (.D(_02050_),
    .DE(_00075_),
    .Q(\w[47][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][3]$_SDFFCE_PN0P_  (.D(_02051_),
    .DE(_00075_),
    .Q(\w[47][3] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][4]$_SDFFCE_PN0P_  (.D(_02052_),
    .DE(_00075_),
    .Q(\w[47][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][5]$_SDFFCE_PN0P_  (.D(_02053_),
    .DE(_00075_),
    .Q(\w[47][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][6]$_SDFFCE_PN0P_  (.D(_02054_),
    .DE(_00075_),
    .Q(\w[47][6] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][7]$_SDFFCE_PN0P_  (.D(_02055_),
    .DE(_00075_),
    .Q(\w[47][7] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][8]$_SDFFCE_PN0P_  (.D(_02056_),
    .DE(_00075_),
    .Q(\w[47][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][9]$_SDFFCE_PN0P_  (.D(_02057_),
    .DE(_00075_),
    .Q(\w[47][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][0]$_SDFFCE_PN0P_  (.D(_02058_),
    .DE(_00106_),
    .Q(\w[48][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][10]$_SDFFCE_PN0P_  (.D(_02059_),
    .DE(_00106_),
    .Q(\w[48][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][11]$_SDFFCE_PN0P_  (.D(_02060_),
    .DE(_00106_),
    .Q(\w[48][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][12]$_SDFFCE_PN0P_  (.D(_02061_),
    .DE(_00106_),
    .Q(\w[48][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][13]$_SDFFCE_PN0P_  (.D(_02062_),
    .DE(_00106_),
    .Q(\w[48][13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][14]$_SDFFCE_PN0P_  (.D(_02063_),
    .DE(_00106_),
    .Q(\w[48][14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][15]$_SDFFCE_PN0P_  (.D(_02064_),
    .DE(_00106_),
    .Q(\w[48][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][16]$_SDFFCE_PN0P_  (.D(_02065_),
    .DE(_00106_),
    .Q(\w[48][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][17]$_SDFFCE_PN0P_  (.D(_02066_),
    .DE(_00106_),
    .Q(\w[48][17] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][18]$_SDFFCE_PN0P_  (.D(_02067_),
    .DE(_00106_),
    .Q(\w[48][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][19]$_SDFFCE_PN0P_  (.D(_02068_),
    .DE(_00106_),
    .Q(\w[48][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][1]$_SDFFCE_PN0P_  (.D(_02069_),
    .DE(_00106_),
    .Q(\w[48][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][20]$_SDFFCE_PN0P_  (.D(_02070_),
    .DE(_00106_),
    .Q(\w[48][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][21]$_SDFFCE_PN0P_  (.D(_02071_),
    .DE(_00106_),
    .Q(\w[48][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][22]$_SDFFCE_PN0P_  (.D(_02072_),
    .DE(_00106_),
    .Q(\w[48][22] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][23]$_SDFFCE_PN0P_  (.D(_02073_),
    .DE(_00106_),
    .Q(\w[48][23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][24]$_SDFFCE_PN0P_  (.D(_02074_),
    .DE(_00106_),
    .Q(\w[48][24] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][25]$_SDFFCE_PN0P_  (.D(_02075_),
    .DE(_00106_),
    .Q(\w[48][25] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][26]$_SDFFCE_PN0P_  (.D(_02076_),
    .DE(_00106_),
    .Q(\w[48][26] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][27]$_SDFFCE_PN0P_  (.D(_02077_),
    .DE(_00106_),
    .Q(\w[48][27] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][28]$_SDFFCE_PN0P_  (.D(_02078_),
    .DE(_00106_),
    .Q(\w[48][28] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][29]$_SDFFCE_PN0P_  (.D(_02079_),
    .DE(_00106_),
    .Q(\w[48][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][2]$_SDFFCE_PN0P_  (.D(_02080_),
    .DE(_00106_),
    .Q(\w[48][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][30]$_SDFFCE_PN0P_  (.D(_02081_),
    .DE(_00106_),
    .Q(\w[48][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][31]$_SDFFCE_PN0P_  (.D(_02082_),
    .DE(_00106_),
    .Q(\w[48][31] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][3]$_SDFFCE_PN0P_  (.D(_02083_),
    .DE(_00106_),
    .Q(\w[48][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][4]$_SDFFCE_PN0P_  (.D(_02084_),
    .DE(_00106_),
    .Q(\w[48][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][5]$_SDFFCE_PN0P_  (.D(_02085_),
    .DE(_00106_),
    .Q(\w[48][5] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][6]$_SDFFCE_PN0P_  (.D(_02086_),
    .DE(_00106_),
    .Q(\w[48][6] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][7]$_SDFFCE_PN0P_  (.D(_02087_),
    .DE(_00106_),
    .Q(\w[48][7] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][8]$_SDFFCE_PN0P_  (.D(_02088_),
    .DE(_00106_),
    .Q(\w[48][8] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][9]$_SDFFCE_PN0P_  (.D(_02089_),
    .DE(_00106_),
    .Q(\w[48][9] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][0]$_SDFFCE_PN0P_  (.D(_02090_),
    .DE(_00074_),
    .Q(\w[49][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][10]$_SDFFCE_PN0P_  (.D(_02091_),
    .DE(_00074_),
    .Q(\w[49][10] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][11]$_SDFFCE_PN0P_  (.D(_02092_),
    .DE(_00074_),
    .Q(\w[49][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][12]$_SDFFCE_PN0P_  (.D(_02093_),
    .DE(_00074_),
    .Q(\w[49][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][13]$_SDFFCE_PN0P_  (.D(_02094_),
    .DE(_00074_),
    .Q(\w[49][13] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][14]$_SDFFCE_PN0P_  (.D(_02095_),
    .DE(_00074_),
    .Q(\w[49][14] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][15]$_SDFFCE_PN0P_  (.D(_02096_),
    .DE(_00074_),
    .Q(\w[49][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][16]$_SDFFCE_PN0P_  (.D(_02097_),
    .DE(_00074_),
    .Q(\w[49][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][17]$_SDFFCE_PN0P_  (.D(_02098_),
    .DE(_00074_),
    .Q(\w[49][17] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][18]$_SDFFCE_PN0P_  (.D(_02099_),
    .DE(_00074_),
    .Q(\w[49][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][19]$_SDFFCE_PN0P_  (.D(_02100_),
    .DE(_00074_),
    .Q(\w[49][19] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][1]$_SDFFCE_PN0P_  (.D(_02101_),
    .DE(_00074_),
    .Q(\w[49][1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][20]$_SDFFCE_PN0P_  (.D(_02102_),
    .DE(_00074_),
    .Q(\w[49][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][21]$_SDFFCE_PN0P_  (.D(_02103_),
    .DE(_00074_),
    .Q(\w[49][21] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][22]$_SDFFCE_PN0P_  (.D(_02104_),
    .DE(_00074_),
    .Q(\w[49][22] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][23]$_SDFFCE_PN0P_  (.D(_02105_),
    .DE(_00074_),
    .Q(\w[49][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][24]$_SDFFCE_PN0P_  (.D(_02106_),
    .DE(_00074_),
    .Q(\w[49][24] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][25]$_SDFFCE_PN0P_  (.D(_02107_),
    .DE(_00074_),
    .Q(\w[49][25] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][26]$_SDFFCE_PN0P_  (.D(_02108_),
    .DE(_00074_),
    .Q(\w[49][26] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][27]$_SDFFCE_PN0P_  (.D(_02109_),
    .DE(_00074_),
    .Q(\w[49][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][28]$_SDFFCE_PN0P_  (.D(_02110_),
    .DE(_00074_),
    .Q(\w[49][28] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][29]$_SDFFCE_PN0P_  (.D(_02111_),
    .DE(_00074_),
    .Q(\w[49][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][2]$_SDFFCE_PN0P_  (.D(_02112_),
    .DE(_00074_),
    .Q(\w[49][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][30]$_SDFFCE_PN0P_  (.D(_02113_),
    .DE(_00074_),
    .Q(\w[49][30] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][31]$_SDFFCE_PN0P_  (.D(_02114_),
    .DE(_00074_),
    .Q(\w[49][31] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][3]$_SDFFCE_PN0P_  (.D(_02115_),
    .DE(_00074_),
    .Q(\w[49][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][4]$_SDFFCE_PN0P_  (.D(_02116_),
    .DE(_00074_),
    .Q(\w[49][4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][5]$_SDFFCE_PN0P_  (.D(_02117_),
    .DE(_00074_),
    .Q(\w[49][5] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][6]$_SDFFCE_PN0P_  (.D(_02118_),
    .DE(_00074_),
    .Q(\w[49][6] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][7]$_SDFFCE_PN0P_  (.D(_02119_),
    .DE(_00074_),
    .Q(\w[49][7] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][8]$_SDFFCE_PN0P_  (.D(_02120_),
    .DE(_00074_),
    .Q(\w[49][8] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][9]$_SDFFCE_PN0P_  (.D(_02121_),
    .DE(_00074_),
    .Q(\w[49][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][0]$_DFFE_PP_  (.D(_00449_),
    .DE(_00105_),
    .Q(\w[4][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][10]$_DFFE_PP_  (.D(_00450_),
    .DE(_00105_),
    .Q(\w[4][10] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][11]$_DFFE_PP_  (.D(_00451_),
    .DE(_00105_),
    .Q(\w[4][11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][12]$_DFFE_PP_  (.D(_00452_),
    .DE(_00105_),
    .Q(\w[4][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][13]$_DFFE_PP_  (.D(_00453_),
    .DE(_00105_),
    .Q(\w[4][13] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][14]$_DFFE_PP_  (.D(_00454_),
    .DE(_00105_),
    .Q(\w[4][14] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][15]$_DFFE_PP_  (.D(_00455_),
    .DE(_00105_),
    .Q(\w[4][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][16]$_DFFE_PP_  (.D(_00456_),
    .DE(_00105_),
    .Q(\w[4][16] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][17]$_DFFE_PP_  (.D(_00457_),
    .DE(_00105_),
    .Q(\w[4][17] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][18]$_DFFE_PP_  (.D(_00458_),
    .DE(_00105_),
    .Q(\w[4][18] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][19]$_DFFE_PP_  (.D(_00459_),
    .DE(_00105_),
    .Q(\w[4][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][1]$_DFFE_PP_  (.D(_00460_),
    .DE(_00105_),
    .Q(\w[4][1] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][20]$_DFFE_PP_  (.D(_00461_),
    .DE(_00105_),
    .Q(\w[4][20] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][21]$_DFFE_PP_  (.D(_00462_),
    .DE(_00105_),
    .Q(\w[4][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][22]$_DFFE_PP_  (.D(_00463_),
    .DE(_00105_),
    .Q(\w[4][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][23]$_DFFE_PP_  (.D(_00464_),
    .DE(_00105_),
    .Q(\w[4][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][24]$_DFFE_PP_  (.D(_00465_),
    .DE(_00105_),
    .Q(\w[4][24] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][25]$_DFFE_PP_  (.D(_00466_),
    .DE(_00105_),
    .Q(\w[4][25] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][26]$_DFFE_PP_  (.D(_00467_),
    .DE(_00105_),
    .Q(\w[4][26] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][27]$_DFFE_PP_  (.D(_00468_),
    .DE(_00105_),
    .Q(\w[4][27] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][28]$_DFFE_PP_  (.D(_00469_),
    .DE(_00105_),
    .Q(\w[4][28] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][29]$_DFFE_PP_  (.D(_00470_),
    .DE(_00105_),
    .Q(\w[4][29] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][2]$_DFFE_PP_  (.D(_00471_),
    .DE(_00105_),
    .Q(\w[4][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][30]$_DFFE_PP_  (.D(_00472_),
    .DE(_00105_),
    .Q(\w[4][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][31]$_DFFE_PP_  (.D(_00473_),
    .DE(_00105_),
    .Q(\w[4][31] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][3]$_DFFE_PP_  (.D(_00474_),
    .DE(_00105_),
    .Q(\w[4][3] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][4]$_DFFE_PP_  (.D(_00475_),
    .DE(_00105_),
    .Q(\w[4][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][5]$_DFFE_PP_  (.D(_00476_),
    .DE(_00105_),
    .Q(\w[4][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][6]$_DFFE_PP_  (.D(_00477_),
    .DE(_00105_),
    .Q(\w[4][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][7]$_DFFE_PP_  (.D(_00478_),
    .DE(_00105_),
    .Q(\w[4][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][8]$_DFFE_PP_  (.D(_00479_),
    .DE(_00105_),
    .Q(\w[4][8] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][9]$_DFFE_PP_  (.D(_00480_),
    .DE(_00105_),
    .Q(\w[4][9] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][0]$_SDFFCE_PN0P_  (.D(_02122_),
    .DE(_00104_),
    .Q(\w[50][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][10]$_SDFFCE_PN0P_  (.D(_02123_),
    .DE(_00104_),
    .Q(\w[50][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][11]$_SDFFCE_PN0P_  (.D(_02124_),
    .DE(_00104_),
    .Q(\w[50][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][12]$_SDFFCE_PN0P_  (.D(_02125_),
    .DE(_00104_),
    .Q(\w[50][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][13]$_SDFFCE_PN0P_  (.D(_02126_),
    .DE(_00104_),
    .Q(\w[50][13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][14]$_SDFFCE_PN0P_  (.D(_02127_),
    .DE(_00104_),
    .Q(\w[50][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][15]$_SDFFCE_PN0P_  (.D(_02128_),
    .DE(_00104_),
    .Q(\w[50][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][16]$_SDFFCE_PN0P_  (.D(_02129_),
    .DE(_00104_),
    .Q(\w[50][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][17]$_SDFFCE_PN0P_  (.D(_02130_),
    .DE(_00104_),
    .Q(\w[50][17] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][18]$_SDFFCE_PN0P_  (.D(_02131_),
    .DE(_00104_),
    .Q(\w[50][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][19]$_SDFFCE_PN0P_  (.D(_02132_),
    .DE(_00104_),
    .Q(\w[50][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][1]$_SDFFCE_PN0P_  (.D(_02133_),
    .DE(_00104_),
    .Q(\w[50][1] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][20]$_SDFFCE_PN0P_  (.D(_02134_),
    .DE(_00104_),
    .Q(\w[50][20] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][21]$_SDFFCE_PN0P_  (.D(_02135_),
    .DE(_00104_),
    .Q(\w[50][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][22]$_SDFFCE_PN0P_  (.D(_02136_),
    .DE(_00104_),
    .Q(\w[50][22] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][23]$_SDFFCE_PN0P_  (.D(_02137_),
    .DE(_00104_),
    .Q(\w[50][23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][24]$_SDFFCE_PN0P_  (.D(_02138_),
    .DE(_00104_),
    .Q(\w[50][24] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][25]$_SDFFCE_PN0P_  (.D(_02139_),
    .DE(_00104_),
    .Q(\w[50][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][26]$_SDFFCE_PN0P_  (.D(_02140_),
    .DE(_00104_),
    .Q(\w[50][26] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][27]$_SDFFCE_PN0P_  (.D(_02141_),
    .DE(_00104_),
    .Q(\w[50][27] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][28]$_SDFFCE_PN0P_  (.D(_02142_),
    .DE(_00104_),
    .Q(\w[50][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][29]$_SDFFCE_PN0P_  (.D(_02143_),
    .DE(_00104_),
    .Q(\w[50][29] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][2]$_SDFFCE_PN0P_  (.D(_02144_),
    .DE(_00104_),
    .Q(\w[50][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][30]$_SDFFCE_PN0P_  (.D(_02145_),
    .DE(_00104_),
    .Q(\w[50][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][31]$_SDFFCE_PN0P_  (.D(_02146_),
    .DE(_00104_),
    .Q(\w[50][31] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][3]$_SDFFCE_PN0P_  (.D(_02147_),
    .DE(_00104_),
    .Q(\w[50][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][4]$_SDFFCE_PN0P_  (.D(_02148_),
    .DE(_00104_),
    .Q(\w[50][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][5]$_SDFFCE_PN0P_  (.D(_02149_),
    .DE(_00104_),
    .Q(\w[50][5] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][6]$_SDFFCE_PN0P_  (.D(_02150_),
    .DE(_00104_),
    .Q(\w[50][6] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][7]$_SDFFCE_PN0P_  (.D(_02151_),
    .DE(_00104_),
    .Q(\w[50][7] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][8]$_SDFFCE_PN0P_  (.D(_02152_),
    .DE(_00104_),
    .Q(\w[50][8] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][9]$_SDFFCE_PN0P_  (.D(_02153_),
    .DE(_00104_),
    .Q(\w[50][9] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][0]$_SDFFCE_PN0P_  (.D(_02154_),
    .DE(_00073_),
    .Q(\w[51][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][10]$_SDFFCE_PN0P_  (.D(_02155_),
    .DE(_00073_),
    .Q(\w[51][10] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][11]$_SDFFCE_PN0P_  (.D(_02156_),
    .DE(_00073_),
    .Q(\w[51][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][12]$_SDFFCE_PN0P_  (.D(_02157_),
    .DE(_00073_),
    .Q(\w[51][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][13]$_SDFFCE_PN0P_  (.D(_02158_),
    .DE(_00073_),
    .Q(\w[51][13] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][14]$_SDFFCE_PN0P_  (.D(_02159_),
    .DE(_00073_),
    .Q(\w[51][14] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][15]$_SDFFCE_PN0P_  (.D(_02160_),
    .DE(_00073_),
    .Q(\w[51][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][16]$_SDFFCE_PN0P_  (.D(_02161_),
    .DE(_00073_),
    .Q(\w[51][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][17]$_SDFFCE_PN0P_  (.D(_02162_),
    .DE(_00073_),
    .Q(\w[51][17] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][18]$_SDFFCE_PN0P_  (.D(_02163_),
    .DE(_00073_),
    .Q(\w[51][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][19]$_SDFFCE_PN0P_  (.D(_02164_),
    .DE(_00073_),
    .Q(\w[51][19] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][1]$_SDFFCE_PN0P_  (.D(_02165_),
    .DE(_00073_),
    .Q(\w[51][1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][20]$_SDFFCE_PN0P_  (.D(_02166_),
    .DE(_00073_),
    .Q(\w[51][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][21]$_SDFFCE_PN0P_  (.D(_02167_),
    .DE(_00073_),
    .Q(\w[51][21] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][22]$_SDFFCE_PN0P_  (.D(_02168_),
    .DE(_00073_),
    .Q(\w[51][22] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][23]$_SDFFCE_PN0P_  (.D(_02169_),
    .DE(_00073_),
    .Q(\w[51][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][24]$_SDFFCE_PN0P_  (.D(_02170_),
    .DE(_00073_),
    .Q(\w[51][24] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][25]$_SDFFCE_PN0P_  (.D(_02171_),
    .DE(_00073_),
    .Q(\w[51][25] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][26]$_SDFFCE_PN0P_  (.D(_02172_),
    .DE(_00073_),
    .Q(\w[51][26] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][27]$_SDFFCE_PN0P_  (.D(_02173_),
    .DE(_00073_),
    .Q(\w[51][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][28]$_SDFFCE_PN0P_  (.D(_02174_),
    .DE(_00073_),
    .Q(\w[51][28] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][29]$_SDFFCE_PN0P_  (.D(_02175_),
    .DE(_00073_),
    .Q(\w[51][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][2]$_SDFFCE_PN0P_  (.D(_02176_),
    .DE(_00073_),
    .Q(\w[51][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][30]$_SDFFCE_PN0P_  (.D(_02177_),
    .DE(_00073_),
    .Q(\w[51][30] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][31]$_SDFFCE_PN0P_  (.D(_02178_),
    .DE(_00073_),
    .Q(\w[51][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][3]$_SDFFCE_PN0P_  (.D(_02179_),
    .DE(_00073_),
    .Q(\w[51][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][4]$_SDFFCE_PN0P_  (.D(_02180_),
    .DE(_00073_),
    .Q(\w[51][4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][5]$_SDFFCE_PN0P_  (.D(_02181_),
    .DE(_00073_),
    .Q(\w[51][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][6]$_SDFFCE_PN0P_  (.D(_02182_),
    .DE(_00073_),
    .Q(\w[51][6] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][7]$_SDFFCE_PN0P_  (.D(_02183_),
    .DE(_00073_),
    .Q(\w[51][7] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][8]$_SDFFCE_PN0P_  (.D(_02184_),
    .DE(_00073_),
    .Q(\w[51][8] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][9]$_SDFFCE_PN0P_  (.D(_02185_),
    .DE(_00073_),
    .Q(\w[51][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][0]$_SDFFCE_PN0P_  (.D(_02186_),
    .DE(_00103_),
    .Q(\w[52][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][10]$_SDFFCE_PN0P_  (.D(_02187_),
    .DE(_00103_),
    .Q(\w[52][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][11]$_SDFFCE_PN0P_  (.D(_02188_),
    .DE(_00103_),
    .Q(\w[52][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][12]$_SDFFCE_PN0P_  (.D(_02189_),
    .DE(_00103_),
    .Q(\w[52][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][13]$_SDFFCE_PN0P_  (.D(_02190_),
    .DE(_00103_),
    .Q(\w[52][13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][14]$_SDFFCE_PN0P_  (.D(_02191_),
    .DE(_00103_),
    .Q(\w[52][14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][15]$_SDFFCE_PN0P_  (.D(_02192_),
    .DE(_00103_),
    .Q(\w[52][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][16]$_SDFFCE_PN0P_  (.D(_02193_),
    .DE(_00103_),
    .Q(\w[52][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][17]$_SDFFCE_PN0P_  (.D(_02194_),
    .DE(_00103_),
    .Q(\w[52][17] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][18]$_SDFFCE_PN0P_  (.D(_02195_),
    .DE(_00103_),
    .Q(\w[52][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][19]$_SDFFCE_PN0P_  (.D(_02196_),
    .DE(_00103_),
    .Q(\w[52][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][1]$_SDFFCE_PN0P_  (.D(_02197_),
    .DE(_00103_),
    .Q(\w[52][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][20]$_SDFFCE_PN0P_  (.D(_02198_),
    .DE(_00103_),
    .Q(\w[52][20] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][21]$_SDFFCE_PN0P_  (.D(_02199_),
    .DE(_00103_),
    .Q(\w[52][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][22]$_SDFFCE_PN0P_  (.D(_02200_),
    .DE(_00103_),
    .Q(\w[52][22] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][23]$_SDFFCE_PN0P_  (.D(_02201_),
    .DE(_00103_),
    .Q(\w[52][23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][24]$_SDFFCE_PN0P_  (.D(_02202_),
    .DE(_00103_),
    .Q(\w[52][24] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][25]$_SDFFCE_PN0P_  (.D(_02203_),
    .DE(_00103_),
    .Q(\w[52][25] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][26]$_SDFFCE_PN0P_  (.D(_02204_),
    .DE(_00103_),
    .Q(\w[52][26] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][27]$_SDFFCE_PN0P_  (.D(_02205_),
    .DE(_00103_),
    .Q(\w[52][27] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][28]$_SDFFCE_PN0P_  (.D(_02206_),
    .DE(_00103_),
    .Q(\w[52][28] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][29]$_SDFFCE_PN0P_  (.D(_02207_),
    .DE(_00103_),
    .Q(\w[52][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][2]$_SDFFCE_PN0P_  (.D(_02208_),
    .DE(_00103_),
    .Q(\w[52][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][30]$_SDFFCE_PN0P_  (.D(_02209_),
    .DE(_00103_),
    .Q(\w[52][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][31]$_SDFFCE_PN0P_  (.D(_02210_),
    .DE(_00103_),
    .Q(\w[52][31] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][3]$_SDFFCE_PN0P_  (.D(_02211_),
    .DE(_00103_),
    .Q(\w[52][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][4]$_SDFFCE_PN0P_  (.D(_02212_),
    .DE(_00103_),
    .Q(\w[52][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][5]$_SDFFCE_PN0P_  (.D(_02213_),
    .DE(_00103_),
    .Q(\w[52][5] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][6]$_SDFFCE_PN0P_  (.D(_02214_),
    .DE(_00103_),
    .Q(\w[52][6] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][7]$_SDFFCE_PN0P_  (.D(_02215_),
    .DE(_00103_),
    .Q(\w[52][7] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][8]$_SDFFCE_PN0P_  (.D(_02216_),
    .DE(_00103_),
    .Q(\w[52][8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][9]$_SDFFCE_PN0P_  (.D(_02217_),
    .DE(_00103_),
    .Q(\w[52][9] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][0]$_SDFFCE_PN0P_  (.D(_02218_),
    .DE(_00072_),
    .Q(\w[53][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][10]$_SDFFCE_PN0P_  (.D(_02219_),
    .DE(_00072_),
    .Q(\w[53][10] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][11]$_SDFFCE_PN0P_  (.D(_02220_),
    .DE(_00072_),
    .Q(\w[53][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][12]$_SDFFCE_PN0P_  (.D(_02221_),
    .DE(_00072_),
    .Q(\w[53][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][13]$_SDFFCE_PN0P_  (.D(_02222_),
    .DE(_00072_),
    .Q(\w[53][13] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][14]$_SDFFCE_PN0P_  (.D(_02223_),
    .DE(_00072_),
    .Q(\w[53][14] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][15]$_SDFFCE_PN0P_  (.D(_02224_),
    .DE(_00072_),
    .Q(\w[53][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][16]$_SDFFCE_PN0P_  (.D(_02225_),
    .DE(_00072_),
    .Q(\w[53][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][17]$_SDFFCE_PN0P_  (.D(_02226_),
    .DE(_00072_),
    .Q(\w[53][17] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][18]$_SDFFCE_PN0P_  (.D(_02227_),
    .DE(_00072_),
    .Q(\w[53][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][19]$_SDFFCE_PN0P_  (.D(_02228_),
    .DE(_00072_),
    .Q(\w[53][19] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][1]$_SDFFCE_PN0P_  (.D(_02229_),
    .DE(_00072_),
    .Q(\w[53][1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][20]$_SDFFCE_PN0P_  (.D(_02230_),
    .DE(_00072_),
    .Q(\w[53][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][21]$_SDFFCE_PN0P_  (.D(_02231_),
    .DE(_00072_),
    .Q(\w[53][21] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][22]$_SDFFCE_PN0P_  (.D(_02232_),
    .DE(_00072_),
    .Q(\w[53][22] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][23]$_SDFFCE_PN0P_  (.D(_02233_),
    .DE(_00072_),
    .Q(\w[53][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][24]$_SDFFCE_PN0P_  (.D(_02234_),
    .DE(_00072_),
    .Q(\w[53][24] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][25]$_SDFFCE_PN0P_  (.D(_02235_),
    .DE(_00072_),
    .Q(\w[53][25] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][26]$_SDFFCE_PN0P_  (.D(_02236_),
    .DE(_00072_),
    .Q(\w[53][26] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][27]$_SDFFCE_PN0P_  (.D(_02237_),
    .DE(_00072_),
    .Q(\w[53][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][28]$_SDFFCE_PN0P_  (.D(_02238_),
    .DE(_00072_),
    .Q(\w[53][28] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][29]$_SDFFCE_PN0P_  (.D(_02239_),
    .DE(_00072_),
    .Q(\w[53][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][2]$_SDFFCE_PN0P_  (.D(_02240_),
    .DE(_00072_),
    .Q(\w[53][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][30]$_SDFFCE_PN0P_  (.D(_02241_),
    .DE(_00072_),
    .Q(\w[53][30] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][31]$_SDFFCE_PN0P_  (.D(_02242_),
    .DE(_00072_),
    .Q(\w[53][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][3]$_SDFFCE_PN0P_  (.D(_02243_),
    .DE(_00072_),
    .Q(\w[53][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][4]$_SDFFCE_PN0P_  (.D(_02244_),
    .DE(_00072_),
    .Q(\w[53][4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][5]$_SDFFCE_PN0P_  (.D(_02245_),
    .DE(_00072_),
    .Q(\w[53][5] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][6]$_SDFFCE_PN0P_  (.D(_02246_),
    .DE(_00072_),
    .Q(\w[53][6] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][7]$_SDFFCE_PN0P_  (.D(_02247_),
    .DE(_00072_),
    .Q(\w[53][7] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][8]$_SDFFCE_PN0P_  (.D(_02248_),
    .DE(_00072_),
    .Q(\w[53][8] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][9]$_SDFFCE_PN0P_  (.D(_02249_),
    .DE(_00072_),
    .Q(\w[53][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][0]$_SDFFCE_PN0P_  (.D(_02250_),
    .DE(_00102_),
    .Q(\w[54][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][10]$_SDFFCE_PN0P_  (.D(_02251_),
    .DE(_00102_),
    .Q(\w[54][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][11]$_SDFFCE_PN0P_  (.D(_02252_),
    .DE(_00102_),
    .Q(\w[54][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][12]$_SDFFCE_PN0P_  (.D(_02253_),
    .DE(_00102_),
    .Q(\w[54][12] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][13]$_SDFFCE_PN0P_  (.D(_02254_),
    .DE(_00102_),
    .Q(\w[54][13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][14]$_SDFFCE_PN0P_  (.D(_02255_),
    .DE(_00102_),
    .Q(\w[54][14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][15]$_SDFFCE_PN0P_  (.D(_02256_),
    .DE(_00102_),
    .Q(\w[54][15] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][16]$_SDFFCE_PN0P_  (.D(_02257_),
    .DE(_00102_),
    .Q(\w[54][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][17]$_SDFFCE_PN0P_  (.D(_02258_),
    .DE(_00102_),
    .Q(\w[54][17] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][18]$_SDFFCE_PN0P_  (.D(_02259_),
    .DE(_00102_),
    .Q(\w[54][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][19]$_SDFFCE_PN0P_  (.D(_02260_),
    .DE(_00102_),
    .Q(\w[54][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][1]$_SDFFCE_PN0P_  (.D(_02261_),
    .DE(_00102_),
    .Q(\w[54][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][20]$_SDFFCE_PN0P_  (.D(_02262_),
    .DE(_00102_),
    .Q(\w[54][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][21]$_SDFFCE_PN0P_  (.D(_02263_),
    .DE(_00102_),
    .Q(\w[54][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][22]$_SDFFCE_PN0P_  (.D(_02264_),
    .DE(_00102_),
    .Q(\w[54][22] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][23]$_SDFFCE_PN0P_  (.D(_02265_),
    .DE(_00102_),
    .Q(\w[54][23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][24]$_SDFFCE_PN0P_  (.D(_02266_),
    .DE(_00102_),
    .Q(\w[54][24] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][25]$_SDFFCE_PN0P_  (.D(_02267_),
    .DE(_00102_),
    .Q(\w[54][25] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][26]$_SDFFCE_PN0P_  (.D(_02268_),
    .DE(_00102_),
    .Q(\w[54][26] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][27]$_SDFFCE_PN0P_  (.D(_02269_),
    .DE(_00102_),
    .Q(\w[54][27] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][28]$_SDFFCE_PN0P_  (.D(_02270_),
    .DE(_00102_),
    .Q(\w[54][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][29]$_SDFFCE_PN0P_  (.D(_02271_),
    .DE(_00102_),
    .Q(\w[54][29] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][2]$_SDFFCE_PN0P_  (.D(_02272_),
    .DE(_00102_),
    .Q(\w[54][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][30]$_SDFFCE_PN0P_  (.D(_02273_),
    .DE(_00102_),
    .Q(\w[54][30] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][31]$_SDFFCE_PN0P_  (.D(_02274_),
    .DE(_00102_),
    .Q(\w[54][31] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][3]$_SDFFCE_PN0P_  (.D(_02275_),
    .DE(_00102_),
    .Q(\w[54][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][4]$_SDFFCE_PN0P_  (.D(_02276_),
    .DE(_00102_),
    .Q(\w[54][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][5]$_SDFFCE_PN0P_  (.D(_02277_),
    .DE(_00102_),
    .Q(\w[54][5] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][6]$_SDFFCE_PN0P_  (.D(_02278_),
    .DE(_00102_),
    .Q(\w[54][6] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][7]$_SDFFCE_PN0P_  (.D(_02279_),
    .DE(_00102_),
    .Q(\w[54][7] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][8]$_SDFFCE_PN0P_  (.D(_02280_),
    .DE(_00102_),
    .Q(\w[54][8] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][9]$_SDFFCE_PN0P_  (.D(_02281_),
    .DE(_00102_),
    .Q(\w[54][9] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][0]$_SDFFCE_PN0P_  (.D(_02282_),
    .DE(net471),
    .Q(\w[55][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][10]$_SDFFCE_PN0P_  (.D(_02283_),
    .DE(_00071_),
    .Q(\w[55][10] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][11]$_SDFFCE_PN0P_  (.D(_02284_),
    .DE(_00071_),
    .Q(\w[55][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][12]$_SDFFCE_PN0P_  (.D(_02285_),
    .DE(net471),
    .Q(\w[55][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][13]$_SDFFCE_PN0P_  (.D(_02286_),
    .DE(_00071_),
    .Q(\w[55][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][14]$_SDFFCE_PN0P_  (.D(_02287_),
    .DE(net471),
    .Q(\w[55][14] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][15]$_SDFFCE_PN0P_  (.D(_02288_),
    .DE(net471),
    .Q(\w[55][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][16]$_SDFFCE_PN0P_  (.D(_02289_),
    .DE(net471),
    .Q(\w[55][16] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][17]$_SDFFCE_PN0P_  (.D(_02290_),
    .DE(net470),
    .Q(\w[55][17] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][18]$_SDFFCE_PN0P_  (.D(_02291_),
    .DE(net470),
    .Q(\w[55][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][19]$_SDFFCE_PN0P_  (.D(_02292_),
    .DE(_00071_),
    .Q(\w[55][19] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][1]$_SDFFCE_PN0P_  (.D(_02293_),
    .DE(net471),
    .Q(\w[55][1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][20]$_SDFFCE_PN0P_  (.D(_02294_),
    .DE(_00071_),
    .Q(\w[55][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][21]$_SDFFCE_PN0P_  (.D(_02295_),
    .DE(_00071_),
    .Q(\w[55][21] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][22]$_SDFFCE_PN0P_  (.D(_02296_),
    .DE(_00071_),
    .Q(\w[55][22] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][23]$_SDFFCE_PN0P_  (.D(_02297_),
    .DE(net470),
    .Q(\w[55][23] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][24]$_SDFFCE_PN0P_  (.D(_02298_),
    .DE(net470),
    .Q(\w[55][24] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][25]$_SDFFCE_PN0P_  (.D(_02299_),
    .DE(net470),
    .Q(\w[55][25] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][26]$_SDFFCE_PN0P_  (.D(_02300_),
    .DE(net470),
    .Q(\w[55][26] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][27]$_SDFFCE_PN0P_  (.D(_02301_),
    .DE(net470),
    .Q(\w[55][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][28]$_SDFFCE_PN0P_  (.D(_02302_),
    .DE(net470),
    .Q(\w[55][28] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][29]$_SDFFCE_PN0P_  (.D(_02303_),
    .DE(_00071_),
    .Q(\w[55][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][2]$_SDFFCE_PN0P_  (.D(_02304_),
    .DE(net470),
    .Q(\w[55][2] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][30]$_SDFFCE_PN0P_  (.D(_02305_),
    .DE(net470),
    .Q(\w[55][30] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][31]$_SDFFCE_PN0P_  (.D(_02306_),
    .DE(net470),
    .Q(\w[55][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][3]$_SDFFCE_PN0P_  (.D(_02307_),
    .DE(net471),
    .Q(\w[55][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][4]$_SDFFCE_PN0P_  (.D(_02308_),
    .DE(net471),
    .Q(\w[55][4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][5]$_SDFFCE_PN0P_  (.D(_02309_),
    .DE(net471),
    .Q(\w[55][5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][6]$_SDFFCE_PN0P_  (.D(_02310_),
    .DE(net470),
    .Q(\w[55][6] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][7]$_SDFFCE_PN0P_  (.D(_02311_),
    .DE(net471),
    .Q(\w[55][7] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][8]$_SDFFCE_PN0P_  (.D(_02312_),
    .DE(net471),
    .Q(\w[55][8] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][9]$_SDFFCE_PN0P_  (.D(_02313_),
    .DE(_00071_),
    .Q(\w[55][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][0]$_SDFFCE_PN0P_  (.D(_02314_),
    .DE(_00101_),
    .Q(\w[56][0] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][10]$_SDFFCE_PN0P_  (.D(_02315_),
    .DE(_00101_),
    .Q(\w[56][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][11]$_SDFFCE_PN0P_  (.D(_02316_),
    .DE(_00101_),
    .Q(\w[56][11] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][12]$_SDFFCE_PN0P_  (.D(_02317_),
    .DE(_00101_),
    .Q(\w[56][12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][13]$_SDFFCE_PN0P_  (.D(_02318_),
    .DE(_00101_),
    .Q(\w[56][13] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][14]$_SDFFCE_PN0P_  (.D(_02319_),
    .DE(_00101_),
    .Q(\w[56][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][15]$_SDFFCE_PN0P_  (.D(_02320_),
    .DE(_00101_),
    .Q(\w[56][15] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][16]$_SDFFCE_PN0P_  (.D(_02321_),
    .DE(_00101_),
    .Q(\w[56][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][17]$_SDFFCE_PN0P_  (.D(_02322_),
    .DE(_00101_),
    .Q(\w[56][17] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][18]$_SDFFCE_PN0P_  (.D(_02323_),
    .DE(_00101_),
    .Q(\w[56][18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][19]$_SDFFCE_PN0P_  (.D(_02324_),
    .DE(_00101_),
    .Q(\w[56][19] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][1]$_SDFFCE_PN0P_  (.D(_02325_),
    .DE(_00101_),
    .Q(\w[56][1] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][20]$_SDFFCE_PN0P_  (.D(_02326_),
    .DE(_00101_),
    .Q(\w[56][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][21]$_SDFFCE_PN0P_  (.D(_02327_),
    .DE(_00101_),
    .Q(\w[56][21] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][22]$_SDFFCE_PN0P_  (.D(_02328_),
    .DE(_00101_),
    .Q(\w[56][22] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][23]$_SDFFCE_PN0P_  (.D(_02329_),
    .DE(_00101_),
    .Q(\w[56][23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][24]$_SDFFCE_PN0P_  (.D(_02330_),
    .DE(_00101_),
    .Q(\w[56][24] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][25]$_SDFFCE_PN0P_  (.D(_02331_),
    .DE(_00101_),
    .Q(\w[56][25] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][26]$_SDFFCE_PN0P_  (.D(_02332_),
    .DE(_00101_),
    .Q(\w[56][26] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][27]$_SDFFCE_PN0P_  (.D(_02333_),
    .DE(_00101_),
    .Q(\w[56][27] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][28]$_SDFFCE_PN0P_  (.D(_02334_),
    .DE(_00101_),
    .Q(\w[56][28] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][29]$_SDFFCE_PN0P_  (.D(_02335_),
    .DE(_00101_),
    .Q(\w[56][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][2]$_SDFFCE_PN0P_  (.D(_02336_),
    .DE(_00101_),
    .Q(\w[56][2] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][30]$_SDFFCE_PN0P_  (.D(_02337_),
    .DE(_00101_),
    .Q(\w[56][30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][31]$_SDFFCE_PN0P_  (.D(_02338_),
    .DE(_00101_),
    .Q(\w[56][31] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][3]$_SDFFCE_PN0P_  (.D(_02339_),
    .DE(_00101_),
    .Q(\w[56][3] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][4]$_SDFFCE_PN0P_  (.D(_02340_),
    .DE(_00101_),
    .Q(\w[56][4] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][5]$_SDFFCE_PN0P_  (.D(_02341_),
    .DE(_00101_),
    .Q(\w[56][5] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][6]$_SDFFCE_PN0P_  (.D(_02342_),
    .DE(_00101_),
    .Q(\w[56][6] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][7]$_SDFFCE_PN0P_  (.D(_02343_),
    .DE(_00101_),
    .Q(\w[56][7] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][8]$_SDFFCE_PN0P_  (.D(_02344_),
    .DE(_00101_),
    .Q(\w[56][8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][9]$_SDFFCE_PN0P_  (.D(_02345_),
    .DE(_00101_),
    .Q(\w[56][9] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][0]$_SDFFCE_PN0P_  (.D(_02346_),
    .DE(_00070_),
    .Q(\w[57][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][10]$_SDFFCE_PN0P_  (.D(_02347_),
    .DE(_00070_),
    .Q(\w[57][10] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][11]$_SDFFCE_PN0P_  (.D(_02348_),
    .DE(_00070_),
    .Q(\w[57][11] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][12]$_SDFFCE_PN0P_  (.D(_02349_),
    .DE(_00070_),
    .Q(\w[57][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][13]$_SDFFCE_PN0P_  (.D(_02350_),
    .DE(_00070_),
    .Q(\w[57][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][14]$_SDFFCE_PN0P_  (.D(_02351_),
    .DE(_00070_),
    .Q(\w[57][14] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][15]$_SDFFCE_PN0P_  (.D(_02352_),
    .DE(_00070_),
    .Q(\w[57][15] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][16]$_SDFFCE_PN0P_  (.D(_02353_),
    .DE(_00070_),
    .Q(\w[57][16] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][17]$_SDFFCE_PN0P_  (.D(_02354_),
    .DE(_00070_),
    .Q(\w[57][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][18]$_SDFFCE_PN0P_  (.D(_02355_),
    .DE(_00070_),
    .Q(\w[57][18] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][19]$_SDFFCE_PN0P_  (.D(_02356_),
    .DE(_00070_),
    .Q(\w[57][19] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][1]$_SDFFCE_PN0P_  (.D(_02357_),
    .DE(_00070_),
    .Q(\w[57][1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][20]$_SDFFCE_PN0P_  (.D(_02358_),
    .DE(_00070_),
    .Q(\w[57][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][21]$_SDFFCE_PN0P_  (.D(_02359_),
    .DE(_00070_),
    .Q(\w[57][21] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][22]$_SDFFCE_PN0P_  (.D(_02360_),
    .DE(_00070_),
    .Q(\w[57][22] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][23]$_SDFFCE_PN0P_  (.D(_02361_),
    .DE(_00070_),
    .Q(\w[57][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][24]$_SDFFCE_PN0P_  (.D(_02362_),
    .DE(_00070_),
    .Q(\w[57][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][25]$_SDFFCE_PN0P_  (.D(_02363_),
    .DE(_00070_),
    .Q(\w[57][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][26]$_SDFFCE_PN0P_  (.D(_02364_),
    .DE(_00070_),
    .Q(\w[57][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][27]$_SDFFCE_PN0P_  (.D(_02365_),
    .DE(_00070_),
    .Q(\w[57][27] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][28]$_SDFFCE_PN0P_  (.D(_02366_),
    .DE(_00070_),
    .Q(\w[57][28] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][29]$_SDFFCE_PN0P_  (.D(_02367_),
    .DE(_00070_),
    .Q(\w[57][29] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][2]$_SDFFCE_PN0P_  (.D(_02368_),
    .DE(_00070_),
    .Q(\w[57][2] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][30]$_SDFFCE_PN0P_  (.D(_02369_),
    .DE(_00070_),
    .Q(\w[57][30] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][31]$_SDFFCE_PN0P_  (.D(_02370_),
    .DE(_00070_),
    .Q(\w[57][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][3]$_SDFFCE_PN0P_  (.D(_02371_),
    .DE(_00070_),
    .Q(\w[57][3] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][4]$_SDFFCE_PN0P_  (.D(_02372_),
    .DE(_00070_),
    .Q(\w[57][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][5]$_SDFFCE_PN0P_  (.D(_02373_),
    .DE(_00070_),
    .Q(\w[57][5] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][6]$_SDFFCE_PN0P_  (.D(_02374_),
    .DE(_00070_),
    .Q(\w[57][6] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][7]$_SDFFCE_PN0P_  (.D(_02375_),
    .DE(_00070_),
    .Q(\w[57][7] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][8]$_SDFFCE_PN0P_  (.D(_02376_),
    .DE(_00070_),
    .Q(\w[57][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][9]$_SDFFCE_PN0P_  (.D(_02377_),
    .DE(_00070_),
    .Q(\w[57][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][0]$_SDFFCE_PN0P_  (.D(_02378_),
    .DE(_00100_),
    .Q(\w[58][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][10]$_SDFFCE_PN0P_  (.D(_02379_),
    .DE(_00100_),
    .Q(\w[58][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][11]$_SDFFCE_PN0P_  (.D(_02380_),
    .DE(_00100_),
    .Q(\w[58][11] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][12]$_SDFFCE_PN0P_  (.D(_02381_),
    .DE(_00100_),
    .Q(\w[58][12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][13]$_SDFFCE_PN0P_  (.D(_02382_),
    .DE(_00100_),
    .Q(\w[58][13] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][14]$_SDFFCE_PN0P_  (.D(_02383_),
    .DE(_00100_),
    .Q(\w[58][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][15]$_SDFFCE_PN0P_  (.D(_02384_),
    .DE(_00100_),
    .Q(\w[58][15] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][16]$_SDFFCE_PN0P_  (.D(_02385_),
    .DE(_00100_),
    .Q(\w[58][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][17]$_SDFFCE_PN0P_  (.D(_02386_),
    .DE(_00100_),
    .Q(\w[58][17] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][18]$_SDFFCE_PN0P_  (.D(_02387_),
    .DE(_00100_),
    .Q(\w[58][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][19]$_SDFFCE_PN0P_  (.D(_02388_),
    .DE(_00100_),
    .Q(\w[58][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][1]$_SDFFCE_PN0P_  (.D(_02389_),
    .DE(_00100_),
    .Q(\w[58][1] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][20]$_SDFFCE_PN0P_  (.D(_02390_),
    .DE(_00100_),
    .Q(\w[58][20] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][21]$_SDFFCE_PN0P_  (.D(_02391_),
    .DE(_00100_),
    .Q(\w[58][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][22]$_SDFFCE_PN0P_  (.D(_02392_),
    .DE(_00100_),
    .Q(\w[58][22] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][23]$_SDFFCE_PN0P_  (.D(_02393_),
    .DE(_00100_),
    .Q(\w[58][23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][24]$_SDFFCE_PN0P_  (.D(_02394_),
    .DE(_00100_),
    .Q(\w[58][24] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][25]$_SDFFCE_PN0P_  (.D(_02395_),
    .DE(_00100_),
    .Q(\w[58][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][26]$_SDFFCE_PN0P_  (.D(_02396_),
    .DE(_00100_),
    .Q(\w[58][26] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][27]$_SDFFCE_PN0P_  (.D(_02397_),
    .DE(_00100_),
    .Q(\w[58][27] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][28]$_SDFFCE_PN0P_  (.D(_02398_),
    .DE(_00100_),
    .Q(\w[58][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][29]$_SDFFCE_PN0P_  (.D(_02399_),
    .DE(_00100_),
    .Q(\w[58][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][2]$_SDFFCE_PN0P_  (.D(_02400_),
    .DE(_00100_),
    .Q(\w[58][2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][30]$_SDFFCE_PN0P_  (.D(_02401_),
    .DE(_00100_),
    .Q(\w[58][30] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][31]$_SDFFCE_PN0P_  (.D(_02402_),
    .DE(_00100_),
    .Q(\w[58][31] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][3]$_SDFFCE_PN0P_  (.D(_02403_),
    .DE(_00100_),
    .Q(\w[58][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][4]$_SDFFCE_PN0P_  (.D(_02404_),
    .DE(_00100_),
    .Q(\w[58][4] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][5]$_SDFFCE_PN0P_  (.D(_02405_),
    .DE(_00100_),
    .Q(\w[58][5] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][6]$_SDFFCE_PN0P_  (.D(_02406_),
    .DE(_00100_),
    .Q(\w[58][6] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][7]$_SDFFCE_PN0P_  (.D(_02407_),
    .DE(_00100_),
    .Q(\w[58][7] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][8]$_SDFFCE_PN0P_  (.D(_02408_),
    .DE(_00100_),
    .Q(\w[58][8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][9]$_SDFFCE_PN0P_  (.D(_02409_),
    .DE(_00100_),
    .Q(\w[58][9] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][0]$_SDFFCE_PN0P_  (.D(_02410_),
    .DE(_00069_),
    .Q(\w[59][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][10]$_SDFFCE_PN0P_  (.D(_02411_),
    .DE(_00069_),
    .Q(\w[59][10] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][11]$_SDFFCE_PN0P_  (.D(_02412_),
    .DE(_00069_),
    .Q(\w[59][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][12]$_SDFFCE_PN0P_  (.D(_02413_),
    .DE(_00069_),
    .Q(\w[59][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][13]$_SDFFCE_PN0P_  (.D(_02414_),
    .DE(_00069_),
    .Q(\w[59][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][14]$_SDFFCE_PN0P_  (.D(_02415_),
    .DE(_00069_),
    .Q(\w[59][14] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][15]$_SDFFCE_PN0P_  (.D(_02416_),
    .DE(_00069_),
    .Q(\w[59][15] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][16]$_SDFFCE_PN0P_  (.D(_02417_),
    .DE(_00069_),
    .Q(\w[59][16] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][17]$_SDFFCE_PN0P_  (.D(_02418_),
    .DE(_00069_),
    .Q(\w[59][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][18]$_SDFFCE_PN0P_  (.D(_02419_),
    .DE(_00069_),
    .Q(\w[59][18] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][19]$_SDFFCE_PN0P_  (.D(_02420_),
    .DE(_00069_),
    .Q(\w[59][19] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][1]$_SDFFCE_PN0P_  (.D(_02421_),
    .DE(_00069_),
    .Q(\w[59][1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][20]$_SDFFCE_PN0P_  (.D(_02422_),
    .DE(_00069_),
    .Q(\w[59][20] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][21]$_SDFFCE_PN0P_  (.D(_02423_),
    .DE(_00069_),
    .Q(\w[59][21] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][22]$_SDFFCE_PN0P_  (.D(_02424_),
    .DE(_00069_),
    .Q(\w[59][22] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][23]$_SDFFCE_PN0P_  (.D(_02425_),
    .DE(_00069_),
    .Q(\w[59][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][24]$_SDFFCE_PN0P_  (.D(_02426_),
    .DE(_00069_),
    .Q(\w[59][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][25]$_SDFFCE_PN0P_  (.D(_02427_),
    .DE(_00069_),
    .Q(\w[59][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][26]$_SDFFCE_PN0P_  (.D(_02428_),
    .DE(_00069_),
    .Q(\w[59][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][27]$_SDFFCE_PN0P_  (.D(_02429_),
    .DE(_00069_),
    .Q(\w[59][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][28]$_SDFFCE_PN0P_  (.D(_02430_),
    .DE(_00069_),
    .Q(\w[59][28] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][29]$_SDFFCE_PN0P_  (.D(_02431_),
    .DE(_00069_),
    .Q(\w[59][29] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][2]$_SDFFCE_PN0P_  (.D(_02432_),
    .DE(_00069_),
    .Q(\w[59][2] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][30]$_SDFFCE_PN0P_  (.D(_02433_),
    .DE(_00069_),
    .Q(\w[59][30] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][31]$_SDFFCE_PN0P_  (.D(_02434_),
    .DE(_00069_),
    .Q(\w[59][31] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][3]$_SDFFCE_PN0P_  (.D(_02435_),
    .DE(_00069_),
    .Q(\w[59][3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][4]$_SDFFCE_PN0P_  (.D(_02436_),
    .DE(_00069_),
    .Q(\w[59][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][5]$_SDFFCE_PN0P_  (.D(_02437_),
    .DE(_00069_),
    .Q(\w[59][5] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][6]$_SDFFCE_PN0P_  (.D(_02438_),
    .DE(_00069_),
    .Q(\w[59][6] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][7]$_SDFFCE_PN0P_  (.D(_02439_),
    .DE(_00069_),
    .Q(\w[59][7] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][8]$_SDFFCE_PN0P_  (.D(_02440_),
    .DE(_00069_),
    .Q(\w[59][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][9]$_SDFFCE_PN0P_  (.D(_02441_),
    .DE(_00069_),
    .Q(\w[59][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][0]$_DFFE_PP_  (.D(_00481_),
    .DE(_00068_),
    .Q(\w[5][0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][10]$_DFFE_PP_  (.D(_00482_),
    .DE(_00068_),
    .Q(\w[5][10] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][11]$_DFFE_PP_  (.D(_00483_),
    .DE(_00068_),
    .Q(\w[5][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][12]$_DFFE_PP_  (.D(_00484_),
    .DE(_00068_),
    .Q(\w[5][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][13]$_DFFE_PP_  (.D(_00485_),
    .DE(_00068_),
    .Q(\w[5][13] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][14]$_DFFE_PP_  (.D(_00486_),
    .DE(_00068_),
    .Q(\w[5][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][15]$_DFFE_PP_  (.D(_00487_),
    .DE(_00068_),
    .Q(\w[5][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][16]$_DFFE_PP_  (.D(_00488_),
    .DE(_00068_),
    .Q(\w[5][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][17]$_DFFE_PP_  (.D(_00489_),
    .DE(_00068_),
    .Q(\w[5][17] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][18]$_DFFE_PP_  (.D(_00490_),
    .DE(_00068_),
    .Q(\w[5][18] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][19]$_DFFE_PP_  (.D(_00491_),
    .DE(_00068_),
    .Q(\w[5][19] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][1]$_DFFE_PP_  (.D(_00492_),
    .DE(_00068_),
    .Q(\w[5][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][20]$_DFFE_PP_  (.D(_00493_),
    .DE(_00068_),
    .Q(\w[5][20] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][21]$_DFFE_PP_  (.D(_00494_),
    .DE(_00068_),
    .Q(\w[5][21] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][22]$_DFFE_PP_  (.D(_00495_),
    .DE(_00068_),
    .Q(\w[5][22] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][23]$_DFFE_PP_  (.D(_00496_),
    .DE(_00068_),
    .Q(\w[5][23] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][24]$_DFFE_PP_  (.D(_00497_),
    .DE(_00068_),
    .Q(\w[5][24] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][25]$_DFFE_PP_  (.D(_00498_),
    .DE(_00068_),
    .Q(\w[5][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][26]$_DFFE_PP_  (.D(_00499_),
    .DE(_00068_),
    .Q(\w[5][26] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][27]$_DFFE_PP_  (.D(_00500_),
    .DE(_00068_),
    .Q(\w[5][27] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][28]$_DFFE_PP_  (.D(_00501_),
    .DE(_00068_),
    .Q(\w[5][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][29]$_DFFE_PP_  (.D(_00502_),
    .DE(_00068_),
    .Q(\w[5][29] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][2]$_DFFE_PP_  (.D(_00503_),
    .DE(_00068_),
    .Q(\w[5][2] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][30]$_DFFE_PP_  (.D(_00504_),
    .DE(_00068_),
    .Q(\w[5][30] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][31]$_DFFE_PP_  (.D(_00505_),
    .DE(_00068_),
    .Q(\w[5][31] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][3]$_DFFE_PP_  (.D(_00506_),
    .DE(_00068_),
    .Q(\w[5][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][4]$_DFFE_PP_  (.D(_00507_),
    .DE(_00068_),
    .Q(\w[5][4] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][5]$_DFFE_PP_  (.D(_00508_),
    .DE(_00068_),
    .Q(\w[5][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][6]$_DFFE_PP_  (.D(_00509_),
    .DE(_00068_),
    .Q(\w[5][6] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][7]$_DFFE_PP_  (.D(_00510_),
    .DE(_00068_),
    .Q(\w[5][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][8]$_DFFE_PP_  (.D(_00511_),
    .DE(_00068_),
    .Q(\w[5][8] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][9]$_DFFE_PP_  (.D(_00512_),
    .DE(_00068_),
    .Q(\w[5][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][0]$_SDFFCE_PN0P_  (.D(_02442_),
    .DE(_00099_),
    .Q(\w[60][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][10]$_SDFFCE_PN0P_  (.D(_02443_),
    .DE(_00099_),
    .Q(\w[60][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][11]$_SDFFCE_PN0P_  (.D(_02444_),
    .DE(_00099_),
    .Q(\w[60][11] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][12]$_SDFFCE_PN0P_  (.D(_02445_),
    .DE(_00099_),
    .Q(\w[60][12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][13]$_SDFFCE_PN0P_  (.D(_02446_),
    .DE(_00099_),
    .Q(\w[60][13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][14]$_SDFFCE_PN0P_  (.D(_02447_),
    .DE(_00099_),
    .Q(\w[60][14] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][15]$_SDFFCE_PN0P_  (.D(_02448_),
    .DE(_00099_),
    .Q(\w[60][15] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][16]$_SDFFCE_PN0P_  (.D(_02449_),
    .DE(_00099_),
    .Q(\w[60][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][17]$_SDFFCE_PN0P_  (.D(_02450_),
    .DE(_00099_),
    .Q(\w[60][17] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][18]$_SDFFCE_PN0P_  (.D(_02451_),
    .DE(_00099_),
    .Q(\w[60][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][19]$_SDFFCE_PN0P_  (.D(_02452_),
    .DE(_00099_),
    .Q(\w[60][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][1]$_SDFFCE_PN0P_  (.D(_02453_),
    .DE(_00099_),
    .Q(\w[60][1] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][20]$_SDFFCE_PN0P_  (.D(_02454_),
    .DE(_00099_),
    .Q(\w[60][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][21]$_SDFFCE_PN0P_  (.D(_02455_),
    .DE(_00099_),
    .Q(\w[60][21] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][22]$_SDFFCE_PN0P_  (.D(_02456_),
    .DE(_00099_),
    .Q(\w[60][22] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][23]$_SDFFCE_PN0P_  (.D(_02457_),
    .DE(_00099_),
    .Q(\w[60][23] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][24]$_SDFFCE_PN0P_  (.D(_02458_),
    .DE(_00099_),
    .Q(\w[60][24] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][25]$_SDFFCE_PN0P_  (.D(_02459_),
    .DE(_00099_),
    .Q(\w[60][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][26]$_SDFFCE_PN0P_  (.D(_02460_),
    .DE(_00099_),
    .Q(\w[60][26] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][27]$_SDFFCE_PN0P_  (.D(_02461_),
    .DE(_00099_),
    .Q(\w[60][27] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][28]$_SDFFCE_PN0P_  (.D(_02462_),
    .DE(_00099_),
    .Q(\w[60][28] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][29]$_SDFFCE_PN0P_  (.D(_02463_),
    .DE(_00099_),
    .Q(\w[60][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][2]$_SDFFCE_PN0P_  (.D(_02464_),
    .DE(_00099_),
    .Q(\w[60][2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][30]$_SDFFCE_PN0P_  (.D(_02465_),
    .DE(_00099_),
    .Q(\w[60][30] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][31]$_SDFFCE_PN0P_  (.D(_02466_),
    .DE(_00099_),
    .Q(\w[60][31] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][3]$_SDFFCE_PN0P_  (.D(_02467_),
    .DE(_00099_),
    .Q(\w[60][3] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][4]$_SDFFCE_PN0P_  (.D(_02468_),
    .DE(_00099_),
    .Q(\w[60][4] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][5]$_SDFFCE_PN0P_  (.D(_02469_),
    .DE(_00099_),
    .Q(\w[60][5] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][6]$_SDFFCE_PN0P_  (.D(_02470_),
    .DE(_00099_),
    .Q(\w[60][6] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][7]$_SDFFCE_PN0P_  (.D(_02471_),
    .DE(_00099_),
    .Q(\w[60][7] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][8]$_SDFFCE_PN0P_  (.D(_02472_),
    .DE(_00099_),
    .Q(\w[60][8] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][9]$_SDFFCE_PN0P_  (.D(_02473_),
    .DE(_00099_),
    .Q(\w[60][9] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][0]$_SDFFCE_PN0P_  (.D(_02474_),
    .DE(_00067_),
    .Q(\w[61][0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][10]$_SDFFCE_PN0P_  (.D(_02475_),
    .DE(_00067_),
    .Q(\w[61][10] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][11]$_SDFFCE_PN0P_  (.D(_02476_),
    .DE(_00067_),
    .Q(\w[61][11] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][12]$_SDFFCE_PN0P_  (.D(_02477_),
    .DE(_00067_),
    .Q(\w[61][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][13]$_SDFFCE_PN0P_  (.D(_02478_),
    .DE(_00067_),
    .Q(\w[61][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][14]$_SDFFCE_PN0P_  (.D(_02479_),
    .DE(_00067_),
    .Q(\w[61][14] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][15]$_SDFFCE_PN0P_  (.D(_02480_),
    .DE(_00067_),
    .Q(\w[61][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][16]$_SDFFCE_PN0P_  (.D(_02481_),
    .DE(_00067_),
    .Q(\w[61][16] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][17]$_SDFFCE_PN0P_  (.D(_02482_),
    .DE(_00067_),
    .Q(\w[61][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][18]$_SDFFCE_PN0P_  (.D(_02483_),
    .DE(_00067_),
    .Q(\w[61][18] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][19]$_SDFFCE_PN0P_  (.D(_02484_),
    .DE(_00067_),
    .Q(\w[61][19] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][1]$_SDFFCE_PN0P_  (.D(_02485_),
    .DE(_00067_),
    .Q(\w[61][1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][20]$_SDFFCE_PN0P_  (.D(_02486_),
    .DE(_00067_),
    .Q(\w[61][20] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][21]$_SDFFCE_PN0P_  (.D(_02487_),
    .DE(_00067_),
    .Q(\w[61][21] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][22]$_SDFFCE_PN0P_  (.D(_02488_),
    .DE(_00067_),
    .Q(\w[61][22] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][23]$_SDFFCE_PN0P_  (.D(_02489_),
    .DE(_00067_),
    .Q(\w[61][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][24]$_SDFFCE_PN0P_  (.D(_02490_),
    .DE(_00067_),
    .Q(\w[61][24] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][25]$_SDFFCE_PN0P_  (.D(_02491_),
    .DE(_00067_),
    .Q(\w[61][25] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][26]$_SDFFCE_PN0P_  (.D(_02492_),
    .DE(_00067_),
    .Q(\w[61][26] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][27]$_SDFFCE_PN0P_  (.D(_02493_),
    .DE(_00067_),
    .Q(\w[61][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][28]$_SDFFCE_PN0P_  (.D(_02494_),
    .DE(_00067_),
    .Q(\w[61][28] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][29]$_SDFFCE_PN0P_  (.D(_02495_),
    .DE(_00067_),
    .Q(\w[61][29] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][2]$_SDFFCE_PN0P_  (.D(_02496_),
    .DE(_00067_),
    .Q(\w[61][2] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][30]$_SDFFCE_PN0P_  (.D(_02497_),
    .DE(_00067_),
    .Q(\w[61][30] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][31]$_SDFFCE_PN0P_  (.D(_02498_),
    .DE(_00067_),
    .Q(\w[61][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][3]$_SDFFCE_PN0P_  (.D(_02499_),
    .DE(_00067_),
    .Q(\w[61][3] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][4]$_SDFFCE_PN0P_  (.D(_02500_),
    .DE(_00067_),
    .Q(\w[61][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][5]$_SDFFCE_PN0P_  (.D(_02501_),
    .DE(_00067_),
    .Q(\w[61][5] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][6]$_SDFFCE_PN0P_  (.D(_02502_),
    .DE(_00067_),
    .Q(\w[61][6] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][7]$_SDFFCE_PN0P_  (.D(_02503_),
    .DE(_00067_),
    .Q(\w[61][7] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][8]$_SDFFCE_PN0P_  (.D(_02504_),
    .DE(_00067_),
    .Q(\w[61][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][9]$_SDFFCE_PN0P_  (.D(_02505_),
    .DE(_00067_),
    .Q(\w[61][9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][0]$_SDFFCE_PN0P_  (.D(_02506_),
    .DE(_00098_),
    .Q(\w[62][0] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][10]$_SDFFCE_PN0P_  (.D(_02507_),
    .DE(_00098_),
    .Q(\w[62][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][11]$_SDFFCE_PN0P_  (.D(_02508_),
    .DE(_00098_),
    .Q(\w[62][11] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][12]$_SDFFCE_PN0P_  (.D(_02509_),
    .DE(_00098_),
    .Q(\w[62][12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][13]$_SDFFCE_PN0P_  (.D(_02510_),
    .DE(_00098_),
    .Q(\w[62][13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][14]$_SDFFCE_PN0P_  (.D(_02511_),
    .DE(_00098_),
    .Q(\w[62][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][15]$_SDFFCE_PN0P_  (.D(_02512_),
    .DE(_00098_),
    .Q(\w[62][15] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][16]$_SDFFCE_PN0P_  (.D(_02513_),
    .DE(_00098_),
    .Q(\w[62][16] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][17]$_SDFFCE_PN0P_  (.D(_02514_),
    .DE(_00098_),
    .Q(\w[62][17] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][18]$_SDFFCE_PN0P_  (.D(_02515_),
    .DE(_00098_),
    .Q(\w[62][18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][19]$_SDFFCE_PN0P_  (.D(_02516_),
    .DE(_00098_),
    .Q(\w[62][19] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][1]$_SDFFCE_PN0P_  (.D(_02517_),
    .DE(_00098_),
    .Q(\w[62][1] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][20]$_SDFFCE_PN0P_  (.D(_02518_),
    .DE(_00098_),
    .Q(\w[62][20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][21]$_SDFFCE_PN0P_  (.D(_02519_),
    .DE(_00098_),
    .Q(\w[62][21] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][22]$_SDFFCE_PN0P_  (.D(_02520_),
    .DE(_00098_),
    .Q(\w[62][22] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][23]$_SDFFCE_PN0P_  (.D(_02521_),
    .DE(_00098_),
    .Q(\w[62][23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][24]$_SDFFCE_PN0P_  (.D(_02522_),
    .DE(_00098_),
    .Q(\w[62][24] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][25]$_SDFFCE_PN0P_  (.D(_02523_),
    .DE(_00098_),
    .Q(\w[62][25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][26]$_SDFFCE_PN0P_  (.D(_02524_),
    .DE(_00098_),
    .Q(\w[62][26] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][27]$_SDFFCE_PN0P_  (.D(_02525_),
    .DE(_00098_),
    .Q(\w[62][27] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][28]$_SDFFCE_PN0P_  (.D(_02526_),
    .DE(_00098_),
    .Q(\w[62][28] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][29]$_SDFFCE_PN0P_  (.D(_02527_),
    .DE(_00098_),
    .Q(\w[62][29] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][2]$_SDFFCE_PN0P_  (.D(_02528_),
    .DE(_00098_),
    .Q(\w[62][2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][30]$_SDFFCE_PN0P_  (.D(_02529_),
    .DE(_00098_),
    .Q(\w[62][30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][31]$_SDFFCE_PN0P_  (.D(_02530_),
    .DE(_00098_),
    .Q(\w[62][31] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][3]$_SDFFCE_PN0P_  (.D(_02531_),
    .DE(_00098_),
    .Q(\w[62][3] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][4]$_SDFFCE_PN0P_  (.D(_02532_),
    .DE(_00098_),
    .Q(\w[62][4] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][5]$_SDFFCE_PN0P_  (.D(_02533_),
    .DE(_00098_),
    .Q(\w[62][5] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][6]$_SDFFCE_PN0P_  (.D(_02534_),
    .DE(_00098_),
    .Q(\w[62][6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][7]$_SDFFCE_PN0P_  (.D(_02535_),
    .DE(_00098_),
    .Q(\w[62][7] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][8]$_SDFFCE_PN0P_  (.D(_02536_),
    .DE(_00098_),
    .Q(\w[62][8] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][9]$_SDFFCE_PN0P_  (.D(_02537_),
    .DE(_00098_),
    .Q(\w[62][9] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][0]$_SDFFCE_PN0P_  (.D(_02538_),
    .DE(_00066_),
    .Q(\w[63][0] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][10]$_SDFFCE_PN0P_  (.D(_02539_),
    .DE(_00066_),
    .Q(\w[63][10] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][11]$_SDFFCE_PN0P_  (.D(_02540_),
    .DE(_00066_),
    .Q(\w[63][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][12]$_SDFFCE_PN0P_  (.D(_02541_),
    .DE(_00066_),
    .Q(\w[63][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][13]$_SDFFCE_PN0P_  (.D(_02542_),
    .DE(_00066_),
    .Q(\w[63][13] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][14]$_SDFFCE_PN0P_  (.D(_02543_),
    .DE(_00066_),
    .Q(\w[63][14] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][15]$_SDFFCE_PN0P_  (.D(_02544_),
    .DE(_00066_),
    .Q(\w[63][15] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][16]$_SDFFCE_PN0P_  (.D(_02545_),
    .DE(_00066_),
    .Q(\w[63][16] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][17]$_SDFFCE_PN0P_  (.D(_02546_),
    .DE(_00066_),
    .Q(\w[63][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][18]$_SDFFCE_PN0P_  (.D(_02547_),
    .DE(_00066_),
    .Q(\w[63][18] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][19]$_SDFFCE_PN0P_  (.D(_02548_),
    .DE(_00066_),
    .Q(\w[63][19] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][1]$_SDFFCE_PN0P_  (.D(_02549_),
    .DE(_00066_),
    .Q(\w[63][1] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][20]$_SDFFCE_PN0P_  (.D(_02550_),
    .DE(_00066_),
    .Q(\w[63][20] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][21]$_SDFFCE_PN0P_  (.D(_02551_),
    .DE(_00066_),
    .Q(\w[63][21] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][22]$_SDFFCE_PN0P_  (.D(_02552_),
    .DE(_00066_),
    .Q(\w[63][22] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][23]$_SDFFCE_PN0P_  (.D(_02553_),
    .DE(_00066_),
    .Q(\w[63][23] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][24]$_SDFFCE_PN0P_  (.D(_02554_),
    .DE(_00066_),
    .Q(\w[63][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][25]$_SDFFCE_PN0P_  (.D(_02555_),
    .DE(_00066_),
    .Q(\w[63][25] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][26]$_SDFFCE_PN0P_  (.D(_02556_),
    .DE(_00066_),
    .Q(\w[63][26] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][27]$_SDFFCE_PN0P_  (.D(_02557_),
    .DE(_00066_),
    .Q(\w[63][27] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][28]$_SDFFCE_PN0P_  (.D(_02558_),
    .DE(_00066_),
    .Q(\w[63][28] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][29]$_SDFFCE_PN0P_  (.D(_02559_),
    .DE(_00066_),
    .Q(\w[63][29] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][2]$_SDFFCE_PN0P_  (.D(_02560_),
    .DE(_00066_),
    .Q(\w[63][2] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][30]$_SDFFCE_PN0P_  (.D(_02561_),
    .DE(_00066_),
    .Q(\w[63][30] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][31]$_SDFFCE_PN0P_  (.D(_02562_),
    .DE(_00066_),
    .Q(\w[63][31] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][3]$_SDFFCE_PN0P_  (.D(_02563_),
    .DE(_00066_),
    .Q(\w[63][3] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][4]$_SDFFCE_PN0P_  (.D(_02564_),
    .DE(_00066_),
    .Q(\w[63][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][5]$_SDFFCE_PN0P_  (.D(_02565_),
    .DE(_00066_),
    .Q(\w[63][5] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][6]$_SDFFCE_PN0P_  (.D(_02566_),
    .DE(_00066_),
    .Q(\w[63][6] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][7]$_SDFFCE_PN0P_  (.D(_02567_),
    .DE(_00066_),
    .Q(\w[63][7] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][8]$_SDFFCE_PN0P_  (.D(_02568_),
    .DE(_00066_),
    .Q(\w[63][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][9]$_SDFFCE_PN0P_  (.D(_02569_),
    .DE(_00066_),
    .Q(\w[63][9] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][0]$_DFFE_PP_  (.D(_00513_),
    .DE(_00097_),
    .Q(\w[6][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][10]$_DFFE_PP_  (.D(_00514_),
    .DE(_00097_),
    .Q(\w[6][10] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][11]$_DFFE_PP_  (.D(_00515_),
    .DE(_00097_),
    .Q(\w[6][11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][12]$_DFFE_PP_  (.D(_00516_),
    .DE(_00097_),
    .Q(\w[6][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][13]$_DFFE_PP_  (.D(_00517_),
    .DE(_00097_),
    .Q(\w[6][13] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][14]$_DFFE_PP_  (.D(_00518_),
    .DE(_00097_),
    .Q(\w[6][14] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][15]$_DFFE_PP_  (.D(_00519_),
    .DE(_00097_),
    .Q(\w[6][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][16]$_DFFE_PP_  (.D(_00520_),
    .DE(_00097_),
    .Q(\w[6][16] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][17]$_DFFE_PP_  (.D(_00521_),
    .DE(_00097_),
    .Q(\w[6][17] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][18]$_DFFE_PP_  (.D(_00522_),
    .DE(_00097_),
    .Q(\w[6][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][19]$_DFFE_PP_  (.D(_00523_),
    .DE(_00097_),
    .Q(\w[6][19] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][1]$_DFFE_PP_  (.D(_00524_),
    .DE(_00097_),
    .Q(\w[6][1] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][20]$_DFFE_PP_  (.D(_00525_),
    .DE(_00097_),
    .Q(\w[6][20] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][21]$_DFFE_PP_  (.D(_00526_),
    .DE(_00097_),
    .Q(\w[6][21] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][22]$_DFFE_PP_  (.D(_00527_),
    .DE(_00097_),
    .Q(\w[6][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][23]$_DFFE_PP_  (.D(_00528_),
    .DE(_00097_),
    .Q(\w[6][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][24]$_DFFE_PP_  (.D(_00529_),
    .DE(_00097_),
    .Q(\w[6][24] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][25]$_DFFE_PP_  (.D(_00530_),
    .DE(_00097_),
    .Q(\w[6][25] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][26]$_DFFE_PP_  (.D(_00531_),
    .DE(_00097_),
    .Q(\w[6][26] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][27]$_DFFE_PP_  (.D(_00532_),
    .DE(_00097_),
    .Q(\w[6][27] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][28]$_DFFE_PP_  (.D(_00533_),
    .DE(_00097_),
    .Q(\w[6][28] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][29]$_DFFE_PP_  (.D(_00534_),
    .DE(_00097_),
    .Q(\w[6][29] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][2]$_DFFE_PP_  (.D(_00535_),
    .DE(_00097_),
    .Q(\w[6][2] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][30]$_DFFE_PP_  (.D(_00536_),
    .DE(_00097_),
    .Q(\w[6][30] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][31]$_DFFE_PP_  (.D(_00537_),
    .DE(_00097_),
    .Q(\w[6][31] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][3]$_DFFE_PP_  (.D(_00538_),
    .DE(_00097_),
    .Q(\w[6][3] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][4]$_DFFE_PP_  (.D(_00539_),
    .DE(_00097_),
    .Q(\w[6][4] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][5]$_DFFE_PP_  (.D(_00540_),
    .DE(_00097_),
    .Q(\w[6][5] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][6]$_DFFE_PP_  (.D(_00541_),
    .DE(_00097_),
    .Q(\w[6][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][7]$_DFFE_PP_  (.D(_00542_),
    .DE(_00097_),
    .Q(\w[6][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][8]$_DFFE_PP_  (.D(_00543_),
    .DE(_00097_),
    .Q(\w[6][8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][9]$_DFFE_PP_  (.D(_00544_),
    .DE(_00097_),
    .Q(\w[6][9] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][0]$_DFFE_PP_  (.D(_00545_),
    .DE(net469),
    .Q(\w[7][0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][10]$_DFFE_PP_  (.D(_00546_),
    .DE(net468),
    .Q(\w[7][10] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][11]$_DFFE_PP_  (.D(_00547_),
    .DE(_00065_),
    .Q(\w[7][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][12]$_DFFE_PP_  (.D(_00548_),
    .DE(net469),
    .Q(\w[7][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][13]$_DFFE_PP_  (.D(_00549_),
    .DE(net468),
    .Q(\w[7][13] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][14]$_DFFE_PP_  (.D(_00550_),
    .DE(net467),
    .Q(\w[7][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][15]$_DFFE_PP_  (.D(_00551_),
    .DE(net469),
    .Q(\w[7][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][16]$_DFFE_PP_  (.D(_00552_),
    .DE(net467),
    .Q(\w[7][16] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][17]$_DFFE_PP_  (.D(_00553_),
    .DE(net467),
    .Q(\w[7][17] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][18]$_DFFE_PP_  (.D(_00554_),
    .DE(net468),
    .Q(\w[7][18] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][19]$_DFFE_PP_  (.D(_00555_),
    .DE(net468),
    .Q(\w[7][19] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][1]$_DFFE_PP_  (.D(_00556_),
    .DE(net469),
    .Q(\w[7][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][20]$_DFFE_PP_  (.D(_00557_),
    .DE(_00065_),
    .Q(\w[7][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][21]$_DFFE_PP_  (.D(_00558_),
    .DE(net468),
    .Q(\w[7][21] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][22]$_DFFE_PP_  (.D(_00559_),
    .DE(net468),
    .Q(\w[7][22] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][23]$_DFFE_PP_  (.D(_00560_),
    .DE(net467),
    .Q(\w[7][23] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][24]$_DFFE_PP_  (.D(_00561_),
    .DE(net467),
    .Q(\w[7][24] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][25]$_DFFE_PP_  (.D(_00562_),
    .DE(net467),
    .Q(\w[7][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][26]$_DFFE_PP_  (.D(_00563_),
    .DE(net467),
    .Q(\w[7][26] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][27]$_DFFE_PP_  (.D(_00564_),
    .DE(net467),
    .Q(\w[7][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][28]$_DFFE_PP_  (.D(_00565_),
    .DE(net468),
    .Q(\w[7][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][29]$_DFFE_PP_  (.D(_00566_),
    .DE(net468),
    .Q(\w[7][29] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][2]$_DFFE_PP_  (.D(_00567_),
    .DE(net467),
    .Q(\w[7][2] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][30]$_DFFE_PP_  (.D(_00568_),
    .DE(net468),
    .Q(\w[7][30] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][31]$_DFFE_PP_  (.D(_00569_),
    .DE(net468),
    .Q(\w[7][31] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][3]$_DFFE_PP_  (.D(_00570_),
    .DE(net469),
    .Q(\w[7][3] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][4]$_DFFE_PP_  (.D(_00571_),
    .DE(net469),
    .Q(\w[7][4] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][5]$_DFFE_PP_  (.D(_00572_),
    .DE(net469),
    .Q(\w[7][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][6]$_DFFE_PP_  (.D(_00573_),
    .DE(net468),
    .Q(\w[7][6] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][7]$_DFFE_PP_  (.D(_00574_),
    .DE(net469),
    .Q(\w[7][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][8]$_DFFE_PP_  (.D(_00575_),
    .DE(net467),
    .Q(\w[7][8] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][9]$_DFFE_PP_  (.D(_00576_),
    .DE(_00065_),
    .Q(\w[7][9] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][0]$_DFFE_PP_  (.D(_00577_),
    .DE(_00096_),
    .Q(\w[8][0] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][10]$_DFFE_PP_  (.D(_00578_),
    .DE(_00096_),
    .Q(\w[8][10] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][11]$_DFFE_PP_  (.D(_00579_),
    .DE(_00096_),
    .Q(\w[8][11] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][12]$_DFFE_PP_  (.D(_00580_),
    .DE(_00096_),
    .Q(\w[8][12] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][13]$_DFFE_PP_  (.D(_00581_),
    .DE(_00096_),
    .Q(\w[8][13] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][14]$_DFFE_PP_  (.D(_00582_),
    .DE(_00096_),
    .Q(\w[8][14] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][15]$_DFFE_PP_  (.D(_00583_),
    .DE(_00096_),
    .Q(\w[8][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][16]$_DFFE_PP_  (.D(_00584_),
    .DE(_00096_),
    .Q(\w[8][16] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][17]$_DFFE_PP_  (.D(_00585_),
    .DE(_00096_),
    .Q(\w[8][17] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][18]$_DFFE_PP_  (.D(_00586_),
    .DE(_00096_),
    .Q(\w[8][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][19]$_DFFE_PP_  (.D(_00587_),
    .DE(_00096_),
    .Q(\w[8][19] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][1]$_DFFE_PP_  (.D(_00588_),
    .DE(_00096_),
    .Q(\w[8][1] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][20]$_DFFE_PP_  (.D(_00589_),
    .DE(_00096_),
    .Q(\w[8][20] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][21]$_DFFE_PP_  (.D(_00590_),
    .DE(_00096_),
    .Q(\w[8][21] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][22]$_DFFE_PP_  (.D(_00591_),
    .DE(_00096_),
    .Q(\w[8][22] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][23]$_DFFE_PP_  (.D(_00592_),
    .DE(_00096_),
    .Q(\w[8][23] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][24]$_DFFE_PP_  (.D(_00593_),
    .DE(_00096_),
    .Q(\w[8][24] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][25]$_DFFE_PP_  (.D(_00594_),
    .DE(_00096_),
    .Q(\w[8][25] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][26]$_DFFE_PP_  (.D(_00595_),
    .DE(_00096_),
    .Q(\w[8][26] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][27]$_DFFE_PP_  (.D(_00596_),
    .DE(_00096_),
    .Q(\w[8][27] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][28]$_DFFE_PP_  (.D(_00597_),
    .DE(_00096_),
    .Q(\w[8][28] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][29]$_DFFE_PP_  (.D(_00598_),
    .DE(_00096_),
    .Q(\w[8][29] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][2]$_DFFE_PP_  (.D(_00599_),
    .DE(_00096_),
    .Q(\w[8][2] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][30]$_DFFE_PP_  (.D(_00600_),
    .DE(_00096_),
    .Q(\w[8][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][31]$_DFFE_PP_  (.D(_00601_),
    .DE(_00096_),
    .Q(\w[8][31] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][3]$_DFFE_PP_  (.D(_00602_),
    .DE(_00096_),
    .Q(\w[8][3] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][4]$_DFFE_PP_  (.D(_00603_),
    .DE(_00096_),
    .Q(\w[8][4] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][5]$_DFFE_PP_  (.D(_00604_),
    .DE(_00096_),
    .Q(\w[8][5] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][6]$_DFFE_PP_  (.D(_00605_),
    .DE(_00096_),
    .Q(\w[8][6] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][7]$_DFFE_PP_  (.D(_00606_),
    .DE(_00096_),
    .Q(\w[8][7] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][8]$_DFFE_PP_  (.D(_00607_),
    .DE(_00096_),
    .Q(\w[8][8] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][9]$_DFFE_PP_  (.D(_00608_),
    .DE(_00096_),
    .Q(\w[8][9] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][0]$_DFFE_PP_  (.D(_00609_),
    .DE(_00064_),
    .Q(\w[9][0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][10]$_DFFE_PP_  (.D(_00610_),
    .DE(_00064_),
    .Q(\w[9][10] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][11]$_DFFE_PP_  (.D(_00611_),
    .DE(_00064_),
    .Q(\w[9][11] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][12]$_DFFE_PP_  (.D(_00612_),
    .DE(_00064_),
    .Q(\w[9][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][13]$_DFFE_PP_  (.D(_00613_),
    .DE(_00064_),
    .Q(\w[9][13] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][14]$_DFFE_PP_  (.D(_00614_),
    .DE(_00064_),
    .Q(\w[9][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][15]$_DFFE_PP_  (.D(_00615_),
    .DE(_00064_),
    .Q(\w[9][15] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][16]$_DFFE_PP_  (.D(_00616_),
    .DE(_00064_),
    .Q(\w[9][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][17]$_DFFE_PP_  (.D(_00617_),
    .DE(_00064_),
    .Q(\w[9][17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][18]$_DFFE_PP_  (.D(_00618_),
    .DE(_00064_),
    .Q(\w[9][18] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][19]$_DFFE_PP_  (.D(_00619_),
    .DE(_00064_),
    .Q(\w[9][19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][1]$_DFFE_PP_  (.D(_00620_),
    .DE(_00064_),
    .Q(\w[9][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][20]$_DFFE_PP_  (.D(_00621_),
    .DE(_00064_),
    .Q(\w[9][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][21]$_DFFE_PP_  (.D(_00622_),
    .DE(_00064_),
    .Q(\w[9][21] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][22]$_DFFE_PP_  (.D(_00623_),
    .DE(_00064_),
    .Q(\w[9][22] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][23]$_DFFE_PP_  (.D(_00624_),
    .DE(_00064_),
    .Q(\w[9][23] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][24]$_DFFE_PP_  (.D(_00625_),
    .DE(_00064_),
    .Q(\w[9][24] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][25]$_DFFE_PP_  (.D(_00626_),
    .DE(_00064_),
    .Q(\w[9][25] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][26]$_DFFE_PP_  (.D(_00627_),
    .DE(_00064_),
    .Q(\w[9][26] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][27]$_DFFE_PP_  (.D(_00628_),
    .DE(_00064_),
    .Q(\w[9][27] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][28]$_DFFE_PP_  (.D(_00629_),
    .DE(_00064_),
    .Q(\w[9][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][29]$_DFFE_PP_  (.D(_00630_),
    .DE(_00064_),
    .Q(\w[9][29] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][2]$_DFFE_PP_  (.D(_00631_),
    .DE(_00064_),
    .Q(\w[9][2] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][30]$_DFFE_PP_  (.D(_00632_),
    .DE(_00064_),
    .Q(\w[9][30] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][31]$_DFFE_PP_  (.D(_00633_),
    .DE(_00064_),
    .Q(\w[9][31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][3]$_DFFE_PP_  (.D(_00634_),
    .DE(_00064_),
    .Q(\w[9][3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][4]$_DFFE_PP_  (.D(_00635_),
    .DE(_00064_),
    .Q(\w[9][4] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][5]$_DFFE_PP_  (.D(_00636_),
    .DE(_00064_),
    .Q(\w[9][5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][6]$_DFFE_PP_  (.D(_00637_),
    .DE(_00064_),
    .Q(\w[9][6] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][7]$_DFFE_PP_  (.D(_00638_),
    .DE(_00064_),
    .Q(\w[9][7] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][8]$_DFFE_PP_  (.D(_00639_),
    .DE(_00064_),
    .Q(\w[9][8] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][9]$_DFFE_PP_  (.D(_00640_),
    .DE(_00064_),
    .Q(\w[9][9] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[0]$_DFF_P_  (.D(_00000_),
    .Q(\hash.CA1.w_i1[0] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[10]$_DFF_P_  (.D(_00001_),
    .Q(\hash.CA1.w_i1[10] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[11]$_DFF_P_  (.D(_00002_),
    .Q(\hash.CA1.w_i1[11] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[12]$_DFF_P_  (.D(_00003_),
    .Q(\hash.CA1.w_i1[12] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[13]$_DFF_P_  (.D(_00004_),
    .Q(\hash.CA1.w_i1[13] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[14]$_DFF_P_  (.D(_00005_),
    .Q(\hash.CA1.w_i1[14] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[15]$_DFF_P_  (.D(_00006_),
    .Q(\hash.CA1.w_i1[15] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[16]$_DFF_P_  (.D(_00007_),
    .Q(\hash.CA1.w_i1[16] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[17]$_DFF_P_  (.D(_00008_),
    .Q(\hash.CA1.w_i1[17] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[18]$_DFF_P_  (.D(_00009_),
    .Q(\hash.CA1.w_i1[18] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[19]$_DFF_P_  (.D(_00010_),
    .Q(\hash.CA1.w_i1[19] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_2 \w_value1[1]$_DFF_P_  (.D(_00011_),
    .Q(\hash.CA1.w_i1[1] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_2 \w_value1[20]$_DFF_P_  (.D(_00012_),
    .Q(\hash.CA1.w_i1[20] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[21]$_DFF_P_  (.D(_00013_),
    .Q(\hash.CA1.w_i1[21] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[22]$_DFF_P_  (.D(_00014_),
    .Q(\hash.CA1.w_i1[22] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[23]$_DFF_P_  (.D(_00015_),
    .Q(\hash.CA1.w_i1[23] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 \w_value1[24]$_DFF_P_  (.D(_00016_),
    .Q(\hash.CA1.w_i1[24] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[25]$_DFF_P_  (.D(_00017_),
    .Q(\hash.CA1.w_i1[25] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[26]$_DFF_P_  (.D(_00018_),
    .Q(\hash.CA1.w_i1[26] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[27]$_DFF_P_  (.D(_00019_),
    .Q(\hash.CA1.w_i1[27] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[28]$_DFF_P_  (.D(_00020_),
    .Q(\hash.CA1.w_i1[28] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_2 \w_value1[29]$_DFF_P_  (.D(_00021_),
    .Q(\hash.CA1.w_i1[29] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[2]$_DFF_P_  (.D(_00022_),
    .Q(\hash.CA1.w_i1[2] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[30]$_DFF_P_  (.D(_00023_),
    .Q(\hash.CA1.w_i1[30] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[31]$_DFF_P_  (.D(_00024_),
    .Q(\hash.CA1.w_i1[31] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[3]$_DFF_P_  (.D(_00025_),
    .Q(\hash.CA1.w_i1[3] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_2 \w_value1[4]$_DFF_P_  (.D(_00026_),
    .Q(\hash.CA1.w_i1[4] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[5]$_DFF_P_  (.D(_00027_),
    .Q(\hash.CA1.w_i1[5] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[6]$_DFF_P_  (.D(_00028_),
    .Q(\hash.CA1.w_i1[6] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[7]$_DFF_P_  (.D(_00029_),
    .Q(\hash.CA1.w_i1[7] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[8]$_DFF_P_  (.D(_00030_),
    .Q(\hash.CA1.w_i1[8] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[9]$_DFF_P_  (.D(_00031_),
    .Q(\hash.CA1.w_i1[9] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[0]$_DFF_P_  (.D(_00032_),
    .Q(\hash.CA1.w_i2[0] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[10]$_DFF_P_  (.D(_00033_),
    .Q(\hash.CA1.w_i2[10] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[11]$_DFF_P_  (.D(_00034_),
    .Q(\hash.CA1.w_i2[11] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[12]$_DFF_P_  (.D(_00035_),
    .Q(\hash.CA1.w_i2[12] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[13]$_DFF_P_  (.D(_00036_),
    .Q(\hash.CA1.w_i2[13] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[14]$_DFF_P_  (.D(_00037_),
    .Q(\hash.CA1.w_i2[14] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[15]$_DFF_P_  (.D(_00038_),
    .Q(\hash.CA1.w_i2[15] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[16]$_DFF_P_  (.D(_00039_),
    .Q(\hash.CA1.w_i2[16] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[17]$_DFF_P_  (.D(_00040_),
    .Q(\hash.CA1.w_i2[17] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[18]$_DFF_P_  (.D(_00041_),
    .Q(\hash.CA1.w_i2[18] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[19]$_DFF_P_  (.D(_00042_),
    .Q(\hash.CA1.w_i2[19] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[1]$_DFF_P_  (.D(_00043_),
    .Q(\hash.CA1.w_i2[1] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[20]$_DFF_P_  (.D(_00044_),
    .Q(\hash.CA1.w_i2[20] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[21]$_DFF_P_  (.D(_00045_),
    .Q(\hash.CA1.w_i2[21] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[22]$_DFF_P_  (.D(_00046_),
    .Q(\hash.CA1.w_i2[22] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[23]$_DFF_P_  (.D(_00047_),
    .Q(\hash.CA1.w_i2[23] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[24]$_DFF_P_  (.D(_00048_),
    .Q(\hash.CA1.w_i2[24] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[25]$_DFF_P_  (.D(_00049_),
    .Q(\hash.CA1.w_i2[25] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[26]$_DFF_P_  (.D(_00050_),
    .Q(\hash.CA1.w_i2[26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[27]$_DFF_P_  (.D(_00051_),
    .Q(\hash.CA1.w_i2[27] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[28]$_DFF_P_  (.D(_00052_),
    .Q(\hash.CA1.w_i2[28] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[29]$_DFF_P_  (.D(_00053_),
    .Q(\hash.CA1.w_i2[29] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[2]$_DFF_P_  (.D(_00054_),
    .Q(\hash.CA1.w_i2[2] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[30]$_DFF_P_  (.D(_00055_),
    .Q(\hash.CA1.w_i2[30] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[31]$_DFF_P_  (.D(_00056_),
    .Q(\hash.CA1.w_i2[31] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[3]$_DFF_P_  (.D(_00057_),
    .Q(\hash.CA1.w_i2[3] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[4]$_DFF_P_  (.D(_00058_),
    .Q(\hash.CA1.w_i2[4] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[5]$_DFF_P_  (.D(_00059_),
    .Q(\hash.CA1.w_i2[5] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 \w_value2[6]$_DFF_P_  (.D(_00060_),
    .Q(\hash.CA1.w_i2[6] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[7]$_DFF_P_  (.D(_00061_),
    .Q(\hash.CA1.w_i2[7] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[8]$_DFF_P_  (.D(_00062_),
    .Q(\hash.CA1.w_i2[8] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[9]$_DFF_P_  (.D(_00063_),
    .Q(\hash.CA1.w_i2[9] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5196 ();
 sky130_fd_sc_hd__buf_12 load_slew453 (.A(net455),
    .X(net453));
 sky130_fd_sc_hd__buf_16 load_slew454 (.A(_10035_),
    .X(net454));
 sky130_fd_sc_hd__buf_16 load_slew455 (.A(_10035_),
    .X(net455));
 sky130_fd_sc_hd__buf_16 max_cap456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_12 wire457 (.A(net459),
    .X(net457));
 sky130_fd_sc_hd__buf_16 load_slew458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_16 load_slew459 (.A(_10564_),
    .X(net459));
 sky130_fd_sc_hd__buf_12 load_slew460 (.A(_10513_),
    .X(net460));
 sky130_fd_sc_hd__buf_16 load_slew461 (.A(net463),
    .X(net461));
 sky130_fd_sc_hd__buf_16 load_slew462 (.A(_10508_),
    .X(net462));
 sky130_fd_sc_hd__buf_12 max_cap463 (.A(_10508_),
    .X(net463));
 sky130_fd_sc_hd__buf_12 wire464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_12 load_slew465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_16 wire466 (.A(_10027_),
    .X(net466));
 sky130_fd_sc_hd__buf_8 wire467 (.A(net469),
    .X(net467));
 sky130_fd_sc_hd__buf_8 load_slew468 (.A(_00065_),
    .X(net468));
 sky130_fd_sc_hd__buf_16 max_cap469 (.A(_00065_),
    .X(net469));
 sky130_fd_sc_hd__buf_16 max_cap470 (.A(_00071_),
    .X(net470));
 sky130_fd_sc_hd__buf_16 max_cap471 (.A(_00071_),
    .X(net471));
 sky130_fd_sc_hd__buf_8 wire472 (.A(_00080_),
    .X(net472));
 sky130_fd_sc_hd__buf_16 max_cap473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_8 wire474 (.A(_00080_),
    .X(net474));
 sky130_fd_sc_hd__buf_12 wire475 (.A(_00088_),
    .X(net475));
 sky130_fd_sc_hd__buf_12 wire476 (.A(_00088_),
    .X(net476));
 sky130_fd_sc_hd__buf_12 load_slew477 (.A(net483),
    .X(net477));
 sky130_fd_sc_hd__buf_12 load_slew478 (.A(net483),
    .X(net478));
 sky130_fd_sc_hd__buf_12 load_slew479 (.A(net483),
    .X(net479));
 sky130_fd_sc_hd__buf_12 load_slew480 (.A(net482),
    .X(net480));
 sky130_fd_sc_hd__buf_16 load_slew481 (.A(_00655_),
    .X(net481));
 sky130_fd_sc_hd__buf_12 load_slew482 (.A(_00655_),
    .X(net482));
 sky130_fd_sc_hd__buf_12 load_slew483 (.A(_00655_),
    .X(net483));
 sky130_fd_sc_hd__buf_16 load_slew484 (.A(net488),
    .X(net484));
 sky130_fd_sc_hd__buf_12 load_slew485 (.A(net487),
    .X(net485));
 sky130_fd_sc_hd__buf_16 load_slew486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_16 load_slew487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_16 load_slew488 (.A(_00657_),
    .X(net488));
 sky130_fd_sc_hd__buf_16 load_slew489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_16 load_slew490 (.A(_10532_),
    .X(net490));
 sky130_fd_sc_hd__buf_16 max_cap491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_16 load_slew492 (.A(_10532_),
    .X(net492));
 sky130_fd_sc_hd__buf_16 load_slew493 (.A(_10503_),
    .X(net493));
 sky130_fd_sc_hd__buf_16 load_slew494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__buf_16 load_slew495 (.A(_10503_),
    .X(net495));
 sky130_fd_sc_hd__buf_16 load_slew496 (.A(net499),
    .X(net496));
 sky130_fd_sc_hd__buf_16 load_slew497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_12 max_cap498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_12 max_cap499 (.A(_10503_),
    .X(net499));
 sky130_fd_sc_hd__buf_16 load_slew500 (.A(net502),
    .X(net500));
 sky130_fd_sc_hd__buf_16 load_slew501 (.A(net503),
    .X(net501));
 sky130_fd_sc_hd__buf_16 load_slew502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_16 load_slew503 (.A(net507),
    .X(net503));
 sky130_fd_sc_hd__buf_12 wire504 (.A(_10499_),
    .X(net504));
 sky130_fd_sc_hd__buf_16 load_slew505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__buf_12 wire506 (.A(_10499_),
    .X(net506));
 sky130_fd_sc_hd__buf_12 load_slew507 (.A(_10499_),
    .X(net507));
 sky130_fd_sc_hd__buf_16 max_cap508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_16 max_cap509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_12 wire510 (.A(_10016_),
    .X(net510));
 sky130_fd_sc_hd__buf_12 max_cap511 (.A(net512),
    .X(net511));
 sky130_fd_sc_hd__buf_12 load_slew512 (.A(_10016_),
    .X(net512));
 sky130_fd_sc_hd__buf_16 wire513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_12 wire514 (.A(_10013_),
    .X(net514));
 sky130_fd_sc_hd__buf_12 load_slew515 (.A(_10013_),
    .X(net515));
 sky130_fd_sc_hd__buf_12 wire516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_12 load_slew517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__buf_12 load_slew518 (.A(_10013_),
    .X(net518));
 sky130_fd_sc_hd__buf_16 load_slew519 (.A(_06210_),
    .X(net519));
 sky130_fd_sc_hd__buf_16 load_slew520 (.A(\hash.reset ),
    .X(net520));
 sky130_fd_sc_hd__buf_16 load_slew521 (.A(net523),
    .X(net521));
 sky130_fd_sc_hd__buf_16 load_slew522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__buf_16 load_slew523 (.A(\hash.reset ),
    .X(net523));
 sky130_fd_sc_hd__buf_16 load_slew524 (.A(\hash.reset ),
    .X(net524));
 sky130_fd_sc_hd__buf_16 wire525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__buf_12 max_length526 (.A(reset_hash),
    .X(net526));
 sky130_fd_sc_hd__buf_16 load_slew527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__buf_16 load_slew528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__buf_16 load_slew529 (.A(net538),
    .X(net529));
 sky130_fd_sc_hd__buf_16 load_slew530 (.A(net538),
    .X(net530));
 sky130_fd_sc_hd__buf_6 load_slew531 (.A(net538),
    .X(net531));
 sky130_fd_sc_hd__buf_8 load_slew532 (.A(done),
    .X(net532));
 sky130_fd_sc_hd__buf_16 load_slew533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_16 load_slew534 (.A(net537),
    .X(net534));
 sky130_fd_sc_hd__buf_16 load_slew535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_8 load_slew536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_16 max_cap537 (.A(done),
    .X(net537));
 sky130_fd_sc_hd__buf_16 max_cap538 (.A(done),
    .X(net538));
 sky130_fd_sc_hd__buf_16 load_slew539 (.A(net544),
    .X(net539));
 sky130_fd_sc_hd__buf_12 load_slew540 (.A(net543),
    .X(net540));
 sky130_fd_sc_hd__buf_16 load_slew541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__buf_16 load_slew542 (.A(net543),
    .X(net542));
 sky130_fd_sc_hd__buf_16 max_cap543 (.A(net544),
    .X(net543));
 sky130_fd_sc_hd__buf_16 load_slew544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__buf_16 load_slew545 (.A(\count_hash2[1] ),
    .X(net545));
 sky130_fd_sc_hd__buf_16 load_slew546 (.A(net548),
    .X(net546));
 sky130_fd_sc_hd__buf_16 wire547 (.A(\count_hash1[1] ),
    .X(net547));
 sky130_fd_sc_hd__buf_12 load_slew548 (.A(\count_hash1[1] ),
    .X(net548));
 sky130_fd_sc_hd__buf_12 load_slew549 (.A(net552),
    .X(net549));
 sky130_fd_sc_hd__buf_12 load_slew550 (.A(net552),
    .X(net550));
 sky130_fd_sc_hd__buf_12 load_slew551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__buf_12 load_slew552 (.A(\count_hash1[1] ),
    .X(net552));
 sky130_fd_sc_hd__buf_16 max_cap553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_16 load_slew554 (.A(\count7_2[5] ),
    .X(net554));
 sky130_fd_sc_hd__buf_16 load_slew555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_16 load_slew556 (.A(\count7_2[4] ),
    .X(net556));
 sky130_fd_sc_hd__buf_12 load_slew557 (.A(net559),
    .X(net557));
 sky130_fd_sc_hd__buf_16 load_slew558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__buf_16 load_slew559 (.A(\count7_2[3] ),
    .X(net559));
 sky130_fd_sc_hd__buf_16 load_slew560 (.A(net566),
    .X(net560));
 sky130_fd_sc_hd__buf_12 load_slew561 (.A(net566),
    .X(net561));
 sky130_fd_sc_hd__buf_12 load_slew562 (.A(net566),
    .X(net562));
 sky130_fd_sc_hd__buf_16 load_slew563 (.A(net565),
    .X(net563));
 sky130_fd_sc_hd__buf_12 load_slew564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__buf_16 load_slew565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_16 load_slew566 (.A(\count7_2[2] ),
    .X(net566));
 sky130_fd_sc_hd__buf_16 load_slew567 (.A(\count7_2[1] ),
    .X(net567));
 sky130_fd_sc_hd__buf_12 load_slew568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__buf_16 load_slew569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_12 load_slew570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__buf_16 load_slew571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__buf_16 load_slew572 (.A(\count7_2[1] ),
    .X(net572));
 sky130_fd_sc_hd__buf_12 load_slew573 (.A(\count7_1[5] ),
    .X(net573));
 sky130_fd_sc_hd__buf_16 load_slew574 (.A(\count7_1[5] ),
    .X(net574));
 sky130_fd_sc_hd__buf_16 wire575 (.A(\count7_1[4] ),
    .X(net575));
 sky130_fd_sc_hd__buf_16 load_slew576 (.A(\count7_1[4] ),
    .X(net576));
 sky130_fd_sc_hd__buf_16 load_slew577 (.A(net579),
    .X(net577));
 sky130_fd_sc_hd__buf_12 load_slew578 (.A(\count7_1[3] ),
    .X(net578));
 sky130_fd_sc_hd__buf_12 load_slew579 (.A(\count7_1[3] ),
    .X(net579));
 sky130_fd_sc_hd__buf_12 load_slew580 (.A(net583),
    .X(net580));
 sky130_fd_sc_hd__buf_16 load_slew581 (.A(net583),
    .X(net581));
 sky130_fd_sc_hd__buf_12 load_slew582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__buf_16 load_slew583 (.A(\count7_1[2] ),
    .X(net583));
 sky130_fd_sc_hd__buf_12 load_slew584 (.A(net586),
    .X(net584));
 sky130_fd_sc_hd__buf_16 load_slew585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__buf_16 load_slew586 (.A(\count7_1[2] ),
    .X(net586));
 sky130_fd_sc_hd__buf_12 load_slew587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__buf_16 wire588 (.A(net590),
    .X(net588));
 sky130_fd_sc_hd__buf_16 load_slew589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__buf_16 wire590 (.A(\count7_1[1] ),
    .X(net590));
 sky130_fd_sc_hd__buf_16 load_slew591 (.A(\count7_1[1] ),
    .X(net591));
 sky130_fd_sc_hd__buf_16 wire592 (.A(\count2_2[5] ),
    .X(net592));
 sky130_fd_sc_hd__buf_16 load_slew593 (.A(\count2_2[5] ),
    .X(net593));
 sky130_fd_sc_hd__buf_16 wire594 (.A(\count2_2[4] ),
    .X(net594));
 sky130_fd_sc_hd__buf_12 load_slew595 (.A(\count2_2[4] ),
    .X(net595));
 sky130_fd_sc_hd__buf_12 load_slew596 (.A(\count2_2[3] ),
    .X(net596));
 sky130_fd_sc_hd__buf_12 load_slew597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__buf_12 load_slew598 (.A(\count2_2[3] ),
    .X(net598));
 sky130_fd_sc_hd__buf_16 load_slew599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_16 wire600 (.A(\count2_2[2] ),
    .X(net600));
 sky130_fd_sc_hd__buf_16 load_slew601 (.A(\count2_2[2] ),
    .X(net601));
 sky130_fd_sc_hd__buf_12 load_slew602 (.A(net604),
    .X(net602));
 sky130_fd_sc_hd__buf_16 load_slew603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__buf_16 load_slew604 (.A(\count2_2[2] ),
    .X(net604));
 sky130_fd_sc_hd__buf_12 load_slew605 (.A(net607),
    .X(net605));
 sky130_fd_sc_hd__buf_16 load_slew606 (.A(\count2_2[1] ),
    .X(net606));
 sky130_fd_sc_hd__buf_12 load_slew607 (.A(\count2_2[1] ),
    .X(net607));
 sky130_fd_sc_hd__buf_16 load_slew608 (.A(\count2_2[1] ),
    .X(net608));
 sky130_fd_sc_hd__buf_16 load_slew609 (.A(\count2_2[1] ),
    .X(net609));
 sky130_fd_sc_hd__buf_12 load_slew610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_16 wire611 (.A(\count2_1[5] ),
    .X(net611));
 sky130_fd_sc_hd__buf_12 load_slew612 (.A(net614),
    .X(net612));
 sky130_fd_sc_hd__buf_12 load_slew613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_12 load_slew614 (.A(\count2_1[4] ),
    .X(net614));
 sky130_fd_sc_hd__buf_12 load_slew615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__buf_16 load_slew616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__buf_16 load_slew617 (.A(\count2_1[3] ),
    .X(net617));
 sky130_fd_sc_hd__buf_16 load_slew618 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__buf_16 load_slew619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__buf_16 load_slew620 (.A(net623),
    .X(net620));
 sky130_fd_sc_hd__buf_16 load_slew621 (.A(net623),
    .X(net621));
 sky130_fd_sc_hd__buf_12 load_slew622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__buf_16 load_slew623 (.A(\count2_1[2] ),
    .X(net623));
 sky130_fd_sc_hd__buf_16 load_slew624 (.A(\count2_1[1] ),
    .X(net624));
 sky130_fd_sc_hd__buf_16 load_slew625 (.A(net628),
    .X(net625));
 sky130_fd_sc_hd__buf_16 load_slew626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__buf_16 wire627 (.A(\count2_1[1] ),
    .X(net627));
 sky130_fd_sc_hd__buf_16 load_slew628 (.A(\count2_1[1] ),
    .X(net628));
 sky130_fd_sc_hd__buf_12 load_slew629 (.A(\count16_2[5] ),
    .X(net629));
 sky130_fd_sc_hd__buf_12 load_slew630 (.A(\count16_2[5] ),
    .X(net630));
 sky130_fd_sc_hd__buf_16 load_slew631 (.A(\count16_2[4] ),
    .X(net631));
 sky130_fd_sc_hd__buf_12 load_slew632 (.A(\count16_2[4] ),
    .X(net632));
 sky130_fd_sc_hd__buf_12 load_slew633 (.A(\count16_2[3] ),
    .X(net633));
 sky130_fd_sc_hd__buf_16 load_slew634 (.A(\count16_2[3] ),
    .X(net634));
 sky130_fd_sc_hd__buf_16 load_slew635 (.A(net638),
    .X(net635));
 sky130_fd_sc_hd__buf_12 load_slew636 (.A(net639),
    .X(net636));
 sky130_fd_sc_hd__buf_16 load_slew637 (.A(net639),
    .X(net637));
 sky130_fd_sc_hd__buf_16 load_slew638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__buf_16 load_slew639 (.A(net641),
    .X(net639));
 sky130_fd_sc_hd__buf_16 load_slew640 (.A(\count16_2[2] ),
    .X(net640));
 sky130_fd_sc_hd__buf_12 load_slew641 (.A(\count16_2[2] ),
    .X(net641));
 sky130_fd_sc_hd__buf_16 load_slew642 (.A(\count16_2[1] ),
    .X(net642));
 sky130_fd_sc_hd__buf_16 load_slew643 (.A(net647),
    .X(net643));
 sky130_fd_sc_hd__buf_12 load_slew644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_16 load_slew645 (.A(net647),
    .X(net645));
 sky130_fd_sc_hd__buf_12 load_slew646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_16 load_slew647 (.A(\count16_2[1] ),
    .X(net647));
 sky130_fd_sc_hd__buf_16 load_slew648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__buf_16 load_slew649 (.A(\count16_1[5] ),
    .X(net649));
 sky130_fd_sc_hd__buf_16 load_slew650 (.A(\count16_1[4] ),
    .X(net650));
 sky130_fd_sc_hd__buf_12 load_slew651 (.A(\count16_1[4] ),
    .X(net651));
 sky130_fd_sc_hd__buf_16 wire652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_16 wire653 (.A(\count16_1[3] ),
    .X(net653));
 sky130_fd_sc_hd__buf_16 load_slew654 (.A(net658),
    .X(net654));
 sky130_fd_sc_hd__buf_12 load_slew655 (.A(net658),
    .X(net655));
 sky130_fd_sc_hd__buf_16 load_slew656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__buf_16 load_slew657 (.A(\count16_1[2] ),
    .X(net657));
 sky130_fd_sc_hd__buf_16 load_slew658 (.A(\count16_1[2] ),
    .X(net658));
 sky130_fd_sc_hd__buf_16 load_slew659 (.A(\count16_1[2] ),
    .X(net659));
 sky130_fd_sc_hd__buf_16 load_slew660 (.A(net663),
    .X(net660));
 sky130_fd_sc_hd__buf_16 load_slew661 (.A(net662),
    .X(net661));
 sky130_fd_sc_hd__buf_16 load_slew662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_16 load_slew663 (.A(\count16_1[1] ),
    .X(net663));
 sky130_fd_sc_hd__buf_12 load_slew664 (.A(\count16_1[1] ),
    .X(net664));
 sky130_fd_sc_hd__buf_12 load_slew665 (.A(\count15_2[5] ),
    .X(net665));
 sky130_fd_sc_hd__buf_12 load_slew666 (.A(\count15_2[5] ),
    .X(net666));
 sky130_fd_sc_hd__buf_16 load_slew667 (.A(\count15_2[4] ),
    .X(net667));
 sky130_fd_sc_hd__buf_16 wire668 (.A(\count15_2[4] ),
    .X(net668));
 sky130_fd_sc_hd__buf_16 wire669 (.A(\count15_2[3] ),
    .X(net669));
 sky130_fd_sc_hd__buf_12 load_slew670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__buf_12 load_slew671 (.A(\count15_2[3] ),
    .X(net671));
 sky130_fd_sc_hd__buf_16 wire672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__buf_16 max_cap673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__buf_16 load_slew674 (.A(\count15_2[2] ),
    .X(net674));
 sky130_fd_sc_hd__buf_16 load_slew675 (.A(net677),
    .X(net675));
 sky130_fd_sc_hd__buf_12 load_slew676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__buf_16 load_slew677 (.A(\count15_2[2] ),
    .X(net677));
 sky130_fd_sc_hd__buf_16 load_slew678 (.A(\count15_2[1] ),
    .X(net678));
 sky130_fd_sc_hd__buf_16 load_slew679 (.A(\count15_2[1] ),
    .X(net679));
 sky130_fd_sc_hd__buf_12 load_slew680 (.A(\count15_2[1] ),
    .X(net680));
 sky130_fd_sc_hd__buf_12 load_slew681 (.A(net682),
    .X(net681));
 sky130_fd_sc_hd__buf_16 load_slew682 (.A(\count15_2[1] ),
    .X(net682));
 sky130_fd_sc_hd__buf_16 load_slew683 (.A(\count15_1[5] ),
    .X(net683));
 sky130_fd_sc_hd__buf_16 load_slew684 (.A(\count15_1[5] ),
    .X(net684));
 sky130_fd_sc_hd__buf_16 wire685 (.A(\count15_1[4] ),
    .X(net685));
 sky130_fd_sc_hd__buf_12 load_slew686 (.A(\count15_1[4] ),
    .X(net686));
 sky130_fd_sc_hd__buf_12 load_slew687 (.A(\count15_1[3] ),
    .X(net687));
 sky130_fd_sc_hd__buf_16 load_slew688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__buf_12 load_slew689 (.A(\count15_1[3] ),
    .X(net689));
 sky130_fd_sc_hd__buf_12 load_slew690 (.A(net692),
    .X(net690));
 sky130_fd_sc_hd__buf_16 load_slew691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_16 load_slew692 (.A(\count15_1[2] ),
    .X(net692));
 sky130_fd_sc_hd__buf_12 load_slew693 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__buf_12 load_slew694 (.A(net696),
    .X(net694));
 sky130_fd_sc_hd__buf_12 load_slew695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__buf_16 load_slew696 (.A(\count15_1[2] ),
    .X(net696));
 sky130_fd_sc_hd__buf_16 load_slew697 (.A(\count15_1[1] ),
    .X(net697));
 sky130_fd_sc_hd__buf_12 load_slew698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__buf_16 load_slew699 (.A(\count15_1[1] ),
    .X(net699));
 sky130_fd_sc_hd__buf_16 load_slew700 (.A(\count15_1[1] ),
    .X(net700));
 sky130_fd_sc_hd__buf_12 load_slew701 (.A(\count15_1[1] ),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(message[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(message[100]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(message[101]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(message[102]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(message[103]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(message[104]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(message[105]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(message[106]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(message[107]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(message[108]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(message[109]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(message[10]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(message[110]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(message[111]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(message[112]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(message[113]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(message[114]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(message[115]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(message[116]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(message[117]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(message[118]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(message[119]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(message[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(message[120]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(message[121]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(message[122]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(message[123]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(message[124]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(message[125]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(message[126]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(message[127]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(message[128]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(message[129]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(message[12]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(message[130]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(message[131]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(message[132]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(message[133]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(message[134]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(message[135]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(message[136]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(message[137]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(message[138]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(message[139]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(message[13]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(message[140]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(message[141]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(message[142]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(message[143]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(message[144]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(message[145]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(message[146]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(message[147]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(message[148]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(message[149]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(message[14]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(message[150]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(message[151]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(message[152]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(message[153]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(message[154]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(message[155]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(message[156]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(message[157]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(message[158]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(message[159]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(message[15]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(message[160]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(message[161]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(message[162]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(message[163]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(message[164]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(message[165]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(message[166]),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input75 (.A(message[167]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(message[168]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(message[169]),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(message[16]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(message[170]),
    .X(net79));
 sky130_fd_sc_hd__buf_4 input80 (.A(message[171]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(message[172]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(message[173]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(message[174]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(message[175]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(message[176]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(message[177]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(message[178]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(message[179]),
    .X(net88));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(message[17]),
    .X(net89));
 sky130_fd_sc_hd__buf_4 input90 (.A(message[180]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(message[181]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(message[182]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(message[183]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(message[184]),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 input95 (.A(message[185]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(message[186]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(message[187]),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 input98 (.A(message[188]),
    .X(net98));
 sky130_fd_sc_hd__dlymetal6s2s_1 input99 (.A(message[189]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(message[18]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(message[190]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(message[191]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(message[192]),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 input104 (.A(message[193]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(message[194]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(message[195]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(message[196]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(message[197]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(message[198]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(message[199]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(message[19]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 input112 (.A(message[1]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(message[200]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(message[201]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(message[202]),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 input116 (.A(message[203]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 input117 (.A(message[204]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(message[205]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(message[206]),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 input120 (.A(message[207]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(message[208]),
    .X(net121));
 sky130_fd_sc_hd__dlymetal6s2s_1 input122 (.A(message[209]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(message[20]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(message[210]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(message[211]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(message[212]),
    .X(net126));
 sky130_fd_sc_hd__dlymetal6s2s_1 input127 (.A(message[213]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(message[214]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(message[215]),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 input130 (.A(message[216]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(message[217]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(message[218]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(message[219]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(message[21]),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 input135 (.A(message[220]),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input136 (.A(message[221]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(message[222]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(message[223]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(message[224]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(message[225]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(message[226]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(message[227]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(message[228]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(message[229]),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 input145 (.A(message[22]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(message[230]),
    .X(net146));
 sky130_fd_sc_hd__dlymetal6s2s_1 input147 (.A(message[231]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(message[232]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(message[233]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(message[234]),
    .X(net150));
 sky130_fd_sc_hd__buf_4 input151 (.A(message[235]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 input152 (.A(message[236]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(message[237]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(message[238]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(message[239]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 input156 (.A(message[23]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(message[240]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(message[241]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(message[242]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(message[243]),
    .X(net160));
 sky130_fd_sc_hd__buf_4 input161 (.A(message[244]),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(message[245]),
    .X(net162));
 sky130_fd_sc_hd__buf_4 input163 (.A(message[246]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(message[247]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(message[248]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(message[249]),
    .X(net166));
 sky130_fd_sc_hd__dlymetal6s2s_1 input167 (.A(message[24]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(message[250]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(message[251]),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 input170 (.A(message[252]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(message[253]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(message[254]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(message[255]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(message[256]),
    .X(net174));
 sky130_fd_sc_hd__buf_4 input175 (.A(message[257]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(message[258]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(message[259]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(message[25]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(message[260]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(message[261]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(message[262]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(message[263]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(message[264]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(message[265]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(message[266]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(message[267]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 input187 (.A(message[268]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(message[269]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(message[26]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(message[270]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(message[271]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 input192 (.A(message[272]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(message[273]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(message[274]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(message[275]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(message[276]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(message[277]),
    .X(net197));
 sky130_fd_sc_hd__buf_2 input198 (.A(message[278]),
    .X(net198));
 sky130_fd_sc_hd__dlymetal6s2s_1 input199 (.A(message[279]),
    .X(net199));
 sky130_fd_sc_hd__dlymetal6s2s_1 input200 (.A(message[27]),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 input201 (.A(message[280]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(message[281]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(message[282]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(message[283]),
    .X(net204));
 sky130_fd_sc_hd__dlymetal6s2s_1 input205 (.A(message[284]),
    .X(net205));
 sky130_fd_sc_hd__dlymetal6s2s_1 input206 (.A(message[285]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 input207 (.A(message[286]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(message[287]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(message[288]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(message[289]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(message[28]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(message[290]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(message[291]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(message[292]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(message[293]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(message[294]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(message[295]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(message[296]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(message[297]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input220 (.A(message[298]),
    .X(net220));
 sky130_fd_sc_hd__buf_4 input221 (.A(message[299]),
    .X(net221));
 sky130_fd_sc_hd__dlymetal6s2s_1 input222 (.A(message[29]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(message[2]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 input224 (.A(message[300]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(message[301]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(message[302]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(message[303]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(message[304]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 input229 (.A(message[305]),
    .X(net229));
 sky130_fd_sc_hd__buf_2 input230 (.A(message[306]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(message[307]),
    .X(net231));
 sky130_fd_sc_hd__buf_4 input232 (.A(message[308]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 input233 (.A(message[309]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(message[30]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 input235 (.A(message[310]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(message[311]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(message[312]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 input238 (.A(message[313]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(message[314]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input240 (.A(message[315]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(message[316]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 input242 (.A(message[317]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(message[318]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(message[319]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 input245 (.A(message[31]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(message[320]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 input247 (.A(message[321]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(message[322]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(message[323]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(message[324]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 input251 (.A(message[325]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(message[326]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(message[327]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input254 (.A(message[328]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 input255 (.A(message[329]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 input256 (.A(message[32]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 input257 (.A(message[330]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 input258 (.A(message[331]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 input259 (.A(message[332]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 input260 (.A(message[333]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 input261 (.A(message[334]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 input262 (.A(message[335]),
    .X(net262));
 sky130_fd_sc_hd__dlymetal6s2s_1 input263 (.A(message[336]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 input264 (.A(message[337]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 input265 (.A(message[338]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 input266 (.A(message[339]),
    .X(net266));
 sky130_fd_sc_hd__dlymetal6s2s_1 input267 (.A(message[33]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 input268 (.A(message[340]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 input269 (.A(message[341]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 input270 (.A(message[342]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 input271 (.A(message[343]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 input272 (.A(message[344]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 input273 (.A(message[345]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 input274 (.A(message[346]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 input275 (.A(message[347]),
    .X(net275));
 sky130_fd_sc_hd__dlymetal6s2s_1 input276 (.A(message[348]),
    .X(net276));
 sky130_fd_sc_hd__dlymetal6s2s_1 input277 (.A(message[349]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 input278 (.A(message[34]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 input279 (.A(message[350]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 input280 (.A(message[351]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 input281 (.A(message[352]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 input282 (.A(message[353]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 input283 (.A(message[354]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 input284 (.A(message[355]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 input285 (.A(message[356]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 input286 (.A(message[357]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 input287 (.A(message[358]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 input288 (.A(message[359]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 input289 (.A(message[35]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input290 (.A(message[360]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 input291 (.A(message[361]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 input292 (.A(message[362]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 input293 (.A(message[363]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 input294 (.A(message[364]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 input295 (.A(message[365]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 input296 (.A(message[366]),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 input297 (.A(message[367]),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 input298 (.A(message[368]),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 input299 (.A(message[369]),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 input300 (.A(message[36]),
    .X(net300));
 sky130_fd_sc_hd__buf_2 input301 (.A(message[370]),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 input302 (.A(message[371]),
    .X(net302));
 sky130_fd_sc_hd__buf_4 input303 (.A(message[372]),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 input304 (.A(message[373]),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 input305 (.A(message[374]),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 input306 (.A(message[375]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 input307 (.A(message[376]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 input308 (.A(message[377]),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 input309 (.A(message[378]),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 input310 (.A(message[379]),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 input311 (.A(message[37]),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 input312 (.A(message[380]),
    .X(net312));
 sky130_fd_sc_hd__buf_4 input313 (.A(message[381]),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 input314 (.A(message[382]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 input315 (.A(message[383]),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 input316 (.A(message[384]),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_4 input317 (.A(message[385]),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 input318 (.A(message[386]),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 input319 (.A(message[387]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 input320 (.A(message[388]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 input321 (.A(message[389]),
    .X(net321));
 sky130_fd_sc_hd__dlymetal6s2s_1 input322 (.A(message[38]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 input323 (.A(message[390]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 input324 (.A(message[391]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 input325 (.A(message[392]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 input326 (.A(message[393]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 input327 (.A(message[394]),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 input328 (.A(message[395]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_2 input329 (.A(message[396]),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 input330 (.A(message[397]),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 input331 (.A(message[398]),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 input332 (.A(message[399]),
    .X(net332));
 sky130_fd_sc_hd__dlymetal6s2s_1 input333 (.A(message[39]),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 input334 (.A(message[3]),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 input335 (.A(message[400]),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 input336 (.A(message[401]),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 input337 (.A(message[402]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 input338 (.A(message[403]),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 input339 (.A(message[404]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 input340 (.A(message[405]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 input341 (.A(message[406]),
    .X(net341));
 sky130_fd_sc_hd__dlymetal6s2s_1 input342 (.A(message[407]),
    .X(net342));
 sky130_fd_sc_hd__dlymetal6s2s_1 input343 (.A(message[408]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 input344 (.A(message[409]),
    .X(net344));
 sky130_fd_sc_hd__dlymetal6s2s_1 input345 (.A(message[40]),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 input346 (.A(message[410]),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_1 input347 (.A(message[411]),
    .X(net347));
 sky130_fd_sc_hd__dlymetal6s2s_1 input348 (.A(message[412]),
    .X(net348));
 sky130_fd_sc_hd__dlymetal6s2s_1 input349 (.A(message[413]),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 input350 (.A(message[414]),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 input351 (.A(message[415]),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 input352 (.A(message[416]),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 input353 (.A(message[417]),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 input354 (.A(message[418]),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 input355 (.A(message[419]),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 input356 (.A(message[41]),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 input357 (.A(message[420]),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 input358 (.A(message[421]),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 input359 (.A(message[422]),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 input360 (.A(message[423]),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 input361 (.A(message[424]),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 input362 (.A(message[425]),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 input363 (.A(message[426]),
    .X(net363));
 sky130_fd_sc_hd__buf_4 input364 (.A(message[427]),
    .X(net364));
 sky130_fd_sc_hd__dlymetal6s2s_1 input365 (.A(message[428]),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 input366 (.A(message[429]),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 input367 (.A(message[42]),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 input368 (.A(message[430]),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 input369 (.A(message[431]),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 input370 (.A(message[432]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 input371 (.A(message[433]),
    .X(net371));
 sky130_fd_sc_hd__buf_2 input372 (.A(message[434]),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 input373 (.A(message[435]),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_4 input374 (.A(message[436]),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 input375 (.A(message[437]),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_4 input376 (.A(message[438]),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 input377 (.A(message[439]),
    .X(net377));
 sky130_fd_sc_hd__buf_4 input378 (.A(message[43]),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 input379 (.A(message[440]),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 input380 (.A(message[441]),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 input381 (.A(message[442]),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 input382 (.A(message[443]),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 input383 (.A(message[444]),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 input384 (.A(message[445]),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_1 input385 (.A(message[446]),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 input386 (.A(message[447]),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 input387 (.A(message[448]),
    .X(net387));
 sky130_fd_sc_hd__buf_4 input388 (.A(message[449]),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 input389 (.A(message[44]),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 input390 (.A(message[450]),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 input391 (.A(message[451]),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 input392 (.A(message[452]),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_2 input393 (.A(message[453]),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 input394 (.A(message[454]),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 input395 (.A(message[455]),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 input396 (.A(message[456]),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 input397 (.A(message[457]),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 input398 (.A(message[458]),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 input399 (.A(message[459]),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 input400 (.A(message[45]),
    .X(net400));
 sky130_fd_sc_hd__dlymetal6s2s_1 input401 (.A(message[460]),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 input402 (.A(message[461]),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 input403 (.A(message[462]),
    .X(net403));
 sky130_fd_sc_hd__dlymetal6s2s_1 input404 (.A(message[463]),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 input405 (.A(message[464]),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 input406 (.A(message[465]),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 input407 (.A(message[466]),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_1 input408 (.A(message[467]),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 input409 (.A(message[468]),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 input410 (.A(message[469]),
    .X(net410));
 sky130_fd_sc_hd__buf_2 input411 (.A(message[46]),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 input412 (.A(message[470]),
    .X(net412));
 sky130_fd_sc_hd__dlymetal6s2s_1 input413 (.A(message[471]),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 input414 (.A(message[472]),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 input415 (.A(message[473]),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 input416 (.A(message[474]),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 input417 (.A(message[475]),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_1 input418 (.A(message[476]),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 input419 (.A(message[477]),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 input420 (.A(message[478]),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_1 input421 (.A(message[479]),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 input422 (.A(message[47]),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 input423 (.A(message[480]),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 input424 (.A(message[481]),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 input425 (.A(message[482]),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 input426 (.A(message[483]),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 input427 (.A(message[484]),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 input428 (.A(message[485]),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 input429 (.A(message[486]),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 input430 (.A(message[487]),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_1 input431 (.A(message[488]),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 input432 (.A(message[489]),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 input433 (.A(message[48]),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 input434 (.A(message[490]),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_4 input435 (.A(message[491]),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 input436 (.A(message[492]),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 input437 (.A(message[493]),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 input438 (.A(message[494]),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 input439 (.A(message[495]),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 input440 (.A(message[496]),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 input441 (.A(message[497]),
    .X(net441));
 sky130_fd_sc_hd__buf_2 input442 (.A(message[498]),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 input443 (.A(message[499]),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 input444 (.A(message[49]),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 input445 (.A(message[4]),
    .X(net445));
 sky130_fd_sc_hd__buf_4 input446 (.A(message[500]),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_2 input447 (.A(message[501]),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_4 input448 (.A(message[502]),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_1 input449 (.A(message[503]),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 input450 (.A(message[504]),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 input451 (.A(message[505]),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 input452 (.A(message[506]),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 input453 (.A(message[507]),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_1 input454 (.A(message[508]),
    .X(net703));
 sky130_fd_sc_hd__buf_4 input455 (.A(message[509]),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_4 input456 (.A(message[50]),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_1 input457 (.A(message[510]),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 input458 (.A(message[511]),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_1 input459 (.A(message[51]),
    .X(net708));
 sky130_fd_sc_hd__buf_4 input460 (.A(message[52]),
    .X(net709));
 sky130_fd_sc_hd__buf_2 input461 (.A(message[53]),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_4 input462 (.A(message[54]),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_1 input463 (.A(message[55]),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_1 input464 (.A(message[56]),
    .X(net713));
 sky130_fd_sc_hd__dlymetal6s2s_1 input465 (.A(message[57]),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_1 input466 (.A(message[58]),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_1 input467 (.A(message[59]),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 input468 (.A(message[5]),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_1 input469 (.A(message[60]),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_2 input470 (.A(message[61]),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_1 input471 (.A(message[62]),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_1 input472 (.A(message[63]),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_1 input473 (.A(message[64]),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_2 input474 (.A(message[65]),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_1 input475 (.A(message[66]),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_1 input476 (.A(message[67]),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_1 input477 (.A(message[68]),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_2 input478 (.A(message[69]),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_1 input479 (.A(message[6]),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_1 input480 (.A(message[70]),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 input481 (.A(message[71]),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_1 input482 (.A(message[72]),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 input483 (.A(message[73]),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 input484 (.A(message[74]),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 input485 (.A(message[75]),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_4 input486 (.A(message[76]),
    .X(net735));
 sky130_fd_sc_hd__dlymetal6s2s_1 input487 (.A(message[77]),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_2 input488 (.A(message[78]),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 input489 (.A(message[79]),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 input490 (.A(message[7]),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_2 input491 (.A(message[80]),
    .X(net740));
 sky130_fd_sc_hd__dlymetal6s2s_1 input492 (.A(message[81]),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 input493 (.A(message[82]),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_1 input494 (.A(message[83]),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 input495 (.A(message[84]),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_1 input496 (.A(message[85]),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 input497 (.A(message[86]),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_2 input498 (.A(message[87]),
    .X(net747));
 sky130_fd_sc_hd__dlymetal6s2s_1 input499 (.A(message[88]),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_1 input500 (.A(message[89]),
    .X(net749));
 sky130_fd_sc_hd__buf_4 input501 (.A(message[8]),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 input502 (.A(message[90]),
    .X(net751));
 sky130_fd_sc_hd__dlymetal6s2s_1 input503 (.A(message[91]),
    .X(net752));
 sky130_fd_sc_hd__dlymetal6s2s_1 input504 (.A(message[92]),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_2 input505 (.A(message[93]),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_1 input506 (.A(message[94]),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_1 input507 (.A(message[95]),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 input508 (.A(message[96]),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_1 input509 (.A(message[97]),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_1 input510 (.A(message[98]),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 input511 (.A(message[99]),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 input512 (.A(message[9]),
    .X(net761));
 sky130_fd_sc_hd__buf_16 input513 (.A(reset),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_1 output514 (.A(net763),
    .X(hashvalue[0]));
 sky130_fd_sc_hd__clkbuf_1 output515 (.A(net764),
    .X(hashvalue[100]));
 sky130_fd_sc_hd__clkbuf_1 output516 (.A(net765),
    .X(hashvalue[101]));
 sky130_fd_sc_hd__clkbuf_1 output517 (.A(net766),
    .X(hashvalue[102]));
 sky130_fd_sc_hd__clkbuf_1 output518 (.A(net767),
    .X(hashvalue[103]));
 sky130_fd_sc_hd__clkbuf_1 output519 (.A(net768),
    .X(hashvalue[104]));
 sky130_fd_sc_hd__clkbuf_1 output520 (.A(net769),
    .X(hashvalue[105]));
 sky130_fd_sc_hd__clkbuf_1 output521 (.A(net770),
    .X(hashvalue[106]));
 sky130_fd_sc_hd__clkbuf_1 output522 (.A(net771),
    .X(hashvalue[107]));
 sky130_fd_sc_hd__clkbuf_1 output523 (.A(net772),
    .X(hashvalue[108]));
 sky130_fd_sc_hd__clkbuf_1 output524 (.A(net773),
    .X(hashvalue[109]));
 sky130_fd_sc_hd__clkbuf_1 output525 (.A(net774),
    .X(hashvalue[10]));
 sky130_fd_sc_hd__clkbuf_1 output526 (.A(net775),
    .X(hashvalue[110]));
 sky130_fd_sc_hd__clkbuf_1 output527 (.A(net776),
    .X(hashvalue[111]));
 sky130_fd_sc_hd__clkbuf_1 output528 (.A(net777),
    .X(hashvalue[112]));
 sky130_fd_sc_hd__clkbuf_1 output529 (.A(net778),
    .X(hashvalue[113]));
 sky130_fd_sc_hd__clkbuf_1 output530 (.A(net779),
    .X(hashvalue[114]));
 sky130_fd_sc_hd__clkbuf_1 output531 (.A(net780),
    .X(hashvalue[115]));
 sky130_fd_sc_hd__clkbuf_1 output532 (.A(net781),
    .X(hashvalue[116]));
 sky130_fd_sc_hd__clkbuf_1 output533 (.A(net782),
    .X(hashvalue[117]));
 sky130_fd_sc_hd__clkbuf_1 output534 (.A(net783),
    .X(hashvalue[118]));
 sky130_fd_sc_hd__clkbuf_1 output535 (.A(net784),
    .X(hashvalue[119]));
 sky130_fd_sc_hd__clkbuf_1 output536 (.A(net785),
    .X(hashvalue[11]));
 sky130_fd_sc_hd__clkbuf_1 output537 (.A(net786),
    .X(hashvalue[120]));
 sky130_fd_sc_hd__clkbuf_1 output538 (.A(net787),
    .X(hashvalue[121]));
 sky130_fd_sc_hd__clkbuf_1 output539 (.A(net788),
    .X(hashvalue[122]));
 sky130_fd_sc_hd__clkbuf_1 output540 (.A(net789),
    .X(hashvalue[123]));
 sky130_fd_sc_hd__clkbuf_1 output541 (.A(net790),
    .X(hashvalue[124]));
 sky130_fd_sc_hd__clkbuf_1 output542 (.A(net791),
    .X(hashvalue[125]));
 sky130_fd_sc_hd__clkbuf_1 output543 (.A(net792),
    .X(hashvalue[126]));
 sky130_fd_sc_hd__clkbuf_1 output544 (.A(net793),
    .X(hashvalue[127]));
 sky130_fd_sc_hd__clkbuf_1 output545 (.A(net794),
    .X(hashvalue[128]));
 sky130_fd_sc_hd__clkbuf_1 output546 (.A(net795),
    .X(hashvalue[129]));
 sky130_fd_sc_hd__clkbuf_1 output547 (.A(net796),
    .X(hashvalue[12]));
 sky130_fd_sc_hd__clkbuf_1 output548 (.A(net797),
    .X(hashvalue[130]));
 sky130_fd_sc_hd__clkbuf_1 output549 (.A(net798),
    .X(hashvalue[131]));
 sky130_fd_sc_hd__clkbuf_1 output550 (.A(net799),
    .X(hashvalue[132]));
 sky130_fd_sc_hd__clkbuf_1 output551 (.A(net800),
    .X(hashvalue[133]));
 sky130_fd_sc_hd__clkbuf_1 output552 (.A(net801),
    .X(hashvalue[134]));
 sky130_fd_sc_hd__clkbuf_1 output553 (.A(net802),
    .X(hashvalue[135]));
 sky130_fd_sc_hd__clkbuf_1 output554 (.A(net803),
    .X(hashvalue[136]));
 sky130_fd_sc_hd__clkbuf_1 output555 (.A(net804),
    .X(hashvalue[137]));
 sky130_fd_sc_hd__clkbuf_1 output556 (.A(net805),
    .X(hashvalue[138]));
 sky130_fd_sc_hd__clkbuf_1 output557 (.A(net806),
    .X(hashvalue[139]));
 sky130_fd_sc_hd__clkbuf_1 output558 (.A(net807),
    .X(hashvalue[13]));
 sky130_fd_sc_hd__clkbuf_1 output559 (.A(net808),
    .X(hashvalue[140]));
 sky130_fd_sc_hd__clkbuf_1 output560 (.A(net809),
    .X(hashvalue[141]));
 sky130_fd_sc_hd__clkbuf_1 output561 (.A(net810),
    .X(hashvalue[142]));
 sky130_fd_sc_hd__clkbuf_1 output562 (.A(net811),
    .X(hashvalue[143]));
 sky130_fd_sc_hd__clkbuf_1 output563 (.A(net812),
    .X(hashvalue[144]));
 sky130_fd_sc_hd__clkbuf_1 output564 (.A(net813),
    .X(hashvalue[145]));
 sky130_fd_sc_hd__clkbuf_1 output565 (.A(net814),
    .X(hashvalue[146]));
 sky130_fd_sc_hd__clkbuf_1 output566 (.A(net815),
    .X(hashvalue[147]));
 sky130_fd_sc_hd__clkbuf_1 output567 (.A(net816),
    .X(hashvalue[148]));
 sky130_fd_sc_hd__clkbuf_1 output568 (.A(net817),
    .X(hashvalue[149]));
 sky130_fd_sc_hd__clkbuf_1 output569 (.A(net818),
    .X(hashvalue[14]));
 sky130_fd_sc_hd__clkbuf_1 output570 (.A(net819),
    .X(hashvalue[150]));
 sky130_fd_sc_hd__clkbuf_1 output571 (.A(net820),
    .X(hashvalue[151]));
 sky130_fd_sc_hd__clkbuf_1 output572 (.A(net821),
    .X(hashvalue[152]));
 sky130_fd_sc_hd__clkbuf_1 output573 (.A(net822),
    .X(hashvalue[153]));
 sky130_fd_sc_hd__clkbuf_1 output574 (.A(net823),
    .X(hashvalue[154]));
 sky130_fd_sc_hd__clkbuf_1 output575 (.A(net824),
    .X(hashvalue[155]));
 sky130_fd_sc_hd__clkbuf_1 output576 (.A(net825),
    .X(hashvalue[156]));
 sky130_fd_sc_hd__clkbuf_1 output577 (.A(net826),
    .X(hashvalue[157]));
 sky130_fd_sc_hd__clkbuf_1 output578 (.A(net827),
    .X(hashvalue[158]));
 sky130_fd_sc_hd__clkbuf_1 output579 (.A(net828),
    .X(hashvalue[159]));
 sky130_fd_sc_hd__clkbuf_1 output580 (.A(net829),
    .X(hashvalue[15]));
 sky130_fd_sc_hd__clkbuf_1 output581 (.A(net830),
    .X(hashvalue[160]));
 sky130_fd_sc_hd__clkbuf_1 output582 (.A(net831),
    .X(hashvalue[161]));
 sky130_fd_sc_hd__clkbuf_1 output583 (.A(net832),
    .X(hashvalue[162]));
 sky130_fd_sc_hd__clkbuf_1 output584 (.A(net833),
    .X(hashvalue[163]));
 sky130_fd_sc_hd__clkbuf_1 output585 (.A(net834),
    .X(hashvalue[164]));
 sky130_fd_sc_hd__clkbuf_1 output586 (.A(net835),
    .X(hashvalue[165]));
 sky130_fd_sc_hd__clkbuf_1 output587 (.A(net836),
    .X(hashvalue[166]));
 sky130_fd_sc_hd__clkbuf_1 output588 (.A(net837),
    .X(hashvalue[167]));
 sky130_fd_sc_hd__clkbuf_1 output589 (.A(net838),
    .X(hashvalue[168]));
 sky130_fd_sc_hd__clkbuf_1 output590 (.A(net839),
    .X(hashvalue[169]));
 sky130_fd_sc_hd__clkbuf_1 output591 (.A(net840),
    .X(hashvalue[16]));
 sky130_fd_sc_hd__clkbuf_1 output592 (.A(net841),
    .X(hashvalue[170]));
 sky130_fd_sc_hd__clkbuf_1 output593 (.A(net842),
    .X(hashvalue[171]));
 sky130_fd_sc_hd__clkbuf_1 output594 (.A(net843),
    .X(hashvalue[172]));
 sky130_fd_sc_hd__clkbuf_1 output595 (.A(net844),
    .X(hashvalue[173]));
 sky130_fd_sc_hd__clkbuf_1 output596 (.A(net845),
    .X(hashvalue[174]));
 sky130_fd_sc_hd__clkbuf_1 output597 (.A(net846),
    .X(hashvalue[175]));
 sky130_fd_sc_hd__clkbuf_1 output598 (.A(net847),
    .X(hashvalue[176]));
 sky130_fd_sc_hd__clkbuf_1 output599 (.A(net848),
    .X(hashvalue[177]));
 sky130_fd_sc_hd__clkbuf_1 output600 (.A(net849),
    .X(hashvalue[178]));
 sky130_fd_sc_hd__clkbuf_1 output601 (.A(net850),
    .X(hashvalue[179]));
 sky130_fd_sc_hd__clkbuf_1 output602 (.A(net851),
    .X(hashvalue[17]));
 sky130_fd_sc_hd__clkbuf_1 output603 (.A(net852),
    .X(hashvalue[180]));
 sky130_fd_sc_hd__clkbuf_1 output604 (.A(net853),
    .X(hashvalue[181]));
 sky130_fd_sc_hd__clkbuf_1 output605 (.A(net854),
    .X(hashvalue[182]));
 sky130_fd_sc_hd__clkbuf_1 output606 (.A(net855),
    .X(hashvalue[183]));
 sky130_fd_sc_hd__clkbuf_1 output607 (.A(net856),
    .X(hashvalue[184]));
 sky130_fd_sc_hd__clkbuf_1 output608 (.A(net857),
    .X(hashvalue[185]));
 sky130_fd_sc_hd__clkbuf_1 output609 (.A(net858),
    .X(hashvalue[186]));
 sky130_fd_sc_hd__clkbuf_1 output610 (.A(net859),
    .X(hashvalue[187]));
 sky130_fd_sc_hd__clkbuf_1 output611 (.A(net860),
    .X(hashvalue[188]));
 sky130_fd_sc_hd__clkbuf_1 output612 (.A(net861),
    .X(hashvalue[189]));
 sky130_fd_sc_hd__clkbuf_1 output613 (.A(net862),
    .X(hashvalue[18]));
 sky130_fd_sc_hd__clkbuf_1 output614 (.A(net863),
    .X(hashvalue[190]));
 sky130_fd_sc_hd__clkbuf_1 output615 (.A(net864),
    .X(hashvalue[191]));
 sky130_fd_sc_hd__clkbuf_1 output616 (.A(net865),
    .X(hashvalue[192]));
 sky130_fd_sc_hd__clkbuf_1 output617 (.A(net866),
    .X(hashvalue[193]));
 sky130_fd_sc_hd__clkbuf_1 output618 (.A(net867),
    .X(hashvalue[194]));
 sky130_fd_sc_hd__clkbuf_1 output619 (.A(net868),
    .X(hashvalue[195]));
 sky130_fd_sc_hd__clkbuf_1 output620 (.A(net869),
    .X(hashvalue[196]));
 sky130_fd_sc_hd__clkbuf_1 output621 (.A(net870),
    .X(hashvalue[197]));
 sky130_fd_sc_hd__clkbuf_1 output622 (.A(net871),
    .X(hashvalue[198]));
 sky130_fd_sc_hd__clkbuf_1 output623 (.A(net872),
    .X(hashvalue[199]));
 sky130_fd_sc_hd__clkbuf_1 output624 (.A(net873),
    .X(hashvalue[19]));
 sky130_fd_sc_hd__clkbuf_1 output625 (.A(net874),
    .X(hashvalue[1]));
 sky130_fd_sc_hd__clkbuf_1 output626 (.A(net875),
    .X(hashvalue[200]));
 sky130_fd_sc_hd__clkbuf_1 output627 (.A(net876),
    .X(hashvalue[201]));
 sky130_fd_sc_hd__clkbuf_1 output628 (.A(net877),
    .X(hashvalue[202]));
 sky130_fd_sc_hd__clkbuf_1 output629 (.A(net878),
    .X(hashvalue[203]));
 sky130_fd_sc_hd__clkbuf_1 output630 (.A(net879),
    .X(hashvalue[204]));
 sky130_fd_sc_hd__clkbuf_1 output631 (.A(net880),
    .X(hashvalue[205]));
 sky130_fd_sc_hd__clkbuf_1 output632 (.A(net881),
    .X(hashvalue[206]));
 sky130_fd_sc_hd__clkbuf_1 output633 (.A(net882),
    .X(hashvalue[207]));
 sky130_fd_sc_hd__clkbuf_1 output634 (.A(net883),
    .X(hashvalue[208]));
 sky130_fd_sc_hd__clkbuf_1 output635 (.A(net884),
    .X(hashvalue[209]));
 sky130_fd_sc_hd__clkbuf_1 output636 (.A(net885),
    .X(hashvalue[20]));
 sky130_fd_sc_hd__clkbuf_1 output637 (.A(net886),
    .X(hashvalue[210]));
 sky130_fd_sc_hd__clkbuf_1 output638 (.A(net887),
    .X(hashvalue[211]));
 sky130_fd_sc_hd__clkbuf_1 output639 (.A(net888),
    .X(hashvalue[212]));
 sky130_fd_sc_hd__clkbuf_1 output640 (.A(net889),
    .X(hashvalue[213]));
 sky130_fd_sc_hd__clkbuf_1 output641 (.A(net890),
    .X(hashvalue[214]));
 sky130_fd_sc_hd__clkbuf_1 output642 (.A(net891),
    .X(hashvalue[215]));
 sky130_fd_sc_hd__clkbuf_1 output643 (.A(net892),
    .X(hashvalue[216]));
 sky130_fd_sc_hd__clkbuf_1 output644 (.A(net893),
    .X(hashvalue[217]));
 sky130_fd_sc_hd__clkbuf_1 output645 (.A(net894),
    .X(hashvalue[218]));
 sky130_fd_sc_hd__clkbuf_1 output646 (.A(net895),
    .X(hashvalue[219]));
 sky130_fd_sc_hd__clkbuf_1 output647 (.A(net896),
    .X(hashvalue[21]));
 sky130_fd_sc_hd__clkbuf_1 output648 (.A(net897),
    .X(hashvalue[220]));
 sky130_fd_sc_hd__clkbuf_1 output649 (.A(net898),
    .X(hashvalue[221]));
 sky130_fd_sc_hd__clkbuf_1 output650 (.A(net899),
    .X(hashvalue[222]));
 sky130_fd_sc_hd__clkbuf_1 output651 (.A(net900),
    .X(hashvalue[223]));
 sky130_fd_sc_hd__clkbuf_1 output652 (.A(net901),
    .X(hashvalue[224]));
 sky130_fd_sc_hd__clkbuf_1 output653 (.A(net902),
    .X(hashvalue[225]));
 sky130_fd_sc_hd__clkbuf_1 output654 (.A(net903),
    .X(hashvalue[226]));
 sky130_fd_sc_hd__clkbuf_1 output655 (.A(net904),
    .X(hashvalue[227]));
 sky130_fd_sc_hd__clkbuf_1 output656 (.A(net905),
    .X(hashvalue[228]));
 sky130_fd_sc_hd__clkbuf_1 output657 (.A(net906),
    .X(hashvalue[229]));
 sky130_fd_sc_hd__clkbuf_1 output658 (.A(net907),
    .X(hashvalue[22]));
 sky130_fd_sc_hd__clkbuf_1 output659 (.A(net908),
    .X(hashvalue[230]));
 sky130_fd_sc_hd__clkbuf_1 output660 (.A(net909),
    .X(hashvalue[231]));
 sky130_fd_sc_hd__clkbuf_1 output661 (.A(net910),
    .X(hashvalue[232]));
 sky130_fd_sc_hd__clkbuf_1 output662 (.A(net911),
    .X(hashvalue[233]));
 sky130_fd_sc_hd__clkbuf_1 output663 (.A(net912),
    .X(hashvalue[234]));
 sky130_fd_sc_hd__clkbuf_1 output664 (.A(net913),
    .X(hashvalue[235]));
 sky130_fd_sc_hd__clkbuf_1 output665 (.A(net914),
    .X(hashvalue[236]));
 sky130_fd_sc_hd__clkbuf_1 output666 (.A(net915),
    .X(hashvalue[237]));
 sky130_fd_sc_hd__clkbuf_1 output667 (.A(net916),
    .X(hashvalue[238]));
 sky130_fd_sc_hd__clkbuf_1 output668 (.A(net917),
    .X(hashvalue[239]));
 sky130_fd_sc_hd__clkbuf_1 output669 (.A(net918),
    .X(hashvalue[23]));
 sky130_fd_sc_hd__clkbuf_1 output670 (.A(net919),
    .X(hashvalue[240]));
 sky130_fd_sc_hd__clkbuf_1 output671 (.A(net920),
    .X(hashvalue[241]));
 sky130_fd_sc_hd__clkbuf_1 output672 (.A(net921),
    .X(hashvalue[242]));
 sky130_fd_sc_hd__clkbuf_1 output673 (.A(net922),
    .X(hashvalue[243]));
 sky130_fd_sc_hd__clkbuf_1 output674 (.A(net923),
    .X(hashvalue[244]));
 sky130_fd_sc_hd__clkbuf_1 output675 (.A(net924),
    .X(hashvalue[245]));
 sky130_fd_sc_hd__clkbuf_1 output676 (.A(net925),
    .X(hashvalue[246]));
 sky130_fd_sc_hd__clkbuf_1 output677 (.A(net926),
    .X(hashvalue[247]));
 sky130_fd_sc_hd__clkbuf_1 output678 (.A(net927),
    .X(hashvalue[248]));
 sky130_fd_sc_hd__clkbuf_1 output679 (.A(net928),
    .X(hashvalue[249]));
 sky130_fd_sc_hd__clkbuf_1 output680 (.A(net929),
    .X(hashvalue[24]));
 sky130_fd_sc_hd__clkbuf_1 output681 (.A(net930),
    .X(hashvalue[250]));
 sky130_fd_sc_hd__clkbuf_1 output682 (.A(net931),
    .X(hashvalue[251]));
 sky130_fd_sc_hd__clkbuf_1 output683 (.A(net932),
    .X(hashvalue[252]));
 sky130_fd_sc_hd__clkbuf_1 output684 (.A(net933),
    .X(hashvalue[253]));
 sky130_fd_sc_hd__clkbuf_1 output685 (.A(net934),
    .X(hashvalue[254]));
 sky130_fd_sc_hd__clkbuf_1 output686 (.A(net935),
    .X(hashvalue[255]));
 sky130_fd_sc_hd__clkbuf_1 output687 (.A(net936),
    .X(hashvalue[25]));
 sky130_fd_sc_hd__clkbuf_1 output688 (.A(net937),
    .X(hashvalue[26]));
 sky130_fd_sc_hd__clkbuf_1 output689 (.A(net938),
    .X(hashvalue[27]));
 sky130_fd_sc_hd__clkbuf_1 output690 (.A(net939),
    .X(hashvalue[28]));
 sky130_fd_sc_hd__clkbuf_1 output691 (.A(net940),
    .X(hashvalue[29]));
 sky130_fd_sc_hd__clkbuf_1 output692 (.A(net941),
    .X(hashvalue[2]));
 sky130_fd_sc_hd__clkbuf_1 output693 (.A(net942),
    .X(hashvalue[30]));
 sky130_fd_sc_hd__clkbuf_1 output694 (.A(net943),
    .X(hashvalue[31]));
 sky130_fd_sc_hd__clkbuf_1 output695 (.A(net944),
    .X(hashvalue[32]));
 sky130_fd_sc_hd__clkbuf_1 output696 (.A(net945),
    .X(hashvalue[33]));
 sky130_fd_sc_hd__clkbuf_1 output697 (.A(net946),
    .X(hashvalue[34]));
 sky130_fd_sc_hd__clkbuf_1 output698 (.A(net947),
    .X(hashvalue[35]));
 sky130_fd_sc_hd__clkbuf_1 output699 (.A(net948),
    .X(hashvalue[36]));
 sky130_fd_sc_hd__clkbuf_1 output700 (.A(net949),
    .X(hashvalue[37]));
 sky130_fd_sc_hd__clkbuf_1 output701 (.A(net950),
    .X(hashvalue[38]));
 sky130_fd_sc_hd__clkbuf_1 output702 (.A(net951),
    .X(hashvalue[39]));
 sky130_fd_sc_hd__clkbuf_1 output703 (.A(net952),
    .X(hashvalue[3]));
 sky130_fd_sc_hd__clkbuf_1 output704 (.A(net953),
    .X(hashvalue[40]));
 sky130_fd_sc_hd__clkbuf_1 output705 (.A(net954),
    .X(hashvalue[41]));
 sky130_fd_sc_hd__clkbuf_1 output706 (.A(net955),
    .X(hashvalue[42]));
 sky130_fd_sc_hd__clkbuf_1 output707 (.A(net956),
    .X(hashvalue[43]));
 sky130_fd_sc_hd__clkbuf_1 output708 (.A(net957),
    .X(hashvalue[44]));
 sky130_fd_sc_hd__clkbuf_1 output709 (.A(net958),
    .X(hashvalue[45]));
 sky130_fd_sc_hd__clkbuf_1 output710 (.A(net959),
    .X(hashvalue[46]));
 sky130_fd_sc_hd__clkbuf_1 output711 (.A(net960),
    .X(hashvalue[47]));
 sky130_fd_sc_hd__clkbuf_1 output712 (.A(net961),
    .X(hashvalue[48]));
 sky130_fd_sc_hd__clkbuf_1 output713 (.A(net962),
    .X(hashvalue[49]));
 sky130_fd_sc_hd__clkbuf_1 output714 (.A(net963),
    .X(hashvalue[4]));
 sky130_fd_sc_hd__clkbuf_1 output715 (.A(net964),
    .X(hashvalue[50]));
 sky130_fd_sc_hd__clkbuf_1 output716 (.A(net965),
    .X(hashvalue[51]));
 sky130_fd_sc_hd__clkbuf_1 output717 (.A(net966),
    .X(hashvalue[52]));
 sky130_fd_sc_hd__clkbuf_1 output718 (.A(net967),
    .X(hashvalue[53]));
 sky130_fd_sc_hd__clkbuf_1 output719 (.A(net968),
    .X(hashvalue[54]));
 sky130_fd_sc_hd__clkbuf_1 output720 (.A(net969),
    .X(hashvalue[55]));
 sky130_fd_sc_hd__clkbuf_1 output721 (.A(net970),
    .X(hashvalue[56]));
 sky130_fd_sc_hd__clkbuf_1 output722 (.A(net971),
    .X(hashvalue[57]));
 sky130_fd_sc_hd__clkbuf_1 output723 (.A(net972),
    .X(hashvalue[58]));
 sky130_fd_sc_hd__clkbuf_1 output724 (.A(net973),
    .X(hashvalue[59]));
 sky130_fd_sc_hd__clkbuf_1 output725 (.A(net974),
    .X(hashvalue[5]));
 sky130_fd_sc_hd__clkbuf_1 output726 (.A(net975),
    .X(hashvalue[60]));
 sky130_fd_sc_hd__clkbuf_1 output727 (.A(net976),
    .X(hashvalue[61]));
 sky130_fd_sc_hd__clkbuf_1 output728 (.A(net977),
    .X(hashvalue[62]));
 sky130_fd_sc_hd__clkbuf_1 output729 (.A(net978),
    .X(hashvalue[63]));
 sky130_fd_sc_hd__clkbuf_1 output730 (.A(net979),
    .X(hashvalue[64]));
 sky130_fd_sc_hd__clkbuf_1 output731 (.A(net980),
    .X(hashvalue[65]));
 sky130_fd_sc_hd__clkbuf_1 output732 (.A(net981),
    .X(hashvalue[66]));
 sky130_fd_sc_hd__clkbuf_1 output733 (.A(net982),
    .X(hashvalue[67]));
 sky130_fd_sc_hd__clkbuf_1 output734 (.A(net983),
    .X(hashvalue[68]));
 sky130_fd_sc_hd__clkbuf_1 output735 (.A(net984),
    .X(hashvalue[69]));
 sky130_fd_sc_hd__clkbuf_1 output736 (.A(net985),
    .X(hashvalue[6]));
 sky130_fd_sc_hd__clkbuf_1 output737 (.A(net986),
    .X(hashvalue[70]));
 sky130_fd_sc_hd__clkbuf_1 output738 (.A(net987),
    .X(hashvalue[71]));
 sky130_fd_sc_hd__clkbuf_1 output739 (.A(net988),
    .X(hashvalue[72]));
 sky130_fd_sc_hd__clkbuf_1 output740 (.A(net989),
    .X(hashvalue[73]));
 sky130_fd_sc_hd__clkbuf_1 output741 (.A(net990),
    .X(hashvalue[74]));
 sky130_fd_sc_hd__clkbuf_1 output742 (.A(net991),
    .X(hashvalue[75]));
 sky130_fd_sc_hd__clkbuf_1 output743 (.A(net992),
    .X(hashvalue[76]));
 sky130_fd_sc_hd__clkbuf_1 output744 (.A(net993),
    .X(hashvalue[77]));
 sky130_fd_sc_hd__clkbuf_1 output745 (.A(net994),
    .X(hashvalue[78]));
 sky130_fd_sc_hd__clkbuf_1 output746 (.A(net995),
    .X(hashvalue[79]));
 sky130_fd_sc_hd__clkbuf_1 output747 (.A(net996),
    .X(hashvalue[7]));
 sky130_fd_sc_hd__clkbuf_1 output748 (.A(net997),
    .X(hashvalue[80]));
 sky130_fd_sc_hd__clkbuf_1 output749 (.A(net998),
    .X(hashvalue[81]));
 sky130_fd_sc_hd__clkbuf_1 output750 (.A(net999),
    .X(hashvalue[82]));
 sky130_fd_sc_hd__clkbuf_1 output751 (.A(net1000),
    .X(hashvalue[83]));
 sky130_fd_sc_hd__clkbuf_1 output752 (.A(net1001),
    .X(hashvalue[84]));
 sky130_fd_sc_hd__clkbuf_1 output753 (.A(net1002),
    .X(hashvalue[85]));
 sky130_fd_sc_hd__clkbuf_1 output754 (.A(net1003),
    .X(hashvalue[86]));
 sky130_fd_sc_hd__clkbuf_1 output755 (.A(net1004),
    .X(hashvalue[87]));
 sky130_fd_sc_hd__clkbuf_1 output756 (.A(net1005),
    .X(hashvalue[88]));
 sky130_fd_sc_hd__clkbuf_1 output757 (.A(net1006),
    .X(hashvalue[89]));
 sky130_fd_sc_hd__clkbuf_1 output758 (.A(net1007),
    .X(hashvalue[8]));
 sky130_fd_sc_hd__clkbuf_1 output759 (.A(net1008),
    .X(hashvalue[90]));
 sky130_fd_sc_hd__clkbuf_1 output760 (.A(net1009),
    .X(hashvalue[91]));
 sky130_fd_sc_hd__clkbuf_1 output761 (.A(net1010),
    .X(hashvalue[92]));
 sky130_fd_sc_hd__clkbuf_1 output762 (.A(net1011),
    .X(hashvalue[93]));
 sky130_fd_sc_hd__clkbuf_1 output763 (.A(net1012),
    .X(hashvalue[94]));
 sky130_fd_sc_hd__clkbuf_1 output764 (.A(net1013),
    .X(hashvalue[95]));
 sky130_fd_sc_hd__clkbuf_1 output765 (.A(net1014),
    .X(hashvalue[96]));
 sky130_fd_sc_hd__clkbuf_1 output766 (.A(net1015),
    .X(hashvalue[97]));
 sky130_fd_sc_hd__clkbuf_1 output767 (.A(net1016),
    .X(hashvalue[98]));
 sky130_fd_sc_hd__clkbuf_1 output768 (.A(net1017),
    .X(hashvalue[99]));
 sky130_fd_sc_hd__clkbuf_1 output769 (.A(net1018),
    .X(hashvalue[9]));
 sky130_fd_sc_hd__clkbuf_1 output770 (.A(net1019),
    .X(ready));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_274_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_275_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_278_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_280_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_282_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload0 (.A(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload1 (.A(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload2 (.A(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload3 (.A(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload5 (.A(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload7 (.A(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload8 (.A(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload10 (.A(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload11 (.A(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload12 (.A(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload13 (.A(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload14 (.A(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload15 (.A(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload16 (.A(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload17 (.A(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload18 (.A(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload19 (.A(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload20 (.A(clknet_leaf_268_clk));
 sky130_fd_sc_hd__bufinv_16 clkload21 (.A(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkinv_2 clkload22 (.A(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload23 (.A(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload24 (.A(clknet_leaf_280_clk));
 sky130_fd_sc_hd__bufinv_16 clkload25 (.A(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload26 (.A(clknet_leaf_282_clk));
 sky130_fd_sc_hd__clkinv_1 clkload27 (.A(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkinv_1 clkload28 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_1 clkload29 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_1 clkload30 (.A(clknet_leaf_253_clk));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkinv_1 clkload32 (.A(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload33 (.A(clknet_leaf_284_clk));
 sky130_fd_sc_hd__bufinv_16 clkload34 (.A(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkinv_1 clkload35 (.A(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkinv_2 clkload36 (.A(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload37 (.A(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkinv_1 clkload38 (.A(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkinv_1 clkload39 (.A(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkinv_2 clkload40 (.A(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkinv_2 clkload41 (.A(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkinv_2 clkload43 (.A(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkinv_2 clkload45 (.A(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkinv_2 clkload46 (.A(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload47 (.A(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkinv_1 clkload48 (.A(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload49 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload51 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkinv_2 clkload52 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkinv_2 clkload53 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload54 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload55 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinv_1 clkload56 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkinv_1 clkload57 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload58 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload59 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload60 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__bufinv_16 clkload61 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__bufinv_16 clkload63 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__bufinv_16 clkload64 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload65 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_2 clkload66 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload67 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkinv_1 clkload68 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkinv_1 clkload69 (.A(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload70 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload71 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload72 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinv_1 clkload73 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload74 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_1 clkload75 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload76 (.A(clknet_leaf_249_clk));
 sky130_fd_sc_hd__bufinv_16 clkload77 (.A(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload78 (.A(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkinv_1 clkload79 (.A(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload80 (.A(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkinv_2 clkload81 (.A(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkinv_2 clkload82 (.A(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkinv_2 clkload83 (.A(clknet_leaf_228_clk));
 sky130_fd_sc_hd__bufinv_16 clkload84 (.A(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkinv_2 clkload85 (.A(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkinv_1 clkload86 (.A(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload87 (.A(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkinv_1 clkload88 (.A(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkinv_1 clkload89 (.A(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload90 (.A(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload91 (.A(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkinv_2 clkload92 (.A(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload93 (.A(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkinv_1 clkload94 (.A(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkinv_2 clkload95 (.A(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkinv_1 clkload96 (.A(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkinv_2 clkload97 (.A(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload98 (.A(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload99 (.A(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkinv_1 clkload100 (.A(clknet_leaf_215_clk));
 sky130_fd_sc_hd__bufinv_16 clkload101 (.A(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkinv_1 clkload102 (.A(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload103 (.A(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkinv_2 clkload104 (.A(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkinv_1 clkload105 (.A(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload106 (.A(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkinv_2 clkload107 (.A(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload108 (.A(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkinv_1 clkload109 (.A(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload110 (.A(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload111 (.A(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload112 (.A(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload113 (.A(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload114 (.A(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload115 (.A(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload116 (.A(clknet_leaf_177_clk));
 sky130_fd_sc_hd__bufinv_16 clkload117 (.A(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkinv_2 clkload118 (.A(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload119 (.A(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload120 (.A(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkinv_2 clkload121 (.A(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkinv_1 clkload122 (.A(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkinv_1 clkload123 (.A(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload124 (.A(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkinv_1 clkload125 (.A(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkinv_2 clkload126 (.A(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkinv_4 clkload127 (.A(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload128 (.A(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkinv_2 clkload129 (.A(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkinv_1 clkload130 (.A(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload131 (.A(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkinv_2 clkload132 (.A(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkinv_2 clkload133 (.A(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload134 (.A(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload135 (.A(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkinv_2 clkload136 (.A(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload137 (.A(clknet_leaf_193_clk));
 sky130_fd_sc_hd__inv_4 clkload138 (.A(clknet_leaf_194_clk));
 sky130_fd_sc_hd__inv_4 clkload139 (.A(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkinv_1 clkload140 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload141 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload142 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinv_2 clkload143 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload144 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkinv_2 clkload145 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_2 clkload146 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload147 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload148 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkinv_2 clkload149 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__bufinv_16 clkload150 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkinv_4 clkload151 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload152 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload153 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__inv_6 clkload154 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__bufinv_16 clkload155 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_1 clkload156 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload157 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkinv_1 clkload158 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkinv_2 clkload159 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_2 clkload160 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload161 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_1 clkload162 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkinv_2 clkload163 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__bufinv_16 clkload164 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkinv_2 clkload165 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload166 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__bufinv_16 clkload167 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__bufinv_16 clkload168 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload169 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkinv_1 clkload170 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__bufinv_16 clkload171 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinv_2 clkload172 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkinv_1 clkload173 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkinv_2 clkload174 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkinv_2 clkload175 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload176 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload177 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkinv_1 clkload178 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkinv_1 clkload179 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkinv_1 clkload180 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinv_2 clkload181 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkinv_2 clkload182 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkinv_2 clkload183 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload184 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkinv_2 clkload185 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkinv_1 clkload186 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload187 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__bufinv_16 clkload188 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__bufinv_16 clkload189 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinv_2 clkload190 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkinv_1 clkload191 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__inv_6 clkload192 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__bufinv_16 clkload193 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_1 clkload194 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkinv_2 clkload195 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkinv_2 clkload196 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkinv_2 clkload197 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkinv_1 clkload198 (.A(clknet_leaf_166_clk));
 sky130_fd_sc_hd__bufinv_16 clkload199 (.A(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload200 (.A(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload201 (.A(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload202 (.A(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload203 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkinv_4 clkload204 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkinv_2 clkload205 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__bufinv_16 clkload206 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkinv_4 clkload207 (.A(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkinv_2 clkload208 (.A(clknet_leaf_169_clk));
 sky130_fd_sc_hd__bufinv_16 clkload209 (.A(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkinv_1 clkload210 (.A(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload211 (.A(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload212 (.A(clknet_leaf_161_clk));
 sky130_fd_sc_hd__bufinv_16 clkload213 (.A(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkinv_2 clkload214 (.A(clknet_leaf_163_clk));
 sky130_fd_sc_hd__bufinv_16 clkload215 (.A(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkinv_4 clkload216 (.A(clknet_leaf_165_clk));
 sky130_fd_sc_hd__bufinv_16 clkload217 (.A(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload218 (.A(clknet_leaf_148_clk));
 sky130_fd_sc_hd__inv_6 clkload219 (.A(clknet_leaf_149_clk));
 sky130_fd_sc_hd__bufinv_16 clkload220 (.A(clknet_leaf_150_clk));
 sky130_fd_sc_hd__inv_6 clkload221 (.A(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload222 (.A(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkinv_4 clkload223 (.A(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload224 (.A(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload225 (.A(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload226 (.A(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload227 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload228 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload229 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkinv_1 clkload230 (.A(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkinv_2 clkload231 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__inv_6 clkload232 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__inv_6 clkload233 (.A(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload234 (.A(clknet_leaf_132_clk));
 sky130_fd_sc_hd__inv_4 clkload235 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload236 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload237 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload238 (.A(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkinv_2 clkload239 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload240 (.A(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload241 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkinv_2 clkload242 (.A(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload243 (.A(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload244 (.A(clknet_leaf_131_clk));
 sky130_fd_sc_hd__bufinv_16 clkload245 (.A(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload246 (.A(clknet_leaf_134_clk));
 sky130_fd_sc_hd__bufinv_16 clkload247 (.A(clknet_leaf_135_clk));
 sky130_fd_sc_hd__bufinv_16 clkload248 (.A(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload249 (.A(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload250 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkinv_4 clkload251 (.A(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload252 (.A(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload253 (.A(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkinv_4 clkload254 (.A(clknet_leaf_140_clk));
 sky130_fd_sc_hd__bufinv_16 clkload255 (.A(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkinv_4 clkload256 (.A(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkinv_2 clkload257 (.A(clknet_leaf_143_clk));
 sky130_fd_sc_hd__nor2_4 clone1 (.A(net1021),
    .B(net523),
    .Y(net1020));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(_06881_),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_2 rebuffer3 (.A(net1033),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer133 (.A(_06895_),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_13399_),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(_13661_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer7 (.A(net1027),
    .X(net1026));
 sky130_fd_sc_hd__or3_2 clone8 (.A(net523),
    .B(net1156),
    .C(net1028),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(_06889_),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(_04681_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(\hash.CA2.S1.X[25] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(\hash.CA2.S1.X[25] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net1081),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1035),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net1036),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net1037),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1038),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1039),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1082),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net1043),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net1046),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net1054),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net1055),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net1056),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net1057),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_2 rebuffer39 (.A(net1062),
    .X(net1058));
 sky130_fd_sc_hd__buf_6 rebuffer40 (.A(_06862_),
    .X(net1108));
 sky130_fd_sc_hd__buf_6 rebuffer8 (.A(_06880_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer126 (.A(\hash.CA2.S1.X[27] ),
    .X(net1149));
 sky130_fd_sc_hd__buf_4 rebuffer43 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net1066),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net1068),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net1070),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(net1071),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__buf_2 rebuffer53 (.A(net1073),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(net1074),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net1075),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net1076),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_2 rebuffer57 (.A(net1077),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net1078),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(net1079),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(net1080),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer61 (.A(\hash.CA2.S1.X[25] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net1083),
    .X(net1081));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer63 (.A(net1106),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net1084),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net1086),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer67 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer68 (.A(net1088),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(\hash.CA2.S1.X[25] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(net1096),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(net1106),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer72 (.A(\hash.CA2.S1.X[6] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer73 (.A(net1091),
    .X(net1092));
 sky130_fd_sc_hd__buf_2 rebuffer74 (.A(net1092),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer75 (.A(\hash.CA2.S1.X[6] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer76 (.A(net1094),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(net1097),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer78 (.A(net1098),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer79 (.A(net1099),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(net1100),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer81 (.A(net1101),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer82 (.A(net1102),
    .X(net1101));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer83 (.A(\hash.CA2.S1.X[25] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer135 (.A(_04573_),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer85 (.A(_04861_),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 rebuffer86 (.A(_04861_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer91 (.A(_06874_),
    .X(net1110));
 sky130_fd_sc_hd__buf_2 rebuffer134 (.A(_06376_),
    .X(net1157));
 sky130_fd_sc_hd__buf_1 rebuffer93 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__buf_2 rebuffer94 (.A(net1109),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer99 (.A(_04782_),
    .X(net1118));
 sky130_fd_sc_hd__buf_8 rebuffer100 (.A(_04782_),
    .X(net1119));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer101 (.A(_04591_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer102 (.A(_04591_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer103 (.A(net1121),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer104 (.A(net1122),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer105 (.A(net1121),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer106 (.A(_04693_),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer107 (.A(_04573_),
    .X(net1126));
 sky130_fd_sc_hd__buf_6 rebuffer108 (.A(\hash.CA1.S0.X[23] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer109 (.A(net1127),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer110 (.A(_04672_),
    .X(net1129));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer111 (.A(_04672_),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer112 (.A(net1130),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer113 (.A(net1130),
    .X(net1132));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer114 (.A(_04652_),
    .X(net1133));
 sky130_fd_sc_hd__buf_2 rebuffer115 (.A(_04652_),
    .X(net1134));
 sky130_fd_sc_hd__buf_8 rebuffer116 (.A(_04652_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer117 (.A(_12252_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer118 (.A(_04733_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer119 (.A(_04762_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer120 (.A(net1138),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer121 (.A(net1139),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer122 (.A(net1140),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer123 (.A(net1141),
    .X(net1142));
 sky130_fd_sc_hd__buf_8 rebuffer1 (.A(\hash.CA2.S1.X[25] ),
    .X(net1106));
 sky130_fd_sc_hd__buf_1 rebuffer41 (.A(_07211_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer87 (.A(_13497_),
    .X(net1114));
 sky130_fd_sc_hd__buf_1 rebuffer88 (.A(_04901_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer127 (.A(\hash.CA2.S1.X[27] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer128 (.A(\hash.CA2.S1.X[27] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer129 (.A(net1151),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer136 (.A(_04824_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer137 (.A(net1159),
    .X(net1160));
 sky130_fd_sc_hd__buf_2 rebuffer138 (.A(_04824_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer139 (.A(net1161),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer140 (.A(net1161),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer141 (.A(_04667_),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer142 (.A(net1164),
    .X(net1165));
 sky130_fd_sc_hd__buf_12 rebuffer143 (.A(_04667_),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer144 (.A(_04643_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer145 (.A(net1167),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer146 (.A(net1168),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer147 (.A(_04643_),
    .X(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00014_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_00031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_00031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_00031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_00031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_00031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_00038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_00060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_00993_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_04261_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_08122_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_11944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_12086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_12134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_00810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_01020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_01024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_09148_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_09148_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_10328_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_11904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_12062_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_12086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_12545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_09148_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_09148_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1296 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1242 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_983 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_908 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_902 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_774 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1254 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1254 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_930 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1044 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1126 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_930 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1290 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1238 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1200 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1300 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1343 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1008 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1020 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1296 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1298 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1344 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1131 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1324 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_842 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_930 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1309 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1343 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1020 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1328 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1328 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1218 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1238 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1326 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1338 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1017 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1303 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1232 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1293 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1347 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1343 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_924 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1267 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1254 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1347 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1332 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_932 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1174 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_930 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1290 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1352 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_780 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1312 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1333 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1281 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1260 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_998 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1020 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1341 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1250 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1266 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1322 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1326 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1221 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1341 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1160 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_780 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1308 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1343 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1292 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1297 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1312 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1322 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1241 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1347 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1232 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1341 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1260 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1286 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1341 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1340 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_780 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1241 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_983 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1150 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1328 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_962 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1316 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1324 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1344 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1281 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_994 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1001 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1234 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1276 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1284 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1292 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_846 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_803 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1232 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1120 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1356 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1276 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1284 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1292 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1347 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1080 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1282 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1333 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_930 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1227 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1274 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_894 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1044 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1347 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1220 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1333 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1064 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1206 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1208 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_872 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1294 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1206 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1214 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1332 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1347 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1293 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1208 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1241 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1356 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1276 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1284 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1160 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1340 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1104 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1164 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1290 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1236 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1324 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_850 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1103 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1142 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1194 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_872 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1263 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_924 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1221 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1218 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_998 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1274 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1267 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_964 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_983 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1221 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1292 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1284 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1221 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1286 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1022 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1197 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1283 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1268 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1283 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1332 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1236 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1317 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1251 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1220 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1262 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1284 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1314 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1322 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1107 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_964 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1262 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1243 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1256 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1270 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_850 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1238 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1210 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1282 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_932 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_998 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1224 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1241 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1274 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1174 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1221 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1208 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1243 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1270 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1284 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1356 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_908 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_930 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1214 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1232 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1077 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1312 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1244 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1263 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1244 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1220 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1144 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1344 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1230 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1284 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1303 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1350 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1064 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1276 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1347 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1311 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1339 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1347 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_946 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1208 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1285 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1316 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1252 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1309 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1271 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1008 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_632 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_948 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1275 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1338 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1202 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1345 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1160 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1355 ();
endmodule
